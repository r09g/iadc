magic
tech sky130A
magscale 1 2
timestamp 1654583406
<< locali >>
rect 68283 100686 68317 100720
rect 68283 100614 68317 100652
rect 68283 100542 68317 100580
rect 68283 100470 68317 100508
rect 68283 100398 68317 100436
rect 68283 100326 68317 100364
rect 68283 100254 68317 100292
rect 68283 100182 68317 100220
rect 68283 100110 68317 100148
rect 68283 100038 68317 100076
rect 68283 99966 68317 100004
rect 68283 99894 68317 99932
rect 68283 99822 68317 99860
rect 68283 99750 68317 99788
rect 68283 99678 68317 99716
rect 68283 99606 68317 99644
rect 68283 99534 68317 99572
rect 68283 99462 68317 99500
rect 68283 99390 68317 99428
rect 68283 99318 68317 99356
rect 68283 99246 68317 99284
rect 68283 99174 68317 99212
rect 68283 99102 68317 99140
rect 68283 99030 68317 99068
rect 68283 98958 68317 98996
rect 68283 98886 68317 98924
rect 68283 98814 68317 98852
rect 68283 98742 68317 98780
rect 68283 98670 68317 98708
rect 68283 98598 68317 98636
rect 68283 98526 68317 98564
rect 68283 98454 68317 98492
rect 68283 98382 68317 98420
rect 68283 98310 68317 98348
rect 68283 98238 68317 98276
rect 68283 98166 68317 98204
rect 68283 98094 68317 98132
rect 68283 98022 68317 98060
rect 68283 97950 68317 97988
rect 68283 97878 68317 97916
rect 68283 97806 68317 97844
rect 68283 97734 68317 97772
rect 68283 97662 68317 97700
rect 68283 97590 68317 97628
rect 68283 97518 68317 97556
rect 68283 97450 68317 97484
rect 57471 84768 57571 84780
rect 57471 84734 57504 84768
rect 57538 84734 57571 84768
rect 57471 84696 57571 84734
rect 57471 84662 57504 84696
rect 57538 84662 57571 84696
rect 57471 84624 57571 84662
rect 57471 84590 57504 84624
rect 57538 84590 57571 84624
rect 57471 84552 57571 84590
rect 57471 84518 57504 84552
rect 57538 84518 57571 84552
rect 57471 84480 57571 84518
rect 57471 84446 57504 84480
rect 57538 84446 57571 84480
rect 57471 84408 57571 84446
rect 57471 84374 57504 84408
rect 57538 84374 57571 84408
rect 57471 84336 57571 84374
rect 57471 84302 57504 84336
rect 57538 84302 57571 84336
rect 57471 84264 57571 84302
rect 57471 84230 57504 84264
rect 57538 84230 57571 84264
rect 57471 84192 57571 84230
rect 57471 84158 57504 84192
rect 57538 84158 57571 84192
rect 57471 84120 57571 84158
rect 57471 84086 57504 84120
rect 57538 84086 57571 84120
rect 57471 84048 57571 84086
rect 57471 84014 57504 84048
rect 57538 84014 57571 84048
rect 57471 83976 57571 84014
rect 57471 83942 57504 83976
rect 57538 83942 57571 83976
rect 57471 83904 57571 83942
rect 57471 83870 57504 83904
rect 57538 83870 57571 83904
rect 57471 83832 57571 83870
rect 57471 83798 57504 83832
rect 57538 83798 57571 83832
rect 57471 83760 57571 83798
rect 57471 83726 57504 83760
rect 57538 83726 57571 83760
rect 57471 83688 57571 83726
rect 57471 83654 57504 83688
rect 57538 83654 57571 83688
rect 57471 83616 57571 83654
rect 57471 83582 57504 83616
rect 57538 83582 57571 83616
rect 57471 83544 57571 83582
rect 57471 83510 57504 83544
rect 57538 83510 57571 83544
rect 57471 83472 57571 83510
rect 57471 83438 57504 83472
rect 57538 83438 57571 83472
rect 57471 83400 57571 83438
rect 57471 83366 57504 83400
rect 57538 83366 57571 83400
rect 57471 83328 57571 83366
rect 57471 83294 57504 83328
rect 57538 83294 57571 83328
rect 57471 83256 57571 83294
rect 57471 83222 57504 83256
rect 57538 83222 57571 83256
rect 57471 83184 57571 83222
rect 57471 83150 57504 83184
rect 57538 83150 57571 83184
rect 57471 83112 57571 83150
rect 57471 83078 57504 83112
rect 57538 83078 57571 83112
rect 57471 83040 57571 83078
rect 57471 83006 57504 83040
rect 57538 83006 57571 83040
rect 57471 82968 57571 83006
rect 57471 82934 57504 82968
rect 57538 82934 57571 82968
rect 57471 82896 57571 82934
rect 57471 82862 57504 82896
rect 57538 82862 57571 82896
rect 57471 82824 57571 82862
rect 57471 82790 57504 82824
rect 57538 82790 57571 82824
rect 57471 82752 57571 82790
rect 57471 82718 57504 82752
rect 57538 82718 57571 82752
rect 57471 82680 57571 82718
rect 57471 82646 57504 82680
rect 57538 82646 57571 82680
rect 57471 82608 57571 82646
rect 57471 82574 57504 82608
rect 57538 82574 57571 82608
rect 57471 82536 57571 82574
rect 57471 82502 57504 82536
rect 57538 82502 57571 82536
rect 57471 82464 57571 82502
rect 57471 82430 57504 82464
rect 57538 82430 57571 82464
rect 57471 82392 57571 82430
rect 57471 82358 57504 82392
rect 57538 82358 57571 82392
rect 57471 82320 57571 82358
rect 57471 82286 57504 82320
rect 57538 82286 57571 82320
rect 57471 82248 57571 82286
rect 57471 82214 57504 82248
rect 57538 82214 57571 82248
rect 57471 82176 57571 82214
rect 57471 82142 57504 82176
rect 57538 82142 57571 82176
rect 57471 82104 57571 82142
rect 57471 82070 57504 82104
rect 57538 82070 57571 82104
rect 57471 82032 57571 82070
rect 57471 81998 57504 82032
rect 57538 81998 57571 82032
rect 57471 81960 57571 81998
rect 57471 81926 57504 81960
rect 57538 81926 57571 81960
rect 57471 81888 57571 81926
rect 57471 81854 57504 81888
rect 57538 81854 57571 81888
rect 57471 81816 57571 81854
rect 57471 81782 57504 81816
rect 57538 81782 57571 81816
rect 57471 81744 57571 81782
rect 57471 81710 57504 81744
rect 57538 81710 57571 81744
rect 57471 81672 57571 81710
rect 57471 81638 57504 81672
rect 57538 81638 57571 81672
rect 57471 81600 57571 81638
rect 57471 81566 57504 81600
rect 57538 81566 57571 81600
rect 57471 81528 57571 81566
rect 57471 81494 57504 81528
rect 57538 81494 57571 81528
rect 57471 81456 57571 81494
rect 57471 81422 57504 81456
rect 57538 81422 57571 81456
rect 57471 81384 57571 81422
rect 57471 81350 57504 81384
rect 57538 81350 57571 81384
rect 57471 81312 57571 81350
rect 57471 81278 57504 81312
rect 57538 81278 57571 81312
rect 57471 81240 57571 81278
rect 57471 81206 57504 81240
rect 57538 81206 57571 81240
rect 57471 81168 57571 81206
rect 57471 81134 57504 81168
rect 57538 81134 57571 81168
rect 57471 81096 57571 81134
rect 57471 81062 57504 81096
rect 57538 81062 57571 81096
rect 57471 81024 57571 81062
rect 57471 80990 57504 81024
rect 57538 80990 57571 81024
rect 57471 80952 57571 80990
rect 57471 80918 57504 80952
rect 57538 80918 57571 80952
rect 57471 80880 57571 80918
rect 57471 80846 57504 80880
rect 57538 80846 57571 80880
rect 57471 80808 57571 80846
rect 57471 80774 57504 80808
rect 57538 80774 57571 80808
rect 57471 80736 57571 80774
rect 57471 80702 57504 80736
rect 57538 80702 57571 80736
rect 57471 80664 57571 80702
rect 57471 80630 57504 80664
rect 57538 80630 57571 80664
rect 57471 80592 57571 80630
rect 57471 80558 57504 80592
rect 57538 80558 57571 80592
rect 57471 80520 57571 80558
rect 57471 80486 57504 80520
rect 57538 80486 57571 80520
rect 57471 80448 57571 80486
rect 57471 80414 57504 80448
rect 57538 80414 57571 80448
rect 57471 80376 57571 80414
rect 57471 80342 57504 80376
rect 57538 80342 57571 80376
rect 57471 80304 57571 80342
rect 57471 80270 57504 80304
rect 57538 80270 57571 80304
rect 57471 80232 57571 80270
rect 57471 80198 57504 80232
rect 57538 80198 57571 80232
rect 57471 80160 57571 80198
rect 57471 80126 57504 80160
rect 57538 80126 57571 80160
rect 57471 80088 57571 80126
rect 57471 80054 57504 80088
rect 57538 80054 57571 80088
rect 57471 80016 57571 80054
rect 57471 79982 57504 80016
rect 57538 79982 57571 80016
rect 57471 79944 57571 79982
rect 57471 79910 57504 79944
rect 57538 79910 57571 79944
rect 57471 79872 57571 79910
rect 57471 79838 57504 79872
rect 57538 79838 57571 79872
rect 57471 79800 57571 79838
rect 57471 79766 57504 79800
rect 57538 79766 57571 79800
rect 57471 79728 57571 79766
rect 57471 79694 57504 79728
rect 57538 79694 57571 79728
rect 57471 79656 57571 79694
rect 57471 79622 57504 79656
rect 57538 79622 57571 79656
rect 57471 79584 57571 79622
rect 57471 79550 57504 79584
rect 57538 79550 57571 79584
rect 57471 79512 57571 79550
rect 57471 79478 57504 79512
rect 57538 79478 57571 79512
rect 57471 79440 57571 79478
rect 57471 79406 57504 79440
rect 57538 79406 57571 79440
rect 57471 79368 57571 79406
rect 57471 79334 57504 79368
rect 57538 79334 57571 79368
rect 57471 79296 57571 79334
rect 57471 79262 57504 79296
rect 57538 79262 57571 79296
rect 57471 79224 57571 79262
rect 57471 79190 57504 79224
rect 57538 79190 57571 79224
rect 57471 79152 57571 79190
rect 57471 79118 57504 79152
rect 57538 79118 57571 79152
rect 57471 79080 57571 79118
rect 57471 79046 57504 79080
rect 57538 79046 57571 79080
rect 57471 79008 57571 79046
rect 57471 78974 57504 79008
rect 57538 78974 57571 79008
rect 57471 78936 57571 78974
rect 57471 78902 57504 78936
rect 57538 78902 57571 78936
rect 57471 78864 57571 78902
rect 57471 78830 57504 78864
rect 57538 78830 57571 78864
rect 57471 78792 57571 78830
rect 57471 78758 57504 78792
rect 57538 78758 57571 78792
rect 57471 78720 57571 78758
rect 57471 78686 57504 78720
rect 57538 78686 57571 78720
rect 57471 78648 57571 78686
rect 57471 78614 57504 78648
rect 57538 78614 57571 78648
rect 57471 78576 57571 78614
rect 57471 78542 57504 78576
rect 57538 78542 57571 78576
rect 57471 78504 57571 78542
rect 57471 78470 57504 78504
rect 57538 78470 57571 78504
rect 57471 78432 57571 78470
rect 57471 78398 57504 78432
rect 57538 78398 57571 78432
rect 57471 78360 57571 78398
rect 57471 78326 57504 78360
rect 57538 78326 57571 78360
rect 57471 78288 57571 78326
rect 57471 78254 57504 78288
rect 57538 78254 57571 78288
rect 57471 78216 57571 78254
rect 57471 78182 57504 78216
rect 57538 78182 57571 78216
rect 57471 78144 57571 78182
rect 57471 78110 57504 78144
rect 57538 78110 57571 78144
rect 57471 78072 57571 78110
rect 57471 78038 57504 78072
rect 57538 78038 57571 78072
rect 57471 78000 57571 78038
rect 57471 77966 57504 78000
rect 57538 77966 57571 78000
rect 57471 77928 57571 77966
rect 57471 77894 57504 77928
rect 57538 77894 57571 77928
rect 57471 77856 57571 77894
rect 57471 77822 57504 77856
rect 57538 77822 57571 77856
rect 57471 77784 57571 77822
rect 57471 77750 57504 77784
rect 57538 77750 57571 77784
rect 57471 77712 57571 77750
rect 57471 77678 57504 77712
rect 57538 77678 57571 77712
rect 57471 77640 57571 77678
rect 57471 77606 57504 77640
rect 57538 77606 57571 77640
rect 57471 77568 57571 77606
rect 57471 77534 57504 77568
rect 57538 77534 57571 77568
rect 57471 77496 57571 77534
rect 57471 77462 57504 77496
rect 57538 77462 57571 77496
rect 57471 77424 57571 77462
rect 57471 77390 57504 77424
rect 57538 77390 57571 77424
rect 57471 77352 57571 77390
rect 57471 77318 57504 77352
rect 57538 77318 57571 77352
rect 57471 77280 57571 77318
rect 57471 77246 57504 77280
rect 57538 77246 57571 77280
rect 57471 77208 57571 77246
rect 57471 77174 57504 77208
rect 57538 77174 57571 77208
rect 57471 77162 57571 77174
rect 51470 75010 56939 75040
rect 51470 74976 51487 75010
rect 51521 74976 51559 75010
rect 51593 74976 51631 75010
rect 51665 74976 51703 75010
rect 51737 74976 51775 75010
rect 51809 74976 51847 75010
rect 51881 74976 51919 75010
rect 51953 74976 51991 75010
rect 52025 74976 52063 75010
rect 52097 74976 52135 75010
rect 52169 74976 52207 75010
rect 52241 74976 52279 75010
rect 52313 74976 52351 75010
rect 52385 74976 52423 75010
rect 52457 74976 52495 75010
rect 52529 74976 52567 75010
rect 52601 74976 52639 75010
rect 52673 74976 52711 75010
rect 52745 74976 52783 75010
rect 52817 74976 52855 75010
rect 52889 74976 52927 75010
rect 52961 74976 52999 75010
rect 53033 74976 53071 75010
rect 53105 74976 53143 75010
rect 53177 74976 53215 75010
rect 53249 74976 53287 75010
rect 53321 74976 53359 75010
rect 53393 74976 53431 75010
rect 53465 74976 53503 75010
rect 53537 74976 53575 75010
rect 53609 74976 53647 75010
rect 53681 74976 53719 75010
rect 53753 74976 53791 75010
rect 53825 74976 53863 75010
rect 53897 74976 53935 75010
rect 53969 74976 54007 75010
rect 54041 74976 54079 75010
rect 54113 74976 54151 75010
rect 54185 74976 54223 75010
rect 54257 74976 54295 75010
rect 54329 74976 54367 75010
rect 54401 74976 54439 75010
rect 54473 74976 54511 75010
rect 54545 74976 54583 75010
rect 54617 74976 54655 75010
rect 54689 74976 54727 75010
rect 54761 74976 54799 75010
rect 54833 74976 54871 75010
rect 54905 74976 54943 75010
rect 54977 74976 55015 75010
rect 55049 74976 55087 75010
rect 55121 74976 55159 75010
rect 55193 74976 55231 75010
rect 55265 74976 55303 75010
rect 55337 74976 55375 75010
rect 55409 74976 55447 75010
rect 55481 74976 55519 75010
rect 55553 74976 55591 75010
rect 55625 74976 55663 75010
rect 55697 74976 55735 75010
rect 55769 74976 55807 75010
rect 55841 74976 55879 75010
rect 55913 74976 55951 75010
rect 55985 74976 56023 75010
rect 56057 74976 56095 75010
rect 56129 74976 56167 75010
rect 56201 74976 56239 75010
rect 56273 74976 56311 75010
rect 56345 74976 56383 75010
rect 56417 74976 56455 75010
rect 56489 74976 56527 75010
rect 56561 74976 56599 75010
rect 56633 74976 56671 75010
rect 56705 74976 56743 75010
rect 56777 74976 56815 75010
rect 56849 74976 56887 75010
rect 56921 74976 56939 75010
rect 51470 74947 56939 74976
rect 57090 74735 57183 74763
rect 57090 74701 57119 74735
rect 57153 74701 57183 74735
rect 57090 74663 57183 74701
rect 57090 74629 57119 74663
rect 57153 74629 57183 74663
rect 57090 74591 57183 74629
rect 57090 74557 57119 74591
rect 57153 74557 57183 74591
rect 57090 74519 57183 74557
rect 57090 74485 57119 74519
rect 57153 74485 57183 74519
rect 57090 74447 57183 74485
rect 57090 74413 57119 74447
rect 57153 74413 57183 74447
rect 57090 74375 57183 74413
rect 57090 74341 57119 74375
rect 57153 74341 57183 74375
rect 57090 74303 57183 74341
rect 57090 74269 57119 74303
rect 57153 74269 57183 74303
rect 57090 74231 57183 74269
rect 57090 74197 57119 74231
rect 57153 74197 57183 74231
rect 57090 74159 57183 74197
rect 57090 74125 57119 74159
rect 57153 74125 57183 74159
rect 57090 74087 57183 74125
rect 57090 74053 57119 74087
rect 57153 74053 57183 74087
rect 57090 74015 57183 74053
rect 57090 73981 57119 74015
rect 57153 73981 57183 74015
rect 57090 73943 57183 73981
rect 57090 73909 57119 73943
rect 57153 73909 57183 73943
rect 57090 73871 57183 73909
rect 57090 73837 57119 73871
rect 57153 73837 57183 73871
rect 57090 73799 57183 73837
rect 57090 73765 57119 73799
rect 57153 73765 57183 73799
rect 57090 73727 57183 73765
rect 57090 73693 57119 73727
rect 57153 73693 57183 73727
rect 57090 73655 57183 73693
rect 57090 73621 57119 73655
rect 57153 73621 57183 73655
rect 57090 73583 57183 73621
rect 57090 73549 57119 73583
rect 57153 73549 57183 73583
rect 57090 73511 57183 73549
rect 57090 73477 57119 73511
rect 57153 73477 57183 73511
rect 57090 73439 57183 73477
rect 30695 73420 30918 73426
rect 30695 73386 30717 73420
rect 30751 73386 30789 73420
rect 30823 73386 30861 73420
rect 30895 73386 30918 73420
rect 30695 73381 30918 73386
rect 57090 73405 57119 73439
rect 57153 73405 57183 73439
rect 57090 73367 57183 73405
rect 57090 73333 57119 73367
rect 57153 73333 57183 73367
rect 57090 73295 57183 73333
rect 57090 73261 57119 73295
rect 57153 73261 57183 73295
rect 57090 73223 57183 73261
rect 57090 73189 57119 73223
rect 57153 73189 57183 73223
rect 57090 73151 57183 73189
rect 57090 73117 57119 73151
rect 57153 73117 57183 73151
rect 57090 73079 57183 73117
rect 57090 73045 57119 73079
rect 57153 73045 57183 73079
rect 57090 73007 57183 73045
rect 57090 72973 57119 73007
rect 57153 72973 57183 73007
rect 57090 72935 57183 72973
rect 57090 72901 57119 72935
rect 57153 72901 57183 72935
rect 57090 72863 57183 72901
rect 57090 72829 57119 72863
rect 57153 72829 57183 72863
rect 57090 72791 57183 72829
rect 57090 72757 57119 72791
rect 57153 72757 57183 72791
rect 57090 72719 57183 72757
rect 57090 72685 57119 72719
rect 57153 72685 57183 72719
rect 57090 72647 57183 72685
rect 57090 72613 57119 72647
rect 57153 72613 57183 72647
rect 57090 72575 57183 72613
rect 57090 72541 57119 72575
rect 57153 72541 57183 72575
rect 57090 72503 57183 72541
rect 57090 72469 57119 72503
rect 57153 72469 57183 72503
rect 57090 72431 57183 72469
rect 57090 72397 57119 72431
rect 57153 72397 57183 72431
rect 57090 72359 57183 72397
rect 57090 72325 57119 72359
rect 57153 72325 57183 72359
rect 57090 72287 57183 72325
rect 57090 72253 57119 72287
rect 57153 72253 57183 72287
rect 57090 72215 57183 72253
rect 57090 72181 57119 72215
rect 57153 72181 57183 72215
rect 57090 72143 57183 72181
rect 57090 72109 57119 72143
rect 57153 72109 57183 72143
rect 57090 72071 57183 72109
rect 57090 72037 57119 72071
rect 57153 72037 57183 72071
rect 57090 71999 57183 72037
rect 57090 71965 57119 71999
rect 57153 71965 57183 71999
rect 57090 71927 57183 71965
rect 57090 71893 57119 71927
rect 57153 71893 57183 71927
rect 57090 71855 57183 71893
rect 57090 71821 57119 71855
rect 57153 71821 57183 71855
rect 57090 71793 57183 71821
rect 57471 69807 57571 69840
rect 57471 69773 57504 69807
rect 57538 69773 57571 69807
rect 57471 69735 57571 69773
rect 57471 69701 57504 69735
rect 57538 69701 57571 69735
rect 57471 69663 57571 69701
rect 57471 69629 57504 69663
rect 57538 69629 57571 69663
rect 57471 69591 57571 69629
rect 57471 69557 57504 69591
rect 57538 69557 57571 69591
rect 57471 69519 57571 69557
rect 57471 69485 57504 69519
rect 57538 69485 57571 69519
rect 57471 69447 57571 69485
rect 57471 69413 57504 69447
rect 57538 69413 57571 69447
rect 57471 69375 57571 69413
rect 57471 69341 57504 69375
rect 57538 69341 57571 69375
rect 57471 69303 57571 69341
rect 57471 69269 57504 69303
rect 57538 69269 57571 69303
rect 57471 69231 57571 69269
rect 57471 69197 57504 69231
rect 57538 69197 57571 69231
rect 57471 69159 57571 69197
rect 57471 69125 57504 69159
rect 57538 69125 57571 69159
rect 57471 69087 57571 69125
rect 57471 69053 57504 69087
rect 57538 69053 57571 69087
rect 57471 69015 57571 69053
rect 57471 68981 57504 69015
rect 57538 68981 57571 69015
rect 57471 68943 57571 68981
rect 57471 68909 57504 68943
rect 57538 68909 57571 68943
rect 57471 68871 57571 68909
rect 57471 68837 57504 68871
rect 57538 68837 57571 68871
rect 98902 68949 98936 68958
rect 98902 68877 98936 68915
rect 57471 68799 57571 68837
rect 57471 68765 57504 68799
rect 57538 68765 57571 68799
rect 98902 68805 98936 68843
rect 57471 68727 57571 68765
rect 57471 68693 57504 68727
rect 57538 68693 57571 68727
rect 98902 68733 98936 68771
rect 100097 68808 100132 68840
rect 100131 68774 100132 68808
rect 99631 68735 99633 68769
rect 99667 68735 99705 68769
rect 99739 68735 99777 68769
rect 99811 68735 99849 68769
rect 99883 68735 99921 68769
rect 99955 68735 99993 68769
rect 100027 68735 100030 68769
rect 100097 68736 100132 68774
rect 100347 68738 100371 68772
rect 100405 68738 100443 68772
rect 100477 68738 100502 68772
rect 57471 68655 57571 68693
rect 57471 68621 57504 68655
rect 57538 68621 57571 68655
rect 57471 68583 57571 68621
rect 98902 68661 98936 68699
rect 100131 68702 100132 68736
rect 100097 68670 100132 68702
rect 98902 68618 98936 68627
rect 57471 68549 57504 68583
rect 57538 68549 57571 68583
rect 57471 68511 57571 68549
rect 57471 68477 57504 68511
rect 57538 68477 57571 68511
rect 57471 68439 57571 68477
rect 57471 68405 57504 68439
rect 57538 68405 57571 68439
rect 57471 68372 57571 68405
rect 98902 67799 98936 67808
rect 98902 67727 98936 67765
rect 98902 67655 98936 67693
rect 98902 67583 98936 67621
rect 100097 67658 100132 67690
rect 100131 67624 100132 67658
rect 99631 67585 99633 67619
rect 99667 67585 99705 67619
rect 99739 67585 99777 67619
rect 99811 67585 99849 67619
rect 99883 67585 99921 67619
rect 99955 67585 99993 67619
rect 100027 67585 100030 67619
rect 100097 67586 100132 67624
rect 100347 67588 100371 67622
rect 100405 67588 100443 67622
rect 100477 67588 100502 67622
rect 98902 67511 98936 67549
rect 100131 67552 100132 67586
rect 100097 67520 100132 67552
rect 98902 67468 98936 67477
rect 57471 65348 57571 65365
rect 57471 65314 57504 65348
rect 57538 65314 57571 65348
rect 57471 65276 57571 65314
rect 57471 65242 57504 65276
rect 57538 65242 57571 65276
rect 57471 65204 57571 65242
rect 57471 65170 57504 65204
rect 57538 65170 57571 65204
rect 57471 65132 57571 65170
rect 98902 65259 98936 65268
rect 98902 65187 98936 65225
rect 57471 65098 57504 65132
rect 57538 65098 57571 65132
rect 98902 65115 98936 65153
rect 57471 65060 57571 65098
rect 57471 65026 57504 65060
rect 57538 65026 57571 65060
rect 98902 65043 98936 65081
rect 100097 65118 100132 65150
rect 100131 65084 100132 65118
rect 99631 65045 99633 65079
rect 99667 65045 99705 65079
rect 99739 65045 99777 65079
rect 99811 65045 99849 65079
rect 99883 65045 99921 65079
rect 99955 65045 99993 65079
rect 100027 65045 100030 65079
rect 100097 65046 100132 65084
rect 100347 65048 100371 65082
rect 100405 65048 100443 65082
rect 100477 65048 100502 65082
rect 57471 64988 57571 65026
rect 57471 64954 57504 64988
rect 57538 64954 57571 64988
rect 57471 64916 57571 64954
rect 98902 64971 98936 65009
rect 100131 65012 100132 65046
rect 100097 64980 100132 65012
rect 98902 64928 98936 64937
rect 57471 64882 57504 64916
rect 57538 64882 57571 64916
rect 57471 64844 57571 64882
rect 57471 64810 57504 64844
rect 57538 64810 57571 64844
rect 57471 64772 57571 64810
rect 57471 64738 57504 64772
rect 57538 64738 57571 64772
rect 57471 64700 57571 64738
rect 57471 64666 57504 64700
rect 57538 64666 57571 64700
rect 57471 64628 57571 64666
rect 57471 64594 57504 64628
rect 57538 64594 57571 64628
rect 57471 64556 57571 64594
rect 57471 64522 57504 64556
rect 57538 64522 57571 64556
rect 57471 64484 57571 64522
rect 57471 64450 57504 64484
rect 57538 64450 57571 64484
rect 57471 64412 57571 64450
rect 57471 64378 57504 64412
rect 57538 64378 57571 64412
rect 57471 64340 57571 64378
rect 57471 64306 57504 64340
rect 57538 64306 57571 64340
rect 57471 64268 57571 64306
rect 57471 64234 57504 64268
rect 57538 64234 57571 64268
rect 57471 64196 57571 64234
rect 57471 64162 57504 64196
rect 57538 64162 57571 64196
rect 57471 64124 57571 64162
rect 57471 64090 57504 64124
rect 57538 64090 57571 64124
rect 57471 64073 57571 64090
rect 98902 63989 98936 63998
rect 98902 63917 98936 63955
rect 98902 63845 98936 63883
rect 51457 63795 56926 63825
rect 51457 63761 51474 63795
rect 51508 63761 51546 63795
rect 51580 63761 51618 63795
rect 51652 63761 51690 63795
rect 51724 63761 51762 63795
rect 51796 63761 51834 63795
rect 51868 63761 51906 63795
rect 51940 63761 51978 63795
rect 52012 63761 52050 63795
rect 52084 63761 52122 63795
rect 52156 63761 52194 63795
rect 52228 63761 52266 63795
rect 52300 63761 52338 63795
rect 52372 63761 52410 63795
rect 52444 63761 52482 63795
rect 52516 63761 52554 63795
rect 52588 63761 52626 63795
rect 52660 63761 52698 63795
rect 52732 63761 52770 63795
rect 52804 63761 52842 63795
rect 52876 63761 52914 63795
rect 52948 63761 52986 63795
rect 53020 63761 53058 63795
rect 53092 63761 53130 63795
rect 53164 63761 53202 63795
rect 53236 63761 53274 63795
rect 53308 63761 53346 63795
rect 53380 63761 53418 63795
rect 53452 63761 53490 63795
rect 53524 63761 53562 63795
rect 53596 63761 53634 63795
rect 53668 63761 53706 63795
rect 53740 63761 53778 63795
rect 53812 63761 53850 63795
rect 53884 63761 53922 63795
rect 53956 63761 53994 63795
rect 54028 63761 54066 63795
rect 54100 63761 54138 63795
rect 54172 63761 54210 63795
rect 54244 63761 54282 63795
rect 54316 63761 54354 63795
rect 54388 63761 54426 63795
rect 54460 63761 54498 63795
rect 54532 63761 54570 63795
rect 54604 63761 54642 63795
rect 54676 63761 54714 63795
rect 54748 63761 54786 63795
rect 54820 63761 54858 63795
rect 54892 63761 54930 63795
rect 54964 63761 55002 63795
rect 55036 63761 55074 63795
rect 55108 63761 55146 63795
rect 55180 63761 55218 63795
rect 55252 63761 55290 63795
rect 55324 63761 55362 63795
rect 55396 63761 55434 63795
rect 55468 63761 55506 63795
rect 55540 63761 55578 63795
rect 55612 63761 55650 63795
rect 55684 63761 55722 63795
rect 55756 63761 55794 63795
rect 55828 63761 55866 63795
rect 55900 63761 55938 63795
rect 55972 63761 56010 63795
rect 56044 63761 56082 63795
rect 56116 63761 56154 63795
rect 56188 63761 56226 63795
rect 56260 63761 56298 63795
rect 56332 63761 56370 63795
rect 56404 63761 56442 63795
rect 56476 63761 56514 63795
rect 56548 63761 56586 63795
rect 56620 63761 56658 63795
rect 56692 63761 56730 63795
rect 56764 63761 56802 63795
rect 56836 63761 56874 63795
rect 56908 63761 56926 63795
rect 98902 63773 98936 63811
rect 100097 63848 100132 63880
rect 100131 63814 100132 63848
rect 99631 63775 99633 63809
rect 99667 63775 99705 63809
rect 99739 63775 99777 63809
rect 99811 63775 99849 63809
rect 99883 63775 99921 63809
rect 99955 63775 99993 63809
rect 100027 63775 100030 63809
rect 100097 63776 100132 63814
rect 100347 63778 100371 63812
rect 100405 63778 100443 63812
rect 100477 63778 100502 63812
rect 51457 63732 56926 63761
rect 98902 63701 98936 63739
rect 100131 63742 100132 63776
rect 100097 63710 100132 63742
rect 98902 63658 98936 63667
rect 25299 63136 25333 63154
rect 25299 63064 25333 63102
rect 25299 62992 25333 63030
rect 25299 62920 25333 62958
rect 25299 62868 25333 62886
rect 25299 62572 25333 62598
rect 25299 62500 25333 62538
rect 25299 62428 25333 62466
rect 25299 62356 25333 62394
rect 25299 62284 25333 62322
rect 25299 62224 25333 62250
rect 57153 40139 57246 40157
rect 57153 40105 57182 40139
rect 57216 40105 57246 40139
rect 57153 40067 57246 40105
rect 57153 40033 57182 40067
rect 57216 40033 57246 40067
rect 57153 39995 57246 40033
rect 57153 39961 57182 39995
rect 57216 39961 57246 39995
rect 57153 39923 57246 39961
rect 57153 39889 57182 39923
rect 57216 39889 57246 39923
rect 57153 39851 57246 39889
rect 57153 39817 57182 39851
rect 57216 39817 57246 39851
rect 57153 39779 57246 39817
rect 57153 39745 57182 39779
rect 57216 39745 57246 39779
rect 57153 39707 57246 39745
rect 57153 39673 57182 39707
rect 57216 39673 57246 39707
rect 57153 39635 57246 39673
rect 57153 39601 57182 39635
rect 57216 39601 57246 39635
rect 57153 39563 57246 39601
rect 57153 39529 57182 39563
rect 57216 39529 57246 39563
rect 57153 39491 57246 39529
rect 57153 39457 57182 39491
rect 57216 39457 57246 39491
rect 57153 39419 57246 39457
rect 57153 39385 57182 39419
rect 57216 39385 57246 39419
rect 57153 39347 57246 39385
rect 57153 39313 57182 39347
rect 57216 39313 57246 39347
rect 57153 39275 57246 39313
rect 57153 39241 57182 39275
rect 57216 39241 57246 39275
rect 57153 39203 57246 39241
rect 57153 39169 57182 39203
rect 57216 39169 57246 39203
rect 57153 39131 57246 39169
rect 57153 39097 57182 39131
rect 57216 39097 57246 39131
rect 57153 39059 57246 39097
rect 57153 39025 57182 39059
rect 57216 39025 57246 39059
rect 57153 38987 57246 39025
rect 57153 38953 57182 38987
rect 57216 38953 57246 38987
rect 57153 38915 57246 38953
rect 57153 38881 57182 38915
rect 57216 38881 57246 38915
rect 57153 38843 57246 38881
rect 57153 38809 57182 38843
rect 57216 38809 57246 38843
rect 57153 38771 57246 38809
rect 57153 38737 57182 38771
rect 57216 38737 57246 38771
rect 57153 38699 57246 38737
rect 57153 38665 57182 38699
rect 57216 38665 57246 38699
rect 57153 38627 57246 38665
rect 57153 38593 57182 38627
rect 57216 38593 57246 38627
rect 57153 38555 57246 38593
rect 57153 38521 57182 38555
rect 57216 38521 57246 38555
rect 57153 38483 57246 38521
rect 57153 38449 57182 38483
rect 57216 38449 57246 38483
rect 68368 40110 68397 40144
rect 68431 40110 68461 40144
rect 68368 40072 68461 40110
rect 68368 40038 68397 40072
rect 68431 40038 68461 40072
rect 68368 40000 68461 40038
rect 68368 39966 68397 40000
rect 68431 39966 68461 40000
rect 68368 39928 68461 39966
rect 68368 39894 68397 39928
rect 68431 39894 68461 39928
rect 68368 39856 68461 39894
rect 68368 39822 68397 39856
rect 68431 39822 68461 39856
rect 68368 39784 68461 39822
rect 68368 39750 68397 39784
rect 68431 39750 68461 39784
rect 68368 39712 68461 39750
rect 68368 39678 68397 39712
rect 68431 39678 68461 39712
rect 68368 39640 68461 39678
rect 68368 39606 68397 39640
rect 68431 39606 68461 39640
rect 68368 39568 68461 39606
rect 68368 39534 68397 39568
rect 68431 39534 68461 39568
rect 68368 39496 68461 39534
rect 68368 39462 68397 39496
rect 68431 39462 68461 39496
rect 68368 39424 68461 39462
rect 68368 39390 68397 39424
rect 68431 39390 68461 39424
rect 68368 39352 68461 39390
rect 68368 39318 68397 39352
rect 68431 39318 68461 39352
rect 68368 39280 68461 39318
rect 68368 39246 68397 39280
rect 68431 39246 68461 39280
rect 68368 39208 68461 39246
rect 68368 39174 68397 39208
rect 68431 39174 68461 39208
rect 68368 39136 68461 39174
rect 68368 39102 68397 39136
rect 68431 39102 68461 39136
rect 68368 39064 68461 39102
rect 68368 39030 68397 39064
rect 68431 39030 68461 39064
rect 68368 38992 68461 39030
rect 68368 38958 68397 38992
rect 68431 38958 68461 38992
rect 68368 38920 68461 38958
rect 68368 38886 68397 38920
rect 68431 38886 68461 38920
rect 68368 38848 68461 38886
rect 68368 38814 68397 38848
rect 68431 38814 68461 38848
rect 68368 38776 68461 38814
rect 68368 38742 68397 38776
rect 68431 38742 68461 38776
rect 68368 38704 68461 38742
rect 68368 38670 68397 38704
rect 68431 38670 68461 38704
rect 68368 38632 68461 38670
rect 68368 38598 68397 38632
rect 68431 38598 68461 38632
rect 68368 38560 68461 38598
rect 68368 38526 68397 38560
rect 68431 38526 68461 38560
rect 68368 38488 68461 38526
rect 68368 38454 68397 38488
rect 68431 38454 68461 38488
rect 57153 38411 57246 38449
rect 57153 38377 57182 38411
rect 57216 38377 57246 38411
rect 57153 38339 57246 38377
rect 57153 38305 57182 38339
rect 57216 38305 57246 38339
rect 57153 38267 57246 38305
rect 57153 38233 57182 38267
rect 57216 38233 57246 38267
rect 57153 38195 57246 38233
rect 57153 38161 57182 38195
rect 57216 38161 57246 38195
rect 57153 38123 57246 38161
rect 57153 38089 57182 38123
rect 57216 38089 57246 38123
rect 57153 38051 57246 38089
rect 57153 38017 57182 38051
rect 57216 38017 57246 38051
rect 57153 37979 57246 38017
rect 57153 37945 57182 37979
rect 57216 37945 57246 37979
rect 57153 37907 57246 37945
rect 57153 37873 57182 37907
rect 57216 37873 57246 37907
rect 57153 37835 57246 37873
rect 57153 37801 57182 37835
rect 57216 37801 57246 37835
rect 57153 37763 57246 37801
rect 57153 37729 57182 37763
rect 57216 37729 57246 37763
rect 57153 37691 57246 37729
rect 57153 37657 57182 37691
rect 57216 37657 57246 37691
rect 57153 37619 57246 37657
rect 57153 37585 57182 37619
rect 57216 37585 57246 37619
rect 57153 37547 57246 37585
rect 57153 37513 57182 37547
rect 57216 37513 57246 37547
rect 57153 37475 57246 37513
rect 57153 37441 57182 37475
rect 57216 37441 57246 37475
rect 57153 37403 57246 37441
rect 57153 37369 57182 37403
rect 57216 37369 57246 37403
rect 57153 37331 57246 37369
rect 57153 37297 57182 37331
rect 57216 37297 57246 37331
rect 57153 37259 57246 37297
rect 57153 37225 57182 37259
rect 57216 37225 57246 37259
rect 57153 37187 57246 37225
rect 57153 37153 57182 37187
rect 57216 37153 57246 37187
rect 57153 37115 57246 37153
rect 57153 37081 57182 37115
rect 57216 37081 57246 37115
rect 57153 37043 57246 37081
rect 57153 37009 57182 37043
rect 57216 37009 57246 37043
rect 68368 37942 68461 37975
rect 68368 37908 68397 37942
rect 68431 37908 68461 37942
rect 68368 37870 68461 37908
rect 68368 37836 68397 37870
rect 68431 37836 68461 37870
rect 68368 37798 68461 37836
rect 68368 37764 68397 37798
rect 68431 37764 68461 37798
rect 68368 37726 68461 37764
rect 68368 37692 68397 37726
rect 68431 37692 68461 37726
rect 68368 37654 68461 37692
rect 68368 37620 68397 37654
rect 68431 37620 68461 37654
rect 68368 37582 68461 37620
rect 68368 37548 68397 37582
rect 68431 37548 68461 37582
rect 68368 37510 68461 37548
rect 68368 37476 68397 37510
rect 68431 37476 68461 37510
rect 68368 37438 68461 37476
rect 68368 37404 68397 37438
rect 68431 37404 68461 37438
rect 68368 37366 68461 37404
rect 68368 37332 68397 37366
rect 68431 37332 68461 37366
rect 68368 37294 68461 37332
rect 68368 37260 68397 37294
rect 68431 37260 68461 37294
rect 68368 37222 68461 37260
rect 68368 37188 68397 37222
rect 68431 37188 68461 37222
rect 68368 37150 68461 37188
rect 68368 37116 68397 37150
rect 68431 37116 68461 37150
rect 68368 37078 68461 37116
rect 68368 37044 68397 37078
rect 68431 37044 68461 37078
rect 68368 37011 68461 37044
rect 57153 36971 57246 37009
rect 57153 36937 57182 36971
rect 57216 36937 57246 36971
rect 57153 36899 57246 36937
rect 57153 36865 57182 36899
rect 57216 36865 57246 36899
rect 57153 36827 57246 36865
rect 57153 36793 57182 36827
rect 57216 36793 57246 36827
rect 57153 36755 57246 36793
rect 57153 36721 57182 36755
rect 57216 36721 57246 36755
rect 57153 36683 57246 36721
rect 57153 36649 57182 36683
rect 57216 36649 57246 36683
rect 57153 36611 57246 36649
rect 57153 36577 57182 36611
rect 57216 36577 57246 36611
rect 57153 36539 57246 36577
rect 57153 36505 57182 36539
rect 57216 36505 57246 36539
rect 57153 36467 57246 36505
rect 57153 36433 57182 36467
rect 57216 36433 57246 36467
rect 57153 36395 57246 36433
rect 57153 36361 57182 36395
rect 57216 36361 57246 36395
rect 57153 36323 57246 36361
rect 57153 36289 57182 36323
rect 57216 36289 57246 36323
rect 57153 36251 57246 36289
rect 57153 36217 57182 36251
rect 57216 36217 57246 36251
rect 57153 36179 57246 36217
rect 57153 36145 57182 36179
rect 57216 36145 57246 36179
rect 57153 36107 57246 36145
rect 57153 36073 57182 36107
rect 57216 36073 57246 36107
rect 57153 36035 57246 36073
rect 57153 36001 57182 36035
rect 57216 36001 57246 36035
rect 57153 35963 57246 36001
rect 57153 35929 57182 35963
rect 57216 35929 57246 35963
rect 57153 35891 57246 35929
rect 57153 35857 57182 35891
rect 57216 35857 57246 35891
rect 57153 35819 57246 35857
rect 57153 35785 57182 35819
rect 57216 35785 57246 35819
rect 57153 35747 57246 35785
rect 57153 35713 57182 35747
rect 57216 35713 57246 35747
rect 57153 35675 57246 35713
rect 57153 35641 57182 35675
rect 57216 35641 57246 35675
rect 57153 35603 57246 35641
rect 57153 35569 57182 35603
rect 57216 35569 57246 35603
rect 57153 35531 57246 35569
rect 57153 35497 57182 35531
rect 57216 35497 57246 35531
rect 57153 35459 57246 35497
rect 57153 35425 57182 35459
rect 57216 35425 57246 35459
rect 57153 35387 57246 35425
rect 57153 35353 57182 35387
rect 57216 35353 57246 35387
rect 57153 35315 57246 35353
rect 68368 36113 68461 36127
rect 68368 36079 68397 36113
rect 68431 36079 68461 36113
rect 68368 36041 68461 36079
rect 68368 36007 68397 36041
rect 68431 36007 68461 36041
rect 68368 35969 68461 36007
rect 68368 35935 68397 35969
rect 68431 35935 68461 35969
rect 68368 35897 68461 35935
rect 68368 35863 68397 35897
rect 68431 35863 68461 35897
rect 68368 35825 68461 35863
rect 68368 35791 68397 35825
rect 68431 35791 68461 35825
rect 68368 35753 68461 35791
rect 68368 35719 68397 35753
rect 68431 35719 68461 35753
rect 68368 35681 68461 35719
rect 68368 35647 68397 35681
rect 68431 35647 68461 35681
rect 68368 35609 68461 35647
rect 68368 35575 68397 35609
rect 68431 35575 68461 35609
rect 68368 35537 68461 35575
rect 68368 35503 68397 35537
rect 68431 35503 68461 35537
rect 68368 35465 68461 35503
rect 68368 35431 68397 35465
rect 68431 35431 68461 35465
rect 68368 35393 68461 35431
rect 68368 35359 68397 35393
rect 68431 35359 68461 35393
rect 68368 35345 68461 35359
rect 57153 35281 57182 35315
rect 57216 35281 57246 35315
rect 57153 35243 57246 35281
rect 57153 35209 57182 35243
rect 57216 35209 57246 35243
rect 57153 35171 57246 35209
rect 57153 35137 57182 35171
rect 57216 35137 57246 35171
rect 57153 35099 57246 35137
rect 57153 35065 57182 35099
rect 57216 35065 57246 35099
rect 57153 35027 57246 35065
rect 57153 34993 57182 35027
rect 57216 34993 57246 35027
rect 57153 34955 57246 34993
rect 57153 34921 57182 34955
rect 57216 34921 57246 34955
rect 57153 34883 57246 34921
rect 57153 34849 57182 34883
rect 57216 34849 57246 34883
rect 57153 34811 57246 34849
rect 57153 34777 57182 34811
rect 57216 34777 57246 34811
rect 57153 34739 57246 34777
rect 57153 34705 57182 34739
rect 57216 34705 57246 34739
rect 57153 34688 57246 34705
rect 63647 34494 68184 34524
rect 63647 34460 63666 34494
rect 63700 34460 63738 34494
rect 63772 34460 63810 34494
rect 63844 34460 63882 34494
rect 63916 34460 63954 34494
rect 63988 34460 64026 34494
rect 64060 34460 64098 34494
rect 64132 34460 64170 34494
rect 64204 34460 64242 34494
rect 64276 34460 64314 34494
rect 64348 34460 64386 34494
rect 64420 34460 64458 34494
rect 64492 34460 64530 34494
rect 64564 34460 64602 34494
rect 64636 34460 64674 34494
rect 64708 34460 64746 34494
rect 64780 34460 64818 34494
rect 64852 34460 64890 34494
rect 64924 34460 64962 34494
rect 64996 34460 65034 34494
rect 65068 34460 65106 34494
rect 65140 34460 65178 34494
rect 65212 34460 65250 34494
rect 65284 34460 65322 34494
rect 65356 34460 65394 34494
rect 65428 34460 65466 34494
rect 65500 34460 65538 34494
rect 65572 34460 65610 34494
rect 65644 34460 65682 34494
rect 65716 34460 65754 34494
rect 65788 34460 65826 34494
rect 65860 34460 65898 34494
rect 65932 34460 65970 34494
rect 66004 34460 66042 34494
rect 66076 34460 66114 34494
rect 66148 34460 66186 34494
rect 66220 34460 66258 34494
rect 66292 34460 66330 34494
rect 66364 34460 66402 34494
rect 66436 34460 66474 34494
rect 66508 34460 66546 34494
rect 66580 34460 66618 34494
rect 66652 34460 66690 34494
rect 66724 34460 66762 34494
rect 66796 34460 66834 34494
rect 66868 34460 66906 34494
rect 66940 34460 66978 34494
rect 67012 34460 67050 34494
rect 67084 34460 67122 34494
rect 67156 34460 67194 34494
rect 67228 34460 67266 34494
rect 67300 34460 67338 34494
rect 67372 34460 67410 34494
rect 67444 34460 67482 34494
rect 67516 34460 67554 34494
rect 67588 34460 67626 34494
rect 67660 34460 67698 34494
rect 67732 34460 67770 34494
rect 67804 34460 67842 34494
rect 67876 34460 67914 34494
rect 67948 34460 67986 34494
rect 68020 34460 68058 34494
rect 68092 34460 68130 34494
rect 68164 34460 68184 34494
rect 63647 34431 68184 34460
<< viali >>
rect 68283 100652 68317 100686
rect 68283 100580 68317 100614
rect 68283 100508 68317 100542
rect 68283 100436 68317 100470
rect 68283 100364 68317 100398
rect 68283 100292 68317 100326
rect 68283 100220 68317 100254
rect 68283 100148 68317 100182
rect 68283 100076 68317 100110
rect 68283 100004 68317 100038
rect 68283 99932 68317 99966
rect 68283 99860 68317 99894
rect 68283 99788 68317 99822
rect 68283 99716 68317 99750
rect 68283 99644 68317 99678
rect 68283 99572 68317 99606
rect 68283 99500 68317 99534
rect 68283 99428 68317 99462
rect 68283 99356 68317 99390
rect 68283 99284 68317 99318
rect 68283 99212 68317 99246
rect 68283 99140 68317 99174
rect 68283 99068 68317 99102
rect 68283 98996 68317 99030
rect 68283 98924 68317 98958
rect 68283 98852 68317 98886
rect 68283 98780 68317 98814
rect 68283 98708 68317 98742
rect 68283 98636 68317 98670
rect 68283 98564 68317 98598
rect 68283 98492 68317 98526
rect 68283 98420 68317 98454
rect 68283 98348 68317 98382
rect 68283 98276 68317 98310
rect 68283 98204 68317 98238
rect 68283 98132 68317 98166
rect 68283 98060 68317 98094
rect 68283 97988 68317 98022
rect 68283 97916 68317 97950
rect 68283 97844 68317 97878
rect 68283 97772 68317 97806
rect 68283 97700 68317 97734
rect 68283 97628 68317 97662
rect 68283 97556 68317 97590
rect 68283 97484 68317 97518
rect 57504 84734 57538 84768
rect 57504 84662 57538 84696
rect 57504 84590 57538 84624
rect 57504 84518 57538 84552
rect 57504 84446 57538 84480
rect 57504 84374 57538 84408
rect 57504 84302 57538 84336
rect 57504 84230 57538 84264
rect 57504 84158 57538 84192
rect 57504 84086 57538 84120
rect 57504 84014 57538 84048
rect 57504 83942 57538 83976
rect 57504 83870 57538 83904
rect 57504 83798 57538 83832
rect 57504 83726 57538 83760
rect 57504 83654 57538 83688
rect 57504 83582 57538 83616
rect 57504 83510 57538 83544
rect 57504 83438 57538 83472
rect 57504 83366 57538 83400
rect 57504 83294 57538 83328
rect 57504 83222 57538 83256
rect 57504 83150 57538 83184
rect 57504 83078 57538 83112
rect 57504 83006 57538 83040
rect 57504 82934 57538 82968
rect 57504 82862 57538 82896
rect 57504 82790 57538 82824
rect 57504 82718 57538 82752
rect 57504 82646 57538 82680
rect 57504 82574 57538 82608
rect 57504 82502 57538 82536
rect 57504 82430 57538 82464
rect 57504 82358 57538 82392
rect 57504 82286 57538 82320
rect 57504 82214 57538 82248
rect 57504 82142 57538 82176
rect 57504 82070 57538 82104
rect 57504 81998 57538 82032
rect 57504 81926 57538 81960
rect 57504 81854 57538 81888
rect 57504 81782 57538 81816
rect 57504 81710 57538 81744
rect 57504 81638 57538 81672
rect 57504 81566 57538 81600
rect 57504 81494 57538 81528
rect 57504 81422 57538 81456
rect 57504 81350 57538 81384
rect 57504 81278 57538 81312
rect 57504 81206 57538 81240
rect 57504 81134 57538 81168
rect 57504 81062 57538 81096
rect 57504 80990 57538 81024
rect 57504 80918 57538 80952
rect 57504 80846 57538 80880
rect 57504 80774 57538 80808
rect 57504 80702 57538 80736
rect 57504 80630 57538 80664
rect 57504 80558 57538 80592
rect 57504 80486 57538 80520
rect 57504 80414 57538 80448
rect 57504 80342 57538 80376
rect 57504 80270 57538 80304
rect 57504 80198 57538 80232
rect 57504 80126 57538 80160
rect 57504 80054 57538 80088
rect 57504 79982 57538 80016
rect 57504 79910 57538 79944
rect 57504 79838 57538 79872
rect 57504 79766 57538 79800
rect 57504 79694 57538 79728
rect 57504 79622 57538 79656
rect 57504 79550 57538 79584
rect 57504 79478 57538 79512
rect 57504 79406 57538 79440
rect 57504 79334 57538 79368
rect 57504 79262 57538 79296
rect 57504 79190 57538 79224
rect 57504 79118 57538 79152
rect 57504 79046 57538 79080
rect 57504 78974 57538 79008
rect 57504 78902 57538 78936
rect 57504 78830 57538 78864
rect 57504 78758 57538 78792
rect 57504 78686 57538 78720
rect 57504 78614 57538 78648
rect 57504 78542 57538 78576
rect 57504 78470 57538 78504
rect 57504 78398 57538 78432
rect 57504 78326 57538 78360
rect 57504 78254 57538 78288
rect 57504 78182 57538 78216
rect 57504 78110 57538 78144
rect 57504 78038 57538 78072
rect 57504 77966 57538 78000
rect 57504 77894 57538 77928
rect 57504 77822 57538 77856
rect 57504 77750 57538 77784
rect 57504 77678 57538 77712
rect 57504 77606 57538 77640
rect 57504 77534 57538 77568
rect 57504 77462 57538 77496
rect 57504 77390 57538 77424
rect 57504 77318 57538 77352
rect 57504 77246 57538 77280
rect 57504 77174 57538 77208
rect 51487 74976 51521 75010
rect 51559 74976 51593 75010
rect 51631 74976 51665 75010
rect 51703 74976 51737 75010
rect 51775 74976 51809 75010
rect 51847 74976 51881 75010
rect 51919 74976 51953 75010
rect 51991 74976 52025 75010
rect 52063 74976 52097 75010
rect 52135 74976 52169 75010
rect 52207 74976 52241 75010
rect 52279 74976 52313 75010
rect 52351 74976 52385 75010
rect 52423 74976 52457 75010
rect 52495 74976 52529 75010
rect 52567 74976 52601 75010
rect 52639 74976 52673 75010
rect 52711 74976 52745 75010
rect 52783 74976 52817 75010
rect 52855 74976 52889 75010
rect 52927 74976 52961 75010
rect 52999 74976 53033 75010
rect 53071 74976 53105 75010
rect 53143 74976 53177 75010
rect 53215 74976 53249 75010
rect 53287 74976 53321 75010
rect 53359 74976 53393 75010
rect 53431 74976 53465 75010
rect 53503 74976 53537 75010
rect 53575 74976 53609 75010
rect 53647 74976 53681 75010
rect 53719 74976 53753 75010
rect 53791 74976 53825 75010
rect 53863 74976 53897 75010
rect 53935 74976 53969 75010
rect 54007 74976 54041 75010
rect 54079 74976 54113 75010
rect 54151 74976 54185 75010
rect 54223 74976 54257 75010
rect 54295 74976 54329 75010
rect 54367 74976 54401 75010
rect 54439 74976 54473 75010
rect 54511 74976 54545 75010
rect 54583 74976 54617 75010
rect 54655 74976 54689 75010
rect 54727 74976 54761 75010
rect 54799 74976 54833 75010
rect 54871 74976 54905 75010
rect 54943 74976 54977 75010
rect 55015 74976 55049 75010
rect 55087 74976 55121 75010
rect 55159 74976 55193 75010
rect 55231 74976 55265 75010
rect 55303 74976 55337 75010
rect 55375 74976 55409 75010
rect 55447 74976 55481 75010
rect 55519 74976 55553 75010
rect 55591 74976 55625 75010
rect 55663 74976 55697 75010
rect 55735 74976 55769 75010
rect 55807 74976 55841 75010
rect 55879 74976 55913 75010
rect 55951 74976 55985 75010
rect 56023 74976 56057 75010
rect 56095 74976 56129 75010
rect 56167 74976 56201 75010
rect 56239 74976 56273 75010
rect 56311 74976 56345 75010
rect 56383 74976 56417 75010
rect 56455 74976 56489 75010
rect 56527 74976 56561 75010
rect 56599 74976 56633 75010
rect 56671 74976 56705 75010
rect 56743 74976 56777 75010
rect 56815 74976 56849 75010
rect 56887 74976 56921 75010
rect 57119 74701 57153 74735
rect 57119 74629 57153 74663
rect 57119 74557 57153 74591
rect 57119 74485 57153 74519
rect 57119 74413 57153 74447
rect 57119 74341 57153 74375
rect 57119 74269 57153 74303
rect 57119 74197 57153 74231
rect 57119 74125 57153 74159
rect 57119 74053 57153 74087
rect 57119 73981 57153 74015
rect 57119 73909 57153 73943
rect 57119 73837 57153 73871
rect 57119 73765 57153 73799
rect 57119 73693 57153 73727
rect 57119 73621 57153 73655
rect 57119 73549 57153 73583
rect 57119 73477 57153 73511
rect 31047 73435 31081 73469
rect 30717 73386 30751 73420
rect 30789 73386 30823 73420
rect 30861 73386 30895 73420
rect 57119 73405 57153 73439
rect 31047 73349 31081 73383
rect 57119 73333 57153 73367
rect 57119 73261 57153 73295
rect 57119 73189 57153 73223
rect 57119 73117 57153 73151
rect 57119 73045 57153 73079
rect 57119 72973 57153 73007
rect 57119 72901 57153 72935
rect 57119 72829 57153 72863
rect 57119 72757 57153 72791
rect 57119 72685 57153 72719
rect 57119 72613 57153 72647
rect 57119 72541 57153 72575
rect 57119 72469 57153 72503
rect 57119 72397 57153 72431
rect 57119 72325 57153 72359
rect 57119 72253 57153 72287
rect 57119 72181 57153 72215
rect 57119 72109 57153 72143
rect 57119 72037 57153 72071
rect 57119 71965 57153 71999
rect 57119 71893 57153 71927
rect 57119 71821 57153 71855
rect 57504 69773 57538 69807
rect 57504 69701 57538 69735
rect 57504 69629 57538 69663
rect 57504 69557 57538 69591
rect 57504 69485 57538 69519
rect 57504 69413 57538 69447
rect 57504 69341 57538 69375
rect 57504 69269 57538 69303
rect 57504 69197 57538 69231
rect 57504 69125 57538 69159
rect 57504 69053 57538 69087
rect 57504 68981 57538 69015
rect 57504 68909 57538 68943
rect 57504 68837 57538 68871
rect 98902 68915 98936 68949
rect 98902 68843 98936 68877
rect 97078 68805 97112 68839
rect 97697 68804 97731 68838
rect 57504 68765 57538 68799
rect 98099 68798 98133 68832
rect 98255 68804 98289 68838
rect 57504 68693 57538 68727
rect 97222 68724 97256 68758
rect 97999 68739 98033 68773
rect 98902 68771 98936 68805
rect 100375 68824 100409 68858
rect 100547 68824 100581 68858
rect 100719 68824 100753 68858
rect 100891 68824 100925 68858
rect 101063 68824 101097 68858
rect 101268 68824 101302 68858
rect 101445 68824 101479 68858
rect 101617 68824 101651 68858
rect 101789 68824 101823 68858
rect 101961 68824 101995 68858
rect 102133 68824 102167 68858
rect 102305 68824 102339 68858
rect 100097 68774 100131 68808
rect 99633 68735 99667 68769
rect 99705 68735 99739 68769
rect 99777 68735 99811 68769
rect 99849 68735 99883 68769
rect 99921 68735 99955 68769
rect 99993 68735 100027 68769
rect 100371 68738 100405 68772
rect 100443 68738 100477 68772
rect 57504 68621 57538 68655
rect 98902 68699 98936 68733
rect 100097 68702 100131 68736
rect 98902 68627 98936 68661
rect 57504 68549 57538 68583
rect 57504 68477 57538 68511
rect 57504 68405 57538 68439
rect 98902 67765 98936 67799
rect 98902 67693 98936 67727
rect 97078 67655 97112 67689
rect 97697 67654 97731 67688
rect 98099 67648 98133 67682
rect 98255 67654 98289 67688
rect 97222 67574 97256 67608
rect 97999 67589 98033 67623
rect 98902 67621 98936 67655
rect 100375 67674 100409 67708
rect 100547 67674 100581 67708
rect 100719 67674 100753 67708
rect 100891 67674 100925 67708
rect 101063 67674 101097 67708
rect 101268 67674 101302 67708
rect 101445 67674 101479 67708
rect 101617 67674 101651 67708
rect 101789 67674 101823 67708
rect 101961 67674 101995 67708
rect 102133 67674 102167 67708
rect 102305 67674 102339 67708
rect 100097 67624 100131 67658
rect 99633 67585 99667 67619
rect 99705 67585 99739 67619
rect 99777 67585 99811 67619
rect 99849 67585 99883 67619
rect 99921 67585 99955 67619
rect 99993 67585 100027 67619
rect 100371 67588 100405 67622
rect 100443 67588 100477 67622
rect 98902 67549 98936 67583
rect 100097 67552 100131 67586
rect 98902 67477 98936 67511
rect 57504 65314 57538 65348
rect 57504 65242 57538 65276
rect 57504 65170 57538 65204
rect 98902 65225 98936 65259
rect 98902 65153 98936 65187
rect 57504 65098 57538 65132
rect 97078 65115 97112 65149
rect 97697 65114 97731 65148
rect 98099 65108 98133 65142
rect 98255 65114 98289 65148
rect 57504 65026 57538 65060
rect 97222 65034 97256 65068
rect 97999 65049 98033 65083
rect 98902 65081 98936 65115
rect 100375 65134 100409 65168
rect 100547 65134 100581 65168
rect 100719 65134 100753 65168
rect 100891 65134 100925 65168
rect 101063 65134 101097 65168
rect 101268 65134 101302 65168
rect 101445 65134 101479 65168
rect 101617 65134 101651 65168
rect 101789 65134 101823 65168
rect 101961 65134 101995 65168
rect 102133 65134 102167 65168
rect 102305 65134 102339 65168
rect 100097 65084 100131 65118
rect 99633 65045 99667 65079
rect 99705 65045 99739 65079
rect 99777 65045 99811 65079
rect 99849 65045 99883 65079
rect 99921 65045 99955 65079
rect 99993 65045 100027 65079
rect 100371 65048 100405 65082
rect 100443 65048 100477 65082
rect 57504 64954 57538 64988
rect 98902 65009 98936 65043
rect 100097 65012 100131 65046
rect 98902 64937 98936 64971
rect 57504 64882 57538 64916
rect 57504 64810 57538 64844
rect 57504 64738 57538 64772
rect 57504 64666 57538 64700
rect 57504 64594 57538 64628
rect 57504 64522 57538 64556
rect 57504 64450 57538 64484
rect 57504 64378 57538 64412
rect 57504 64306 57538 64340
rect 57504 64234 57538 64268
rect 57504 64162 57538 64196
rect 57504 64090 57538 64124
rect 98902 63955 98936 63989
rect 98902 63883 98936 63917
rect 97078 63845 97112 63879
rect 97697 63844 97731 63878
rect 98099 63838 98133 63872
rect 98255 63844 98289 63878
rect 51474 63761 51508 63795
rect 51546 63761 51580 63795
rect 51618 63761 51652 63795
rect 51690 63761 51724 63795
rect 51762 63761 51796 63795
rect 51834 63761 51868 63795
rect 51906 63761 51940 63795
rect 51978 63761 52012 63795
rect 52050 63761 52084 63795
rect 52122 63761 52156 63795
rect 52194 63761 52228 63795
rect 52266 63761 52300 63795
rect 52338 63761 52372 63795
rect 52410 63761 52444 63795
rect 52482 63761 52516 63795
rect 52554 63761 52588 63795
rect 52626 63761 52660 63795
rect 52698 63761 52732 63795
rect 52770 63761 52804 63795
rect 52842 63761 52876 63795
rect 52914 63761 52948 63795
rect 52986 63761 53020 63795
rect 53058 63761 53092 63795
rect 53130 63761 53164 63795
rect 53202 63761 53236 63795
rect 53274 63761 53308 63795
rect 53346 63761 53380 63795
rect 53418 63761 53452 63795
rect 53490 63761 53524 63795
rect 53562 63761 53596 63795
rect 53634 63761 53668 63795
rect 53706 63761 53740 63795
rect 53778 63761 53812 63795
rect 53850 63761 53884 63795
rect 53922 63761 53956 63795
rect 53994 63761 54028 63795
rect 54066 63761 54100 63795
rect 54138 63761 54172 63795
rect 54210 63761 54244 63795
rect 54282 63761 54316 63795
rect 54354 63761 54388 63795
rect 54426 63761 54460 63795
rect 54498 63761 54532 63795
rect 54570 63761 54604 63795
rect 54642 63761 54676 63795
rect 54714 63761 54748 63795
rect 54786 63761 54820 63795
rect 54858 63761 54892 63795
rect 54930 63761 54964 63795
rect 55002 63761 55036 63795
rect 55074 63761 55108 63795
rect 55146 63761 55180 63795
rect 55218 63761 55252 63795
rect 55290 63761 55324 63795
rect 55362 63761 55396 63795
rect 55434 63761 55468 63795
rect 55506 63761 55540 63795
rect 55578 63761 55612 63795
rect 55650 63761 55684 63795
rect 55722 63761 55756 63795
rect 55794 63761 55828 63795
rect 55866 63761 55900 63795
rect 55938 63761 55972 63795
rect 56010 63761 56044 63795
rect 56082 63761 56116 63795
rect 56154 63761 56188 63795
rect 56226 63761 56260 63795
rect 56298 63761 56332 63795
rect 56370 63761 56404 63795
rect 56442 63761 56476 63795
rect 56514 63761 56548 63795
rect 56586 63761 56620 63795
rect 56658 63761 56692 63795
rect 56730 63761 56764 63795
rect 56802 63761 56836 63795
rect 56874 63761 56908 63795
rect 97222 63764 97256 63798
rect 97999 63779 98033 63813
rect 98902 63811 98936 63845
rect 100375 63864 100409 63898
rect 100547 63864 100581 63898
rect 100719 63864 100753 63898
rect 100891 63864 100925 63898
rect 101063 63864 101097 63898
rect 101268 63864 101302 63898
rect 101445 63864 101479 63898
rect 101617 63864 101651 63898
rect 101789 63864 101823 63898
rect 101961 63864 101995 63898
rect 102133 63864 102167 63898
rect 102305 63864 102339 63898
rect 100097 63814 100131 63848
rect 99633 63775 99667 63809
rect 99705 63775 99739 63809
rect 99777 63775 99811 63809
rect 99849 63775 99883 63809
rect 99921 63775 99955 63809
rect 99993 63775 100027 63809
rect 100371 63778 100405 63812
rect 100443 63778 100477 63812
rect 98902 63739 98936 63773
rect 100097 63742 100131 63776
rect 98902 63667 98936 63701
rect 25299 63102 25333 63136
rect 25299 63030 25333 63064
rect 25299 62958 25333 62992
rect 25299 62886 25333 62920
rect 25299 62538 25333 62572
rect 25299 62466 25333 62500
rect 25299 62394 25333 62428
rect 25299 62322 25333 62356
rect 25299 62250 25333 62284
rect 57182 40105 57216 40139
rect 57182 40033 57216 40067
rect 57182 39961 57216 39995
rect 57182 39889 57216 39923
rect 57182 39817 57216 39851
rect 57182 39745 57216 39779
rect 57182 39673 57216 39707
rect 57182 39601 57216 39635
rect 57182 39529 57216 39563
rect 57182 39457 57216 39491
rect 57182 39385 57216 39419
rect 57182 39313 57216 39347
rect 57182 39241 57216 39275
rect 57182 39169 57216 39203
rect 57182 39097 57216 39131
rect 57182 39025 57216 39059
rect 57182 38953 57216 38987
rect 57182 38881 57216 38915
rect 57182 38809 57216 38843
rect 57182 38737 57216 38771
rect 57182 38665 57216 38699
rect 57182 38593 57216 38627
rect 57182 38521 57216 38555
rect 57182 38449 57216 38483
rect 68397 40110 68431 40144
rect 68397 40038 68431 40072
rect 68397 39966 68431 40000
rect 68397 39894 68431 39928
rect 68397 39822 68431 39856
rect 68397 39750 68431 39784
rect 68397 39678 68431 39712
rect 68397 39606 68431 39640
rect 68397 39534 68431 39568
rect 68397 39462 68431 39496
rect 68397 39390 68431 39424
rect 68397 39318 68431 39352
rect 68397 39246 68431 39280
rect 68397 39174 68431 39208
rect 68397 39102 68431 39136
rect 68397 39030 68431 39064
rect 68397 38958 68431 38992
rect 68397 38886 68431 38920
rect 68397 38814 68431 38848
rect 68397 38742 68431 38776
rect 68397 38670 68431 38704
rect 68397 38598 68431 38632
rect 68397 38526 68431 38560
rect 68397 38454 68431 38488
rect 57182 38377 57216 38411
rect 57182 38305 57216 38339
rect 57182 38233 57216 38267
rect 57182 38161 57216 38195
rect 57182 38089 57216 38123
rect 57182 38017 57216 38051
rect 57182 37945 57216 37979
rect 57182 37873 57216 37907
rect 57182 37801 57216 37835
rect 57182 37729 57216 37763
rect 57182 37657 57216 37691
rect 57182 37585 57216 37619
rect 57182 37513 57216 37547
rect 57182 37441 57216 37475
rect 57182 37369 57216 37403
rect 57182 37297 57216 37331
rect 57182 37225 57216 37259
rect 57182 37153 57216 37187
rect 57182 37081 57216 37115
rect 57182 37009 57216 37043
rect 68397 37908 68431 37942
rect 68397 37836 68431 37870
rect 68397 37764 68431 37798
rect 68397 37692 68431 37726
rect 68397 37620 68431 37654
rect 68397 37548 68431 37582
rect 68397 37476 68431 37510
rect 68397 37404 68431 37438
rect 68397 37332 68431 37366
rect 68397 37260 68431 37294
rect 68397 37188 68431 37222
rect 68397 37116 68431 37150
rect 68397 37044 68431 37078
rect 57182 36937 57216 36971
rect 57182 36865 57216 36899
rect 57182 36793 57216 36827
rect 57182 36721 57216 36755
rect 57182 36649 57216 36683
rect 57182 36577 57216 36611
rect 57182 36505 57216 36539
rect 57182 36433 57216 36467
rect 57182 36361 57216 36395
rect 57182 36289 57216 36323
rect 57182 36217 57216 36251
rect 57182 36145 57216 36179
rect 57182 36073 57216 36107
rect 57182 36001 57216 36035
rect 57182 35929 57216 35963
rect 57182 35857 57216 35891
rect 57182 35785 57216 35819
rect 57182 35713 57216 35747
rect 57182 35641 57216 35675
rect 57182 35569 57216 35603
rect 57182 35497 57216 35531
rect 57182 35425 57216 35459
rect 57182 35353 57216 35387
rect 68397 36079 68431 36113
rect 68397 36007 68431 36041
rect 68397 35935 68431 35969
rect 68397 35863 68431 35897
rect 68397 35791 68431 35825
rect 68397 35719 68431 35753
rect 68397 35647 68431 35681
rect 68397 35575 68431 35609
rect 68397 35503 68431 35537
rect 68397 35431 68431 35465
rect 68397 35359 68431 35393
rect 57182 35281 57216 35315
rect 57182 35209 57216 35243
rect 57182 35137 57216 35171
rect 57182 35065 57216 35099
rect 57182 34993 57216 35027
rect 57182 34921 57216 34955
rect 57182 34849 57216 34883
rect 57182 34777 57216 34811
rect 57182 34705 57216 34739
rect 63666 34460 63700 34494
rect 63738 34460 63772 34494
rect 63810 34460 63844 34494
rect 63882 34460 63916 34494
rect 63954 34460 63988 34494
rect 64026 34460 64060 34494
rect 64098 34460 64132 34494
rect 64170 34460 64204 34494
rect 64242 34460 64276 34494
rect 64314 34460 64348 34494
rect 64386 34460 64420 34494
rect 64458 34460 64492 34494
rect 64530 34460 64564 34494
rect 64602 34460 64636 34494
rect 64674 34460 64708 34494
rect 64746 34460 64780 34494
rect 64818 34460 64852 34494
rect 64890 34460 64924 34494
rect 64962 34460 64996 34494
rect 65034 34460 65068 34494
rect 65106 34460 65140 34494
rect 65178 34460 65212 34494
rect 65250 34460 65284 34494
rect 65322 34460 65356 34494
rect 65394 34460 65428 34494
rect 65466 34460 65500 34494
rect 65538 34460 65572 34494
rect 65610 34460 65644 34494
rect 65682 34460 65716 34494
rect 65754 34460 65788 34494
rect 65826 34460 65860 34494
rect 65898 34460 65932 34494
rect 65970 34460 66004 34494
rect 66042 34460 66076 34494
rect 66114 34460 66148 34494
rect 66186 34460 66220 34494
rect 66258 34460 66292 34494
rect 66330 34460 66364 34494
rect 66402 34460 66436 34494
rect 66474 34460 66508 34494
rect 66546 34460 66580 34494
rect 66618 34460 66652 34494
rect 66690 34460 66724 34494
rect 66762 34460 66796 34494
rect 66834 34460 66868 34494
rect 66906 34460 66940 34494
rect 66978 34460 67012 34494
rect 67050 34460 67084 34494
rect 67122 34460 67156 34494
rect 67194 34460 67228 34494
rect 67266 34460 67300 34494
rect 67338 34460 67372 34494
rect 67410 34460 67444 34494
rect 67482 34460 67516 34494
rect 67554 34460 67588 34494
rect 67626 34460 67660 34494
rect 67698 34460 67732 34494
rect 67770 34460 67804 34494
rect 67842 34460 67876 34494
rect 67914 34460 67948 34494
rect 67986 34460 68020 34494
rect 68058 34460 68092 34494
rect 68130 34460 68164 34494
<< metal1 >>
rect 41674 102134 41930 102162
rect 41674 101954 41712 102134
rect 41892 101954 41930 102134
rect 41674 101926 41930 101954
rect 69690 102105 69946 102133
rect 40235 100740 40356 100745
rect 40235 100688 40269 100740
rect 40321 100688 40356 100740
rect 40235 100676 40356 100688
rect 40235 100624 40269 100676
rect 40321 100624 40356 100676
rect 40235 100612 40356 100624
rect 40235 100560 40269 100612
rect 40321 100560 40356 100612
rect 40235 100548 40356 100560
rect 40235 100496 40269 100548
rect 40321 100496 40356 100548
rect 40235 100484 40356 100496
rect 40235 100432 40269 100484
rect 40321 100432 40356 100484
rect 40235 100420 40356 100432
rect 40235 100368 40269 100420
rect 40321 100368 40356 100420
rect 40235 100356 40356 100368
rect 40235 100304 40269 100356
rect 40321 100304 40356 100356
rect 40235 100292 40356 100304
rect 40235 100240 40269 100292
rect 40321 100240 40356 100292
rect 40235 100228 40356 100240
rect 40235 100176 40269 100228
rect 40321 100176 40356 100228
rect 40235 100164 40356 100176
rect 40235 100112 40269 100164
rect 40321 100112 40356 100164
rect 40235 100100 40356 100112
rect 40235 100048 40269 100100
rect 40321 100048 40356 100100
rect 40235 100036 40356 100048
rect 40235 99984 40269 100036
rect 40321 99984 40356 100036
rect 40235 99972 40356 99984
rect 40235 99920 40269 99972
rect 40321 99920 40356 99972
rect 40235 99908 40356 99920
rect 40235 99856 40269 99908
rect 40321 99856 40356 99908
rect 40235 99844 40356 99856
rect 40235 99792 40269 99844
rect 40321 99792 40356 99844
rect 40235 99780 40356 99792
rect 40235 99728 40269 99780
rect 40321 99728 40356 99780
rect 40235 99716 40356 99728
rect 40235 99664 40269 99716
rect 40321 99664 40356 99716
rect 40235 99652 40356 99664
rect 40235 99600 40269 99652
rect 40321 99600 40356 99652
rect 40235 99588 40356 99600
rect 40235 99536 40269 99588
rect 40321 99536 40356 99588
rect 40235 99524 40356 99536
rect 40235 99472 40269 99524
rect 40321 99472 40356 99524
rect 40235 99460 40356 99472
rect 40235 99408 40269 99460
rect 40321 99408 40356 99460
rect 40235 99396 40356 99408
rect 40235 99344 40269 99396
rect 40321 99344 40356 99396
rect 40235 99332 40356 99344
rect 40235 99280 40269 99332
rect 40321 99280 40356 99332
rect 40235 99268 40356 99280
rect 41741 99277 41869 101926
rect 69690 101925 69728 102105
rect 69908 101925 69946 102105
rect 69690 101897 69946 101925
rect 81740 102106 81996 102134
rect 81740 101926 81778 102106
rect 81958 101926 81996 102106
rect 81740 101898 81996 101926
rect 68271 100754 68461 100828
rect 43236 100746 43357 100751
rect 43236 100694 43270 100746
rect 43322 100694 43357 100746
rect 43236 100682 43357 100694
rect 43236 100630 43270 100682
rect 43322 100630 43357 100682
rect 43236 100618 43357 100630
rect 43236 100566 43270 100618
rect 43322 100566 43357 100618
rect 43236 100554 43357 100566
rect 43236 100502 43270 100554
rect 43322 100502 43357 100554
rect 43236 100490 43357 100502
rect 43236 100438 43270 100490
rect 43322 100438 43357 100490
rect 43236 100426 43357 100438
rect 43236 100374 43270 100426
rect 43322 100374 43357 100426
rect 43236 100362 43357 100374
rect 43236 100310 43270 100362
rect 43322 100310 43357 100362
rect 43236 100298 43357 100310
rect 43236 100246 43270 100298
rect 43322 100246 43357 100298
rect 43236 100234 43357 100246
rect 43236 100182 43270 100234
rect 43322 100182 43357 100234
rect 43236 100170 43357 100182
rect 43236 100118 43270 100170
rect 43322 100118 43357 100170
rect 43236 100106 43357 100118
rect 43236 100054 43270 100106
rect 43322 100054 43357 100106
rect 43236 100042 43357 100054
rect 43236 99990 43270 100042
rect 43322 99990 43357 100042
rect 43236 99978 43357 99990
rect 43236 99926 43270 99978
rect 43322 99926 43357 99978
rect 43236 99914 43357 99926
rect 43236 99862 43270 99914
rect 43322 99862 43357 99914
rect 43236 99850 43357 99862
rect 43236 99798 43270 99850
rect 43322 99798 43357 99850
rect 43236 99786 43357 99798
rect 43236 99734 43270 99786
rect 43322 99734 43357 99786
rect 43236 99722 43357 99734
rect 43236 99670 43270 99722
rect 43322 99670 43357 99722
rect 43236 99658 43357 99670
rect 43236 99606 43270 99658
rect 43322 99606 43357 99658
rect 43236 99594 43357 99606
rect 43236 99542 43270 99594
rect 43322 99542 43357 99594
rect 43236 99530 43357 99542
rect 43236 99478 43270 99530
rect 43322 99478 43357 99530
rect 43236 99466 43357 99478
rect 43236 99414 43270 99466
rect 43322 99414 43357 99466
rect 43236 99402 43357 99414
rect 43236 99350 43270 99402
rect 43322 99350 43357 99402
rect 43236 99338 43357 99350
rect 43236 99286 43270 99338
rect 43322 99286 43357 99338
rect 40235 99216 40269 99268
rect 40321 99216 40356 99268
rect 40235 99204 40356 99216
rect 40235 99152 40269 99204
rect 40321 99152 40356 99204
rect 40235 99140 40356 99152
rect 40235 99088 40269 99140
rect 40321 99088 40356 99140
rect 40235 99076 40356 99088
rect 40235 99024 40269 99076
rect 40321 99024 40356 99076
rect 40235 99012 40356 99024
rect 40235 98960 40269 99012
rect 40321 98960 40356 99012
rect 40235 98948 40356 98960
rect 40235 98896 40269 98948
rect 40321 98896 40356 98948
rect 40235 98884 40356 98896
rect 40235 98832 40269 98884
rect 40321 98832 40356 98884
rect 40235 98820 40356 98832
rect 43236 99274 43357 99286
rect 43236 99222 43270 99274
rect 43322 99222 43357 99274
rect 43236 99210 43357 99222
rect 43236 99158 43270 99210
rect 43322 99158 43357 99210
rect 43236 99146 43357 99158
rect 43236 99094 43270 99146
rect 43322 99094 43357 99146
rect 43236 99082 43357 99094
rect 43236 99030 43270 99082
rect 43322 99030 43357 99082
rect 43236 99018 43357 99030
rect 43236 98966 43270 99018
rect 43322 98966 43357 99018
rect 43236 98954 43357 98966
rect 43236 98902 43270 98954
rect 43322 98902 43357 98954
rect 43236 98890 43357 98902
rect 43236 98838 43270 98890
rect 43322 98838 43357 98890
rect 43236 98826 43357 98838
rect 40235 98768 40269 98820
rect 40321 98768 40356 98820
rect 40235 98756 40356 98768
rect 40235 98704 40269 98756
rect 40321 98704 40356 98756
rect 40235 98692 40356 98704
rect 40235 98640 40269 98692
rect 40321 98640 40356 98692
rect 40235 98628 40356 98640
rect 40235 98576 40269 98628
rect 40321 98576 40356 98628
rect 40235 98564 40356 98576
rect 40235 98512 40269 98564
rect 40321 98512 40356 98564
rect 40235 98500 40356 98512
rect 40235 98448 40269 98500
rect 40321 98448 40356 98500
rect 40235 98436 40356 98448
rect 40235 98384 40269 98436
rect 40321 98384 40356 98436
rect 40235 98372 40356 98384
rect 40235 98320 40269 98372
rect 40321 98320 40356 98372
rect 40235 98308 40356 98320
rect 40235 98256 40269 98308
rect 40321 98256 40356 98308
rect 40235 98244 40356 98256
rect 40235 98192 40269 98244
rect 40321 98192 40356 98244
rect 40235 98180 40356 98192
rect 40235 98128 40269 98180
rect 40321 98128 40356 98180
rect 40235 98116 40356 98128
rect 40235 98064 40269 98116
rect 40321 98064 40356 98116
rect 40235 98052 40356 98064
rect 40235 98000 40269 98052
rect 40321 98000 40356 98052
rect 40235 97988 40356 98000
rect 40235 97936 40269 97988
rect 40321 97936 40356 97988
rect 40235 97924 40356 97936
rect 40235 97872 40269 97924
rect 40321 97872 40356 97924
rect 40235 97860 40356 97872
rect 40235 97808 40269 97860
rect 40321 97808 40356 97860
rect 40235 97796 40356 97808
rect 40235 97744 40269 97796
rect 40321 97744 40356 97796
rect 40235 97732 40356 97744
rect 40235 97680 40269 97732
rect 40321 97680 40356 97732
rect 40235 97668 40356 97680
rect 40235 97616 40269 97668
rect 40321 97616 40356 97668
rect 40235 97604 40356 97616
rect 40235 97552 40269 97604
rect 40321 97552 40356 97604
rect 40235 97540 40356 97552
rect 40235 97488 40269 97540
rect 40321 97488 40356 97540
rect 40235 97476 40356 97488
rect 40235 97424 40269 97476
rect 40321 97424 40356 97476
rect 40235 97420 40356 97424
rect 41741 95980 41869 98823
rect 43236 98774 43270 98826
rect 43322 98774 43357 98826
rect 43236 98762 43357 98774
rect 43236 98710 43270 98762
rect 43322 98710 43357 98762
rect 43236 98698 43357 98710
rect 43236 98646 43270 98698
rect 43322 98646 43357 98698
rect 43236 98634 43357 98646
rect 43236 98582 43270 98634
rect 43322 98582 43357 98634
rect 43236 98570 43357 98582
rect 43236 98518 43270 98570
rect 43322 98518 43357 98570
rect 43236 98506 43357 98518
rect 43236 98454 43270 98506
rect 43322 98454 43357 98506
rect 43236 98442 43357 98454
rect 43236 98390 43270 98442
rect 43322 98390 43357 98442
rect 43236 98378 43357 98390
rect 43236 98326 43270 98378
rect 43322 98326 43357 98378
rect 43236 98314 43357 98326
rect 43236 98262 43270 98314
rect 43322 98262 43357 98314
rect 43236 98250 43357 98262
rect 43236 98198 43270 98250
rect 43322 98198 43357 98250
rect 43236 98186 43357 98198
rect 43236 98134 43270 98186
rect 43322 98134 43357 98186
rect 43236 98122 43357 98134
rect 43236 98070 43270 98122
rect 43322 98070 43357 98122
rect 43236 98058 43357 98070
rect 43236 98006 43270 98058
rect 43322 98006 43357 98058
rect 43236 97994 43357 98006
rect 43236 97942 43270 97994
rect 43322 97942 43357 97994
rect 43236 97930 43357 97942
rect 43236 97878 43270 97930
rect 43322 97878 43357 97930
rect 43236 97866 43357 97878
rect 43236 97814 43270 97866
rect 43322 97814 43357 97866
rect 43236 97802 43357 97814
rect 43236 97750 43270 97802
rect 43322 97750 43357 97802
rect 43236 97738 43357 97750
rect 43236 97686 43270 97738
rect 43322 97686 43357 97738
rect 43236 97674 43357 97686
rect 43236 97622 43270 97674
rect 43322 97622 43357 97674
rect 43236 97610 43357 97622
rect 43236 97558 43270 97610
rect 43322 97558 43357 97610
rect 43236 97546 43357 97558
rect 43236 97494 43270 97546
rect 43322 97494 43357 97546
rect 43236 97482 43357 97494
rect 43236 97430 43270 97482
rect 43322 97430 43357 97482
rect 43236 97426 43357 97430
rect 68227 100742 68461 100754
rect 68227 97426 68243 100742
rect 68359 97426 68461 100742
rect 68227 97414 68461 97426
rect 68271 97342 68461 97414
rect 69754 97041 69872 101897
rect 71228 100755 71376 100767
rect 71228 97439 71244 100755
rect 71360 97439 71376 100755
rect 71228 97427 71376 97439
rect 40420 95818 40504 95824
rect 41815 95821 41899 95827
rect 40420 95766 40436 95818
rect 40488 95766 40504 95818
rect 40420 95760 40504 95766
rect 41598 95814 41682 95820
rect 41598 95762 41614 95814
rect 41666 95762 41682 95814
rect 41815 95769 41831 95821
rect 41883 95769 41899 95821
rect 41815 95763 41899 95769
rect 42949 95818 43033 95824
rect 42949 95766 42965 95818
rect 43017 95766 43033 95818
rect 41598 95756 41682 95762
rect 42949 95760 43033 95766
rect 40530 94314 40614 94320
rect 40530 94262 40546 94314
rect 40598 94262 40614 94314
rect 40530 94256 40614 94262
rect 41644 94300 41728 94306
rect 41644 94248 41660 94300
rect 41712 94248 41728 94300
rect 41644 94242 41728 94248
rect 41857 94301 41941 94307
rect 41857 94249 41873 94301
rect 41925 94249 41941 94301
rect 41857 94243 41941 94249
rect 43021 94301 43105 94307
rect 43021 94249 43037 94301
rect 43089 94249 43105 94301
rect 43021 94243 43105 94249
rect 41662 92516 41746 92537
rect 41662 92464 41678 92516
rect 41730 92464 41746 92516
rect 41662 92452 41746 92464
rect 41662 92400 41678 92452
rect 41730 92400 41746 92452
rect 41662 92388 41746 92400
rect 41662 92336 41678 92388
rect 41730 92336 41746 92388
rect 41662 92324 41746 92336
rect 41121 92263 41214 92283
rect 41121 92211 41141 92263
rect 41193 92211 41214 92263
rect 41121 92199 41214 92211
rect 41121 92147 41141 92199
rect 41193 92147 41214 92199
rect 41662 92272 41678 92324
rect 41730 92272 41746 92324
rect 41662 92260 41746 92272
rect 41662 92208 41678 92260
rect 41730 92208 41746 92260
rect 41662 92188 41746 92208
rect 42205 92266 42298 92286
rect 42205 92214 42225 92266
rect 42277 92214 42298 92266
rect 42205 92202 42298 92214
rect 41121 92127 41214 92147
rect 42205 92150 42225 92202
rect 42277 92150 42298 92202
rect 42205 92130 42298 92150
rect 40507 91629 40591 91635
rect 42780 91634 42864 91640
rect 40507 91577 40523 91629
rect 40575 91577 40591 91629
rect 40507 91571 40591 91577
rect 41662 91623 41746 91629
rect 41662 91571 41678 91623
rect 41730 91571 41746 91623
rect 42780 91582 42796 91634
rect 42848 91582 42864 91634
rect 42780 91576 42864 91582
rect 41662 91565 41746 91571
rect 40971 77020 41099 90348
rect 42312 77622 42440 90360
rect 47200 87418 47662 87424
rect 47200 87366 47213 87418
rect 47265 87366 47277 87418
rect 47329 87366 47341 87418
rect 47393 87366 47405 87418
rect 47457 87366 47469 87418
rect 47521 87366 47533 87418
rect 47585 87366 47597 87418
rect 47649 87366 47662 87418
rect 47200 87360 47662 87366
rect 47857 87360 48114 87424
rect 49011 87420 49473 87426
rect 49011 87368 49024 87420
rect 49076 87368 49088 87420
rect 49140 87368 49152 87420
rect 49204 87368 49216 87420
rect 49268 87368 49280 87420
rect 49332 87368 49344 87420
rect 49396 87368 49408 87420
rect 49460 87368 49473 87420
rect 49011 87362 49473 87368
rect 47958 86910 48022 87360
rect 49667 87354 49906 87418
rect 50806 87416 51268 87422
rect 50806 87364 50819 87416
rect 50871 87364 50883 87416
rect 50935 87364 50947 87416
rect 50999 87364 51011 87416
rect 51063 87364 51075 87416
rect 51127 87364 51139 87416
rect 51191 87364 51203 87416
rect 51255 87364 51268 87416
rect 50806 87358 51268 87364
rect 51471 87359 51702 87423
rect 52605 87414 53067 87420
rect 52605 87362 52618 87414
rect 52670 87362 52682 87414
rect 52734 87362 52746 87414
rect 52798 87362 52810 87414
rect 52862 87362 52874 87414
rect 52926 87362 52938 87414
rect 52990 87362 53002 87414
rect 53054 87362 53067 87414
rect 49753 86910 49817 87354
rect 50145 87198 50405 87228
rect 50145 87018 50185 87198
rect 50365 87018 50405 87198
rect 50145 86988 50405 87018
rect 50237 86910 50301 86988
rect 51553 86910 51617 87359
rect 52605 87356 53067 87362
rect 53262 87357 53522 87421
rect 54396 87418 54858 87424
rect 54396 87366 54409 87418
rect 54461 87366 54473 87418
rect 54525 87366 54537 87418
rect 54589 87366 54601 87418
rect 54653 87366 54665 87418
rect 54717 87366 54729 87418
rect 54781 87366 54793 87418
rect 54845 87366 54858 87418
rect 54396 87360 54858 87366
rect 55065 87361 55300 87425
rect 56198 87414 56660 87420
rect 56198 87362 56211 87414
rect 56263 87362 56275 87414
rect 56327 87362 56339 87414
rect 56391 87362 56403 87414
rect 56455 87362 56467 87414
rect 56519 87362 56531 87414
rect 56583 87362 56595 87414
rect 56647 87362 56660 87414
rect 53356 86910 53420 87357
rect 55160 86910 55224 87361
rect 56198 87356 56660 87362
rect 56873 87360 57092 87424
rect 56956 87163 57020 87360
rect 57841 87224 58391 87254
rect 57841 87163 57866 87224
rect 56956 87099 57866 87163
rect 56956 86910 57020 87099
rect 57841 87044 57866 87099
rect 58366 87044 58391 87224
rect 57841 87014 58391 87044
rect 47958 86846 57020 86910
rect 57431 84830 57623 84849
rect 50227 78618 50291 78619
rect 48527 78611 48611 78617
rect 48527 78559 48543 78611
rect 48595 78559 48611 78611
rect 48527 78553 48611 78559
rect 50218 78612 50302 78618
rect 50218 78560 50234 78612
rect 50286 78560 50302 78612
rect 50218 78554 50302 78560
rect 51923 78611 52007 78617
rect 51923 78559 51939 78611
rect 51991 78559 52007 78611
rect 47380 78419 47642 78425
rect 48537 78423 48601 78553
rect 50227 78425 50291 78554
rect 51923 78553 52007 78559
rect 53719 78611 53803 78617
rect 53719 78559 53735 78611
rect 53787 78559 53803 78611
rect 53719 78553 53803 78559
rect 55548 78611 55632 78617
rect 55548 78559 55564 78611
rect 55616 78559 55632 78611
rect 55548 78553 55632 78559
rect 47380 78367 47421 78419
rect 47473 78367 47485 78419
rect 47537 78367 47549 78419
rect 47601 78367 47642 78419
rect 47380 78361 47642 78367
rect 47864 78359 48603 78423
rect 49175 78418 49437 78424
rect 49175 78366 49216 78418
rect 49268 78366 49280 78418
rect 49332 78366 49344 78418
rect 49396 78366 49437 78418
rect 49175 78360 49437 78366
rect 49659 78361 50291 78425
rect 50975 78420 51237 78426
rect 51933 78425 51997 78553
rect 50975 78368 51016 78420
rect 51068 78368 51080 78420
rect 51132 78368 51144 78420
rect 51196 78368 51237 78420
rect 50975 78362 51237 78368
rect 51462 78361 51997 78425
rect 52773 78419 53035 78425
rect 53729 78423 53793 78553
rect 52773 78367 52814 78419
rect 52866 78367 52878 78419
rect 52930 78367 52942 78419
rect 52994 78367 53035 78419
rect 52773 78361 53035 78367
rect 53262 78361 53793 78423
rect 54571 78420 54833 78426
rect 55558 78424 55622 78553
rect 54571 78368 54612 78420
rect 54664 78368 54676 78420
rect 54728 78368 54740 78420
rect 54792 78368 54833 78420
rect 54571 78362 54833 78368
rect 55067 78360 55622 78424
rect 56374 78419 56636 78425
rect 56374 78367 56415 78419
rect 56467 78367 56479 78419
rect 56531 78367 56543 78419
rect 56595 78367 56636 78419
rect 56374 78361 56636 78367
rect 56869 78420 57344 78426
rect 56869 78368 57276 78420
rect 57328 78368 57344 78420
rect 56869 78362 57344 78368
rect 42301 77616 42449 77622
rect 42301 77564 42317 77616
rect 42369 77564 42381 77616
rect 42433 77564 42449 77616
rect 42301 77558 42449 77564
rect 49534 77616 49618 77622
rect 49534 77564 49550 77616
rect 49602 77564 49618 77616
rect 49534 77558 49618 77564
rect 50095 77616 50243 77622
rect 50095 77564 50111 77616
rect 50163 77564 50175 77616
rect 50227 77564 50243 77616
rect 50095 77558 50243 77564
rect 42312 77542 42440 77558
rect 57431 77162 57469 84830
rect 57585 77162 57623 84830
rect 57431 77143 57623 77162
rect 67261 84834 67655 84858
rect 40971 77008 47974 77020
rect 40971 76956 47702 77008
rect 47754 76956 47766 77008
rect 47818 76956 47974 77008
rect 40971 76945 47974 76956
rect 48230 75243 48334 75271
rect 48230 75191 48256 75243
rect 48308 75191 48334 75243
rect 48230 75179 48334 75191
rect 48230 75127 48256 75179
rect 48308 75127 48334 75179
rect 48230 75115 48334 75127
rect 48230 75063 48256 75115
rect 48308 75063 48334 75115
rect 48230 75036 48334 75063
rect 51396 75086 53216 75088
rect 47686 74953 48404 74959
rect 47686 74901 47702 74953
rect 47754 74901 47766 74953
rect 47818 74901 48404 74953
rect 47686 74895 48404 74901
rect 49550 74951 50243 74957
rect 49550 74899 50111 74951
rect 50163 74899 50175 74951
rect 50227 74899 50243 74951
rect 51396 74906 51416 75086
rect 53196 75046 53216 75086
rect 53722 75065 54568 75096
rect 53722 75046 53735 75065
rect 53196 75010 53735 75046
rect 54555 75046 54568 75065
rect 55429 75055 56339 75086
rect 55429 75046 55442 75055
rect 54555 75010 55442 75046
rect 56326 75046 56339 75055
rect 56326 75010 56951 75046
rect 53196 74976 53215 75010
rect 53249 74976 53287 75010
rect 53321 74976 53359 75010
rect 53393 74976 53431 75010
rect 53465 74976 53503 75010
rect 53537 74976 53575 75010
rect 53609 74976 53647 75010
rect 53681 74976 53719 75010
rect 54555 74976 54583 75010
rect 54617 74976 54655 75010
rect 54689 74976 54727 75010
rect 54761 74976 54799 75010
rect 54833 74976 54871 75010
rect 54905 74976 54943 75010
rect 54977 74976 55015 75010
rect 55049 74976 55087 75010
rect 55121 74976 55159 75010
rect 55193 74976 55231 75010
rect 55265 74976 55303 75010
rect 55337 74976 55375 75010
rect 55409 74976 55442 75010
rect 56345 74976 56383 75010
rect 56417 74976 56455 75010
rect 56489 74976 56527 75010
rect 56561 74976 56599 75010
rect 56633 74976 56671 75010
rect 56705 74976 56743 75010
rect 56777 74976 56815 75010
rect 56849 74976 56887 75010
rect 56921 74976 56951 75010
rect 53196 74949 53735 74976
rect 54555 74949 55442 74976
rect 53196 74941 55442 74949
rect 53196 74906 53216 74941
rect 53722 74918 54568 74941
rect 55429 74939 55442 74941
rect 56326 74941 56951 74976
rect 56326 74939 56339 74941
rect 55429 74908 56339 74939
rect 51396 74905 53216 74906
rect 49550 74893 50243 74899
rect 48210 74792 48324 74813
rect 48210 74740 48241 74792
rect 48293 74740 48324 74792
rect 57006 74783 57225 74796
rect 48210 74728 48324 74740
rect 48210 74676 48241 74728
rect 48293 74676 48324 74728
rect 48210 74664 48324 74676
rect 48210 74612 48241 74664
rect 48293 74612 48324 74664
rect 48210 74600 48324 74612
rect 48210 74548 48241 74600
rect 48293 74548 48324 74600
rect 48210 74536 48324 74548
rect 48210 74484 48241 74536
rect 48293 74484 48324 74536
rect 48210 74472 48324 74484
rect 48210 74420 48241 74472
rect 48293 74420 48324 74472
rect 48210 74400 48324 74420
rect 51152 74736 51356 74742
rect 30014 73736 30378 73742
rect 30014 73684 30042 73736
rect 30094 73684 30106 73736
rect 30158 73684 30170 73736
rect 30222 73684 30234 73736
rect 30286 73684 30298 73736
rect 30350 73684 30378 73736
rect 30014 73678 30378 73684
rect 31035 73469 31093 73490
rect 31035 73446 31047 73469
rect 31024 73440 31047 73446
rect 31081 73446 31093 73469
rect 31081 73440 31108 73446
rect 30676 73429 30947 73435
rect 30676 73377 30689 73429
rect 30741 73420 30753 73429
rect 30805 73420 30817 73429
rect 30869 73420 30881 73429
rect 30751 73386 30753 73420
rect 30741 73377 30753 73386
rect 30805 73377 30817 73386
rect 30869 73377 30881 73386
rect 30933 73377 30947 73429
rect 31024 73388 31040 73440
rect 31092 73388 31108 73440
rect 31024 73383 31108 73388
rect 31024 73382 31047 73383
rect 30676 73371 30947 73377
rect 31035 73349 31047 73382
rect 31081 73382 31108 73383
rect 31081 73349 31093 73382
rect 31035 73317 31093 73349
rect 31100 73194 31464 73200
rect 31100 73142 31128 73194
rect 31180 73142 31192 73194
rect 31244 73142 31256 73194
rect 31308 73142 31320 73194
rect 31372 73142 31384 73194
rect 31436 73142 31464 73194
rect 31100 73136 31464 73142
rect 51152 71804 51164 74736
rect 51344 71804 51356 74736
rect 51152 71798 51356 71804
rect 57006 71787 57025 74783
rect 57205 71787 57225 74783
rect 57006 71774 57225 71787
rect 67261 71662 67272 84834
rect 67644 71662 67655 84834
rect 67261 71639 67655 71662
rect 51160 70294 51382 70296
rect 29997 67318 30114 67335
rect 29997 67266 30029 67318
rect 30081 67266 30114 67318
rect 29997 67254 30114 67266
rect 29997 67202 30029 67254
rect 30081 67202 30114 67254
rect 29997 67190 30114 67202
rect 29997 67138 30029 67190
rect 30081 67138 30114 67190
rect 29997 67126 30114 67138
rect 29997 67074 30029 67126
rect 30081 67074 30114 67126
rect 29997 67062 30114 67074
rect 29997 67010 30029 67062
rect 30081 67010 30114 67062
rect 43615 67077 43699 67083
rect 43615 67025 43631 67077
rect 43683 67025 43699 67077
rect 43615 67019 43699 67025
rect 29997 66998 30114 67010
rect 29997 66946 30029 66998
rect 30081 66946 30114 66998
rect 29997 66934 30114 66946
rect 29997 66882 30029 66934
rect 30081 66882 30114 66934
rect 29997 66870 30114 66882
rect 29997 66818 30029 66870
rect 30081 66818 30114 66870
rect 29997 66801 30114 66818
rect 30002 66177 30109 66191
rect 30002 66125 30029 66177
rect 30081 66125 30109 66177
rect 30002 66113 30109 66125
rect 30002 66061 30029 66113
rect 30081 66061 30109 66113
rect 30002 66049 30109 66061
rect 30002 65997 30029 66049
rect 30081 65997 30109 66049
rect 30002 65985 30109 65997
rect 30002 65933 30029 65985
rect 30081 65933 30109 65985
rect 30002 65921 30109 65933
rect 30002 65869 30029 65921
rect 30081 65869 30109 65921
rect 30002 65857 30109 65869
rect 30002 65805 30029 65857
rect 30081 65805 30109 65857
rect 30002 65793 30109 65805
rect 30002 65741 30029 65793
rect 30081 65741 30109 65793
rect 30002 65729 30109 65741
rect 30002 65677 30029 65729
rect 30081 65677 30109 65729
rect 30002 65665 30109 65677
rect 30002 65613 30029 65665
rect 30081 65613 30109 65665
rect 30002 65601 30109 65613
rect 30002 65549 30029 65601
rect 30081 65549 30109 65601
rect 30002 65537 30109 65549
rect 30002 65485 30029 65537
rect 30081 65485 30109 65537
rect 30002 65473 30109 65485
rect 30002 65421 30029 65473
rect 30081 65421 30109 65473
rect 30002 65409 30109 65421
rect 30002 65357 30029 65409
rect 30081 65357 30109 65409
rect 30002 65345 30109 65357
rect 30002 65293 30029 65345
rect 30081 65293 30109 65345
rect 30002 65281 30109 65293
rect 30002 65229 30029 65281
rect 30081 65229 30109 65281
rect 30002 65217 30109 65229
rect 30002 65165 30029 65217
rect 30081 65165 30109 65217
rect 30002 65153 30109 65165
rect 30002 65101 30029 65153
rect 30081 65101 30109 65153
rect 30002 65089 30109 65101
rect 30002 65037 30029 65089
rect 30081 65037 30109 65089
rect 30002 65024 30109 65037
rect 30007 64651 30114 64665
rect 30007 64599 30034 64651
rect 30086 64599 30114 64651
rect 30007 64587 30114 64599
rect 30007 64535 30034 64587
rect 30086 64535 30114 64587
rect 30007 64523 30114 64535
rect 30007 64471 30034 64523
rect 30086 64471 30114 64523
rect 30007 64459 30114 64471
rect 30007 64407 30034 64459
rect 30086 64407 30114 64459
rect 30007 64395 30114 64407
rect 30007 64343 30034 64395
rect 30086 64343 30114 64395
rect 30007 64331 30114 64343
rect 30007 64279 30034 64331
rect 30086 64279 30114 64331
rect 30007 64267 30114 64279
rect 30007 64215 30034 64267
rect 30086 64215 30114 64267
rect 30007 64203 30114 64215
rect 30007 64151 30034 64203
rect 30086 64151 30114 64203
rect 30007 64139 30114 64151
rect 30007 64087 30034 64139
rect 30086 64087 30114 64139
rect 30007 64075 30114 64087
rect 30007 64023 30034 64075
rect 30086 64023 30114 64075
rect 30007 64011 30114 64023
rect 30007 63959 30034 64011
rect 30086 63959 30114 64011
rect 30007 63947 30114 63959
rect 30007 63895 30034 63947
rect 30086 63895 30114 63947
rect 30007 63883 30114 63895
rect 30007 63831 30034 63883
rect 30086 63831 30114 63883
rect 30007 63819 30114 63831
rect 30007 63767 30034 63819
rect 30086 63767 30114 63819
rect 30007 63755 30114 63767
rect 30007 63703 30034 63755
rect 30086 63703 30114 63755
rect 30007 63691 30114 63703
rect 30007 63639 30034 63691
rect 30086 63639 30114 63691
rect 30007 63627 30114 63639
rect 30007 63575 30034 63627
rect 30086 63575 30114 63627
rect 30007 63563 30114 63575
rect 30007 63511 30034 63563
rect 30086 63511 30114 63563
rect 30007 63498 30114 63511
rect 38201 63542 38297 63559
rect 38201 63490 38223 63542
rect 38275 63490 38297 63542
rect 38201 63478 38297 63490
rect 38201 63426 38223 63478
rect 38275 63426 38297 63478
rect 38201 63414 38297 63426
rect 38201 63362 38223 63414
rect 38275 63362 38297 63414
rect 38201 63350 38297 63362
rect 38201 63298 38223 63350
rect 38275 63298 38297 63350
rect 38201 63286 38297 63298
rect 38201 63234 38223 63286
rect 38275 63234 38297 63286
rect 38201 63222 38297 63234
rect 25272 63172 25356 63188
rect 25272 63120 25288 63172
rect 25340 63120 25356 63172
rect 38201 63170 38223 63222
rect 38275 63170 38297 63222
rect 25948 63148 26012 63163
rect 25272 63108 25299 63120
rect 25333 63108 25356 63120
rect 25545 63114 26012 63148
rect 38201 63158 38297 63170
rect 25272 63056 25288 63108
rect 25340 63056 25356 63108
rect 25272 63044 25299 63056
rect 25333 63044 25356 63056
rect 25272 63029 25288 63044
rect 25263 62995 25288 63029
rect 25272 62992 25288 62995
rect 25340 63029 25356 63044
rect 25340 62995 25384 63029
rect 25340 62992 25356 62995
rect 25272 62980 25299 62992
rect 25333 62980 25356 62992
rect 25272 62928 25288 62980
rect 25340 62928 25356 62980
rect 25272 62920 25356 62928
rect 25272 62916 25299 62920
rect 25333 62916 25356 62920
rect 25272 62864 25288 62916
rect 25340 62864 25356 62916
rect 25948 62908 26012 63114
rect 25541 62874 26012 62908
rect 25272 62849 25356 62864
rect 25273 62617 25357 62635
rect 25273 62565 25289 62617
rect 25341 62565 25357 62617
rect 25948 62592 26012 62874
rect 25273 62553 25299 62565
rect 25333 62553 25357 62565
rect 25541 62558 26012 62592
rect 25273 62501 25289 62553
rect 25341 62501 25357 62553
rect 25273 62500 25357 62501
rect 25273 62489 25299 62500
rect 25333 62489 25357 62500
rect 25273 62437 25289 62489
rect 25341 62437 25357 62489
rect 25273 62429 25357 62437
rect 25263 62428 25360 62429
rect 25263 62425 25299 62428
rect 25333 62425 25360 62428
rect 25263 62395 25289 62425
rect 25273 62373 25289 62395
rect 25341 62395 25360 62425
rect 25341 62373 25357 62395
rect 25273 62361 25357 62373
rect 25273 62309 25289 62361
rect 25341 62309 25357 62361
rect 25273 62297 25357 62309
rect 25273 62245 25289 62297
rect 25341 62245 25357 62297
rect 25948 62278 26012 62558
rect 30002 63140 30106 63142
rect 30002 63088 30028 63140
rect 30080 63088 30106 63140
rect 30002 63076 30106 63088
rect 30002 63024 30028 63076
rect 30080 63024 30106 63076
rect 30002 63012 30106 63024
rect 30002 62960 30028 63012
rect 30080 62960 30106 63012
rect 30002 62948 30106 62960
rect 30002 62896 30028 62948
rect 30080 62896 30106 62948
rect 30002 62884 30106 62896
rect 30002 62832 30028 62884
rect 30080 62832 30106 62884
rect 30002 62820 30106 62832
rect 30002 62768 30028 62820
rect 30080 62768 30106 62820
rect 30002 62756 30106 62768
rect 30002 62704 30028 62756
rect 30080 62704 30106 62756
rect 30002 62692 30106 62704
rect 30002 62640 30028 62692
rect 30080 62640 30106 62692
rect 30002 62628 30106 62640
rect 30002 62576 30028 62628
rect 30080 62576 30106 62628
rect 30002 62564 30106 62576
rect 30002 62512 30028 62564
rect 30080 62512 30106 62564
rect 30002 62500 30106 62512
rect 30002 62448 30028 62500
rect 30080 62448 30106 62500
rect 30002 62436 30106 62448
rect 27470 62429 27954 62435
rect 27470 62377 27494 62429
rect 27546 62377 27558 62429
rect 27610 62377 27622 62429
rect 27674 62377 27686 62429
rect 27738 62377 27750 62429
rect 27802 62377 27814 62429
rect 27866 62377 27878 62429
rect 27930 62377 27954 62429
rect 27470 62371 27954 62377
rect 30002 62384 30028 62436
rect 30080 62384 30106 62436
rect 30002 62372 30106 62384
rect 30002 62320 30028 62372
rect 30080 62320 30106 62372
rect 30002 62308 30106 62320
rect 25935 62272 27390 62278
rect 25935 62264 26070 62272
rect 25273 62233 25357 62245
rect 25273 62181 25289 62233
rect 25341 62181 25357 62233
rect 25541 62230 26070 62264
rect 25935 62220 26070 62230
rect 26122 62220 26134 62272
rect 26186 62220 27390 62272
rect 30002 62256 30028 62308
rect 30080 62256 30106 62308
rect 30002 62254 30106 62256
rect 38201 63106 38223 63158
rect 38275 63106 38297 63158
rect 38201 63094 38297 63106
rect 38201 63042 38223 63094
rect 38275 63042 38297 63094
rect 38201 63030 38297 63042
rect 38201 62978 38223 63030
rect 38275 62978 38297 63030
rect 38201 62966 38297 62978
rect 38201 62914 38223 62966
rect 38275 62914 38297 62966
rect 38201 62902 38297 62914
rect 38201 62850 38223 62902
rect 38275 62850 38297 62902
rect 38201 62838 38297 62850
rect 38201 62786 38223 62838
rect 38275 62786 38297 62838
rect 38201 62774 38297 62786
rect 38201 62722 38223 62774
rect 38275 62722 38297 62774
rect 38201 62710 38297 62722
rect 38201 62658 38223 62710
rect 38275 62658 38297 62710
rect 38201 62646 38297 62658
rect 38201 62594 38223 62646
rect 38275 62594 38297 62646
rect 38201 62582 38297 62594
rect 38201 62530 38223 62582
rect 38275 62530 38297 62582
rect 38201 62518 38297 62530
rect 38201 62466 38223 62518
rect 38275 62466 38297 62518
rect 38201 62454 38297 62466
rect 38201 62402 38223 62454
rect 38275 62402 38297 62454
rect 38201 62390 38297 62402
rect 38201 62338 38223 62390
rect 38275 62338 38297 62390
rect 38201 62326 38297 62338
rect 38201 62274 38223 62326
rect 38275 62274 38297 62326
rect 38201 62262 38297 62274
rect 25935 62214 27390 62220
rect 25273 62163 25357 62181
rect 38201 62210 38223 62262
rect 38275 62210 38297 62262
rect 38201 62198 38297 62210
rect 38201 62146 38223 62198
rect 38275 62146 38297 62198
rect 38201 62134 38297 62146
rect 38201 62082 38223 62134
rect 38275 62082 38297 62134
rect 38201 62070 38297 62082
rect 38201 62018 38223 62070
rect 38275 62018 38297 62070
rect 38201 62006 38297 62018
rect 38201 61954 38223 62006
rect 38275 61954 38297 62006
rect 38201 61942 38297 61954
rect 38201 61890 38223 61942
rect 38275 61890 38297 61942
rect 38201 61878 38297 61890
rect 38201 61826 38223 61878
rect 38275 61826 38297 61878
rect 38201 61814 38297 61826
rect 38201 61762 38223 61814
rect 38275 61762 38297 61814
rect 38201 61750 38297 61762
rect 38201 61698 38223 61750
rect 38275 61698 38297 61750
rect 38201 61686 38297 61698
rect 38201 61634 38223 61686
rect 38275 61634 38297 61686
rect 38201 61622 38297 61634
rect 21566 61562 21822 61590
rect 21566 61382 21604 61562
rect 21784 61497 21822 61562
rect 38201 61570 38223 61622
rect 38275 61570 38297 61622
rect 38201 61558 38297 61570
rect 38201 61506 38223 61558
rect 38275 61506 38297 61558
rect 21784 61491 27398 61497
rect 21784 61439 26901 61491
rect 26953 61439 26965 61491
rect 27017 61439 27398 61491
rect 21784 61433 27398 61439
rect 38201 61494 38297 61506
rect 38201 61442 38223 61494
rect 38275 61442 38297 61494
rect 21784 61382 21822 61433
rect 21566 61354 21822 61382
rect 38201 61430 38297 61442
rect 38201 61378 38223 61430
rect 38275 61378 38297 61430
rect 30005 61373 30109 61375
rect 27432 61339 27961 61345
rect 27432 61287 27446 61339
rect 27498 61287 27510 61339
rect 27562 61287 27574 61339
rect 27626 61287 27638 61339
rect 27690 61287 27702 61339
rect 27754 61287 27766 61339
rect 27818 61287 27830 61339
rect 27882 61287 27894 61339
rect 27946 61287 27961 61339
rect 27432 61281 27961 61287
rect 30005 61321 30031 61373
rect 30083 61321 30109 61373
rect 30005 61309 30109 61321
rect 30005 61257 30031 61309
rect 30083 61257 30109 61309
rect 30005 61245 30109 61257
rect 30005 61193 30031 61245
rect 30083 61193 30109 61245
rect 30005 61181 30109 61193
rect 30005 61129 30031 61181
rect 30083 61129 30109 61181
rect 30005 61117 30109 61129
rect 30005 61065 30031 61117
rect 30083 61065 30109 61117
rect 30005 61053 30109 61065
rect 30005 61001 30031 61053
rect 30083 61001 30109 61053
rect 30005 60989 30109 61001
rect 30005 60937 30031 60989
rect 30083 60937 30109 60989
rect 30005 60925 30109 60937
rect 30005 60873 30031 60925
rect 30083 60873 30109 60925
rect 30005 60861 30109 60873
rect 30005 60809 30031 60861
rect 30083 60809 30109 60861
rect 30005 60797 30109 60809
rect 30005 60745 30031 60797
rect 30083 60745 30109 60797
rect 30005 60733 30109 60745
rect 30005 60681 30031 60733
rect 30083 60681 30109 60733
rect 30005 60669 30109 60681
rect 30005 60617 30031 60669
rect 30083 60617 30109 60669
rect 30005 60605 30109 60617
rect 30005 60553 30031 60605
rect 30083 60553 30109 60605
rect 30005 60541 30109 60553
rect 30005 60489 30031 60541
rect 30083 60489 30109 60541
rect 30005 60487 30109 60489
rect 38201 61366 38297 61378
rect 38201 61314 38223 61366
rect 38275 61314 38297 61366
rect 38201 61302 38297 61314
rect 38201 61250 38223 61302
rect 38275 61250 38297 61302
rect 38201 61238 38297 61250
rect 38201 61186 38223 61238
rect 38275 61186 38297 61238
rect 38201 61174 38297 61186
rect 38201 61122 38223 61174
rect 38275 61122 38297 61174
rect 38201 61110 38297 61122
rect 38201 61058 38223 61110
rect 38275 61058 38297 61110
rect 38201 61046 38297 61058
rect 38201 60994 38223 61046
rect 38275 60994 38297 61046
rect 38201 60982 38297 60994
rect 38201 60930 38223 60982
rect 38275 60930 38297 60982
rect 38201 60918 38297 60930
rect 38201 60866 38223 60918
rect 38275 60866 38297 60918
rect 38201 60854 38297 60866
rect 38201 60802 38223 60854
rect 38275 60802 38297 60854
rect 38201 60790 38297 60802
rect 38201 60738 38223 60790
rect 38275 60738 38297 60790
rect 38201 60726 38297 60738
rect 38201 60674 38223 60726
rect 38275 60674 38297 60726
rect 38201 60662 38297 60674
rect 38201 60610 38223 60662
rect 38275 60610 38297 60662
rect 38201 60598 38297 60610
rect 38201 60546 38223 60598
rect 38275 60546 38297 60598
rect 38201 60534 38297 60546
rect 38201 60482 38223 60534
rect 38275 60482 38297 60534
rect 38201 60470 38297 60482
rect 38201 60418 38223 60470
rect 38275 60418 38297 60470
rect 38201 60406 38297 60418
rect 38201 60354 38223 60406
rect 38275 60354 38297 60406
rect 38201 60342 38297 60354
rect 38201 60290 38223 60342
rect 38275 60290 38297 60342
rect 38201 60278 38297 60290
rect 38201 60226 38223 60278
rect 38275 60226 38297 60278
rect 38201 60214 38297 60226
rect 30007 60164 30108 60182
rect 30007 60112 30031 60164
rect 30083 60112 30108 60164
rect 38201 60162 38223 60214
rect 38275 60162 38297 60214
rect 38201 60146 38297 60162
rect 30007 60100 30108 60112
rect 30007 60048 30031 60100
rect 30083 60048 30108 60100
rect 30007 60036 30108 60048
rect 30007 59984 30031 60036
rect 30083 59984 30108 60036
rect 30007 59972 30108 59984
rect 30007 59920 30031 59972
rect 30083 59920 30108 59972
rect 30007 59908 30108 59920
rect 30007 59856 30031 59908
rect 30083 59856 30108 59908
rect 30007 59844 30108 59856
rect 30007 59792 30031 59844
rect 30083 59792 30108 59844
rect 30007 59780 30108 59792
rect 30007 59728 30031 59780
rect 30083 59728 30108 59780
rect 30007 59716 30108 59728
rect 30007 59664 30031 59716
rect 30083 59664 30108 59716
rect 30007 59652 30108 59664
rect 30007 59600 30031 59652
rect 30083 59600 30108 59652
rect 30007 59588 30108 59600
rect 30007 59536 30031 59588
rect 30083 59536 30108 59588
rect 30007 59524 30108 59536
rect 30007 59472 30031 59524
rect 30083 59472 30108 59524
rect 30007 59460 30108 59472
rect 30007 59408 30031 59460
rect 30083 59408 30108 59460
rect 30007 59396 30108 59408
rect 30007 59344 30031 59396
rect 30083 59344 30108 59396
rect 30007 59332 30108 59344
rect 30007 59280 30031 59332
rect 30083 59280 30108 59332
rect 30007 59268 30108 59280
rect 30007 59216 30031 59268
rect 30083 59216 30108 59268
rect 30007 59204 30108 59216
rect 30007 59152 30031 59204
rect 30083 59152 30108 59204
rect 30007 59140 30108 59152
rect 30007 59088 30031 59140
rect 30083 59088 30108 59140
rect 30007 59076 30108 59088
rect 30007 59024 30031 59076
rect 30083 59024 30108 59076
rect 30007 59007 30108 59024
rect 30005 58686 30104 58713
rect 30005 58634 30028 58686
rect 30080 58634 30104 58686
rect 30005 58622 30104 58634
rect 30005 58570 30028 58622
rect 30080 58570 30104 58622
rect 30005 58558 30104 58570
rect 30005 58506 30028 58558
rect 30080 58506 30104 58558
rect 30005 58494 30104 58506
rect 30005 58442 30028 58494
rect 30080 58442 30104 58494
rect 30005 58430 30104 58442
rect 30005 58378 30028 58430
rect 30080 58378 30104 58430
rect 30005 58366 30104 58378
rect 30005 58314 30028 58366
rect 30080 58314 30104 58366
rect 30005 58302 30104 58314
rect 30005 58250 30028 58302
rect 30080 58250 30104 58302
rect 30005 58238 30104 58250
rect 30005 58186 30028 58238
rect 30080 58186 30104 58238
rect 30005 58174 30104 58186
rect 30005 58122 30028 58174
rect 30080 58122 30104 58174
rect 30005 58110 30104 58122
rect 30005 58058 30028 58110
rect 30080 58058 30104 58110
rect 30005 58046 30104 58058
rect 30005 57994 30028 58046
rect 30080 57994 30104 58046
rect 30005 57982 30104 57994
rect 30005 57930 30028 57982
rect 30080 57930 30104 57982
rect 30005 57918 30104 57930
rect 30005 57866 30028 57918
rect 30080 57866 30104 57918
rect 30005 57854 30104 57866
rect 30005 57802 30028 57854
rect 30080 57802 30104 57854
rect 30005 57790 30104 57802
rect 30005 57738 30028 57790
rect 30080 57738 30104 57790
rect 30005 57726 30104 57738
rect 30005 57674 30028 57726
rect 30080 57674 30104 57726
rect 30005 57662 30104 57674
rect 30005 57610 30028 57662
rect 30080 57610 30104 57662
rect 30005 57598 30104 57610
rect 30005 57546 30028 57598
rect 30080 57546 30104 57598
rect 30005 57520 30104 57546
rect 30000 56904 30099 56921
rect 30000 56852 30023 56904
rect 30075 56852 30099 56904
rect 30000 56840 30099 56852
rect 30000 56788 30023 56840
rect 30075 56788 30099 56840
rect 30000 56776 30099 56788
rect 30000 56724 30023 56776
rect 30075 56724 30099 56776
rect 30000 56712 30099 56724
rect 30000 56660 30023 56712
rect 30075 56660 30099 56712
rect 30000 56648 30099 56660
rect 30000 56596 30023 56648
rect 30075 56596 30099 56648
rect 30000 56584 30099 56596
rect 30000 56532 30023 56584
rect 30075 56532 30099 56584
rect 30000 56520 30099 56532
rect 30000 56468 30023 56520
rect 30075 56468 30099 56520
rect 30000 56456 30099 56468
rect 30000 56404 30023 56456
rect 30075 56404 30099 56456
rect 30000 56387 30099 56404
rect 43625 53351 43689 67019
rect 44391 66414 44475 66420
rect 44391 66362 44407 66414
rect 44459 66362 44475 66414
rect 44391 66356 44475 66362
rect 44401 53774 44465 66356
rect 51160 63842 51181 70294
rect 51361 63842 51382 70294
rect 67264 70149 67655 70150
rect 57428 69865 57662 69866
rect 57187 69387 57251 69388
rect 56525 69335 57251 69387
rect 51160 63841 51382 63842
rect 50105 63827 50233 63828
rect 47686 63821 47834 63827
rect 47686 63769 47702 63821
rect 47754 63769 47766 63821
rect 47818 63769 47834 63821
rect 47686 63763 47834 63769
rect 50095 63821 50243 63827
rect 50095 63769 50111 63821
rect 50163 63769 50175 63821
rect 50227 63769 50243 63821
rect 50095 63763 50243 63769
rect 47696 58692 47824 63763
rect 47696 58640 47731 58692
rect 47783 58640 47824 58692
rect 47696 54327 47824 58640
rect 50105 57195 50233 63763
rect 51400 63688 51432 63868
rect 56924 63688 56956 63868
rect 57187 62588 57251 69335
rect 57428 68341 57455 69865
rect 57635 68341 57662 69865
rect 57428 68340 57662 68341
rect 57436 65403 57616 65405
rect 57436 63879 57468 65403
rect 57584 63879 57616 65403
rect 64176 65328 64294 67034
rect 57436 63877 57616 63879
rect 59597 62873 59699 62903
rect 59597 62821 59622 62873
rect 59674 62821 59699 62873
rect 59597 62809 59699 62821
rect 59597 62757 59622 62809
rect 59674 62757 59699 62809
rect 59597 62745 59699 62757
rect 59597 62693 59622 62745
rect 59674 62693 59699 62745
rect 59597 62664 59699 62693
rect 62455 62590 62519 64460
rect 57177 62582 57261 62588
rect 57177 62530 57193 62582
rect 57245 62530 57261 62582
rect 57177 62524 57261 62530
rect 58314 62582 58398 62588
rect 58314 62530 58330 62582
rect 58382 62530 58398 62582
rect 58314 62524 58398 62530
rect 59533 62584 59794 62590
rect 59533 62532 59726 62584
rect 59778 62532 59794 62584
rect 59533 62526 59794 62532
rect 62445 62584 62529 62590
rect 62445 62532 62461 62584
rect 62513 62532 62529 62584
rect 62445 62526 62529 62532
rect 57187 61673 57251 62524
rect 59599 62416 59718 62442
rect 59599 62364 59632 62416
rect 59684 62364 59718 62416
rect 59599 62352 59718 62364
rect 59599 62300 59632 62352
rect 59684 62300 59718 62352
rect 59599 62288 59718 62300
rect 59599 62236 59632 62288
rect 59684 62236 59718 62288
rect 59599 62224 59718 62236
rect 59599 62172 59632 62224
rect 59684 62172 59718 62224
rect 62455 62177 62519 62526
rect 59599 62160 59718 62172
rect 59599 62108 59632 62160
rect 59684 62108 59718 62160
rect 62445 62171 62529 62177
rect 62445 62119 62461 62171
rect 62513 62119 62529 62171
rect 62445 62113 62529 62119
rect 59599 62096 59718 62108
rect 59599 62044 59632 62096
rect 59684 62044 59718 62096
rect 59599 62018 59718 62044
rect 57177 61667 57261 61673
rect 57177 61615 57193 61667
rect 57245 61615 57261 61667
rect 57177 61609 57261 61615
rect 60511 61667 60595 61673
rect 60511 61615 60527 61667
rect 60579 61615 60595 61667
rect 60511 61609 60595 61615
rect 57187 60838 57251 61609
rect 59728 61223 59812 61229
rect 59728 61171 59744 61223
rect 59796 61171 59812 61223
rect 59252 61167 59336 61171
rect 59252 61115 59268 61167
rect 59320 61115 59336 61167
rect 59728 61165 59812 61171
rect 59252 61103 59336 61115
rect 59252 61051 59268 61103
rect 59320 61051 59336 61103
rect 59252 61039 59336 61051
rect 59252 60987 59268 61039
rect 59320 60987 59336 61039
rect 59252 60975 59336 60987
rect 59252 60923 59268 60975
rect 59320 60923 59336 60975
rect 59252 60920 59336 60923
rect 59738 60838 59802 61165
rect 57177 60832 57261 60838
rect 57177 60780 57193 60832
rect 57245 60780 57261 60832
rect 57177 60774 57261 60780
rect 57967 60832 58051 60838
rect 57967 60780 57983 60832
rect 58035 60780 58051 60832
rect 57967 60774 58051 60780
rect 59334 60774 59802 60838
rect 57187 60772 57251 60774
rect 59253 60667 59337 60690
rect 59253 60615 59269 60667
rect 59321 60615 59337 60667
rect 59253 60603 59337 60615
rect 59253 60551 59269 60603
rect 59321 60551 59337 60603
rect 59253 60539 59337 60551
rect 59253 60487 59269 60539
rect 59321 60487 59337 60539
rect 59253 60475 59337 60487
rect 59253 60423 59269 60475
rect 59321 60423 59337 60475
rect 59253 60411 59337 60423
rect 59253 60359 59269 60411
rect 59321 60359 59337 60411
rect 59253 60347 59337 60359
rect 59253 60295 59269 60347
rect 59321 60295 59337 60347
rect 59253 60272 59337 60295
rect 60022 60107 60447 60110
rect 60022 60055 60048 60107
rect 60100 60055 60112 60107
rect 60164 60055 60176 60107
rect 60228 60055 60240 60107
rect 60292 60055 60304 60107
rect 60356 60055 60368 60107
rect 60420 60055 60447 60107
rect 60022 60052 60447 60055
rect 60521 59972 60585 61609
rect 63795 61229 63859 64471
rect 64176 63232 64412 65328
rect 67264 63889 67305 70149
rect 67613 63889 67655 70149
rect 69636 63232 69872 97041
rect 81750 90723 81986 101898
rect 81844 89763 81890 90723
rect 74514 88760 74600 88765
rect 74514 88708 74531 88760
rect 74583 88708 74600 88760
rect 74514 88696 74600 88708
rect 74514 88644 74531 88696
rect 74583 88644 74600 88696
rect 74514 88632 74600 88644
rect 74514 88580 74531 88632
rect 74583 88580 74600 88632
rect 74514 88568 74600 88580
rect 74514 88516 74531 88568
rect 74583 88516 74600 88568
rect 74514 88504 74600 88516
rect 74514 88452 74531 88504
rect 74583 88452 74600 88504
rect 74514 88440 74600 88452
rect 74514 88388 74531 88440
rect 74583 88388 74600 88440
rect 74514 88376 74600 88388
rect 74514 88324 74531 88376
rect 74583 88324 74600 88376
rect 74514 88312 74600 88324
rect 74514 88260 74531 88312
rect 74583 88260 74600 88312
rect 74514 88248 74600 88260
rect 74514 88196 74531 88248
rect 74583 88196 74600 88248
rect 74514 88191 74600 88196
rect 81042 88760 81128 88765
rect 81042 88708 81059 88760
rect 81111 88708 81128 88760
rect 81042 88696 81128 88708
rect 81042 88644 81059 88696
rect 81111 88644 81128 88696
rect 81042 88632 81128 88644
rect 81042 88580 81059 88632
rect 81111 88580 81128 88632
rect 81042 88568 81128 88580
rect 81042 88516 81059 88568
rect 81111 88516 81128 88568
rect 81042 88504 81128 88516
rect 81042 88452 81059 88504
rect 81111 88452 81128 88504
rect 81042 88440 81128 88452
rect 81042 88388 81059 88440
rect 81111 88388 81128 88440
rect 81042 88376 81128 88388
rect 81042 88324 81059 88376
rect 81111 88324 81128 88376
rect 81042 88312 81128 88324
rect 81042 88260 81059 88312
rect 81111 88260 81128 88312
rect 81042 88248 81128 88260
rect 81042 88196 81059 88248
rect 81111 88196 81128 88248
rect 81042 88191 81128 88196
rect 88658 88760 88744 88765
rect 88658 88708 88675 88760
rect 88727 88708 88744 88760
rect 88658 88696 88744 88708
rect 88658 88644 88675 88696
rect 88727 88644 88744 88696
rect 88658 88632 88744 88644
rect 88658 88580 88675 88632
rect 88727 88580 88744 88632
rect 88658 88568 88744 88580
rect 88658 88516 88675 88568
rect 88727 88516 88744 88568
rect 88658 88504 88744 88516
rect 88658 88452 88675 88504
rect 88727 88452 88744 88504
rect 88658 88440 88744 88452
rect 88658 88388 88675 88440
rect 88727 88388 88744 88440
rect 88658 88376 88744 88388
rect 88658 88324 88675 88376
rect 88727 88324 88744 88376
rect 88658 88312 88744 88324
rect 88658 88260 88675 88312
rect 88727 88260 88744 88312
rect 88658 88248 88744 88260
rect 88658 88196 88675 88248
rect 88727 88196 88744 88248
rect 88658 88191 88744 88196
rect 75059 86757 75145 86762
rect 75059 86705 75076 86757
rect 75128 86705 75145 86757
rect 75059 86693 75145 86705
rect 75059 86641 75076 86693
rect 75128 86641 75145 86693
rect 75059 86629 75145 86641
rect 75059 86577 75076 86629
rect 75128 86577 75145 86629
rect 75059 86565 75145 86577
rect 75059 86513 75076 86565
rect 75128 86513 75145 86565
rect 75059 86501 75145 86513
rect 75059 86449 75076 86501
rect 75128 86449 75145 86501
rect 75059 86437 75145 86449
rect 75059 86385 75076 86437
rect 75128 86385 75145 86437
rect 75059 86373 75145 86385
rect 75059 86321 75076 86373
rect 75128 86321 75145 86373
rect 75059 86309 75145 86321
rect 75059 86257 75076 86309
rect 75128 86257 75145 86309
rect 75059 86245 75145 86257
rect 75059 86193 75076 86245
rect 75128 86193 75145 86245
rect 75059 86188 75145 86193
rect 76147 86757 76233 86762
rect 76147 86705 76164 86757
rect 76216 86705 76233 86757
rect 76147 86693 76233 86705
rect 76147 86641 76164 86693
rect 76216 86641 76233 86693
rect 76147 86629 76233 86641
rect 76147 86577 76164 86629
rect 76216 86577 76233 86629
rect 76147 86565 76233 86577
rect 76147 86513 76164 86565
rect 76216 86513 76233 86565
rect 76147 86501 76233 86513
rect 76147 86449 76164 86501
rect 76216 86449 76233 86501
rect 76147 86437 76233 86449
rect 76147 86385 76164 86437
rect 76216 86385 76233 86437
rect 76147 86373 76233 86385
rect 76147 86321 76164 86373
rect 76216 86321 76233 86373
rect 76147 86309 76233 86321
rect 76147 86257 76164 86309
rect 76216 86257 76233 86309
rect 76147 86245 76233 86257
rect 76147 86193 76164 86245
rect 76216 86193 76233 86245
rect 76147 86188 76233 86193
rect 78323 86757 78409 86762
rect 78323 86705 78340 86757
rect 78392 86705 78409 86757
rect 78323 86693 78409 86705
rect 78323 86641 78340 86693
rect 78392 86641 78409 86693
rect 78323 86629 78409 86641
rect 78323 86577 78340 86629
rect 78392 86577 78409 86629
rect 78323 86565 78409 86577
rect 78323 86513 78340 86565
rect 78392 86513 78409 86565
rect 78323 86501 78409 86513
rect 78323 86449 78340 86501
rect 78392 86449 78409 86501
rect 78323 86437 78409 86449
rect 78323 86385 78340 86437
rect 78392 86385 78409 86437
rect 78323 86373 78409 86385
rect 78323 86321 78340 86373
rect 78392 86321 78409 86373
rect 78323 86309 78409 86321
rect 78323 86257 78340 86309
rect 78392 86257 78409 86309
rect 78323 86245 78409 86257
rect 78323 86193 78340 86245
rect 78392 86193 78409 86245
rect 78323 86188 78409 86193
rect 79411 86757 79497 86762
rect 79411 86705 79428 86757
rect 79480 86705 79497 86757
rect 79411 86693 79497 86705
rect 79411 86641 79428 86693
rect 79480 86641 79497 86693
rect 79411 86629 79497 86641
rect 79411 86577 79428 86629
rect 79480 86577 79497 86629
rect 79411 86565 79497 86577
rect 79411 86513 79428 86565
rect 79480 86513 79497 86565
rect 79411 86501 79497 86513
rect 79411 86449 79428 86501
rect 79480 86449 79497 86501
rect 79411 86437 79497 86449
rect 79411 86385 79428 86437
rect 79480 86385 79497 86437
rect 79411 86373 79497 86385
rect 79411 86321 79428 86373
rect 79480 86321 79497 86373
rect 79411 86309 79497 86321
rect 79411 86257 79428 86309
rect 79480 86257 79497 86309
rect 79411 86245 79497 86257
rect 79411 86193 79428 86245
rect 79480 86193 79497 86245
rect 79411 86188 79497 86193
rect 80499 86757 80585 86762
rect 80499 86705 80516 86757
rect 80568 86705 80585 86757
rect 80499 86693 80585 86705
rect 80499 86641 80516 86693
rect 80568 86641 80585 86693
rect 80499 86629 80585 86641
rect 80499 86577 80516 86629
rect 80568 86577 80585 86629
rect 80499 86565 80585 86577
rect 80499 86513 80516 86565
rect 80568 86513 80585 86565
rect 80499 86501 80585 86513
rect 80499 86449 80516 86501
rect 80568 86449 80585 86501
rect 80499 86437 80585 86449
rect 80499 86385 80516 86437
rect 80568 86385 80585 86437
rect 80499 86373 80585 86385
rect 80499 86321 80516 86373
rect 80568 86321 80585 86373
rect 80499 86309 80585 86321
rect 80499 86257 80516 86309
rect 80568 86257 80585 86309
rect 80499 86245 80585 86257
rect 80499 86193 80516 86245
rect 80568 86193 80585 86245
rect 80499 86188 80585 86193
rect 81587 86757 81673 86762
rect 81587 86705 81604 86757
rect 81656 86705 81673 86757
rect 81587 86693 81673 86705
rect 81587 86641 81604 86693
rect 81656 86641 81673 86693
rect 81587 86629 81673 86641
rect 81587 86577 81604 86629
rect 81656 86577 81673 86629
rect 81587 86565 81673 86577
rect 81587 86513 81604 86565
rect 81656 86513 81673 86565
rect 81587 86501 81673 86513
rect 81587 86449 81604 86501
rect 81656 86449 81673 86501
rect 81587 86437 81673 86449
rect 81587 86385 81604 86437
rect 81656 86385 81673 86437
rect 81587 86373 81673 86385
rect 81587 86321 81604 86373
rect 81656 86321 81673 86373
rect 81587 86309 81673 86321
rect 81587 86257 81604 86309
rect 81656 86257 81673 86309
rect 81587 86245 81673 86257
rect 81587 86193 81604 86245
rect 81656 86193 81673 86245
rect 81587 86188 81673 86193
rect 82675 86757 82761 86762
rect 82675 86705 82692 86757
rect 82744 86705 82761 86757
rect 82675 86693 82761 86705
rect 82675 86641 82692 86693
rect 82744 86641 82761 86693
rect 82675 86629 82761 86641
rect 82675 86577 82692 86629
rect 82744 86577 82761 86629
rect 82675 86565 82761 86577
rect 82675 86513 82692 86565
rect 82744 86513 82761 86565
rect 82675 86501 82761 86513
rect 82675 86449 82692 86501
rect 82744 86449 82761 86501
rect 82675 86437 82761 86449
rect 82675 86385 82692 86437
rect 82744 86385 82761 86437
rect 82675 86373 82761 86385
rect 82675 86321 82692 86373
rect 82744 86321 82761 86373
rect 82675 86309 82761 86321
rect 82675 86257 82692 86309
rect 82744 86257 82761 86309
rect 82675 86245 82761 86257
rect 82675 86193 82692 86245
rect 82744 86193 82761 86245
rect 82675 86188 82761 86193
rect 83763 86757 83849 86762
rect 83763 86705 83780 86757
rect 83832 86705 83849 86757
rect 83763 86693 83849 86705
rect 83763 86641 83780 86693
rect 83832 86641 83849 86693
rect 83763 86629 83849 86641
rect 83763 86577 83780 86629
rect 83832 86577 83849 86629
rect 83763 86565 83849 86577
rect 83763 86513 83780 86565
rect 83832 86513 83849 86565
rect 83763 86501 83849 86513
rect 83763 86449 83780 86501
rect 83832 86449 83849 86501
rect 83763 86437 83849 86449
rect 83763 86385 83780 86437
rect 83832 86385 83849 86437
rect 83763 86373 83849 86385
rect 83763 86321 83780 86373
rect 83832 86321 83849 86373
rect 83763 86309 83849 86321
rect 83763 86257 83780 86309
rect 83832 86257 83849 86309
rect 83763 86245 83849 86257
rect 83763 86193 83780 86245
rect 83832 86193 83849 86245
rect 83763 86188 83849 86193
rect 85939 86757 86025 86762
rect 85939 86705 85956 86757
rect 86008 86705 86025 86757
rect 85939 86693 86025 86705
rect 85939 86641 85956 86693
rect 86008 86641 86025 86693
rect 85939 86629 86025 86641
rect 85939 86577 85956 86629
rect 86008 86577 86025 86629
rect 85939 86565 86025 86577
rect 85939 86513 85956 86565
rect 86008 86513 86025 86565
rect 85939 86501 86025 86513
rect 85939 86449 85956 86501
rect 86008 86449 86025 86501
rect 85939 86437 86025 86449
rect 85939 86385 85956 86437
rect 86008 86385 86025 86437
rect 85939 86373 86025 86385
rect 85939 86321 85956 86373
rect 86008 86321 86025 86373
rect 85939 86309 86025 86321
rect 85939 86257 85956 86309
rect 86008 86257 86025 86309
rect 85939 86245 86025 86257
rect 85939 86193 85956 86245
rect 86008 86193 86025 86245
rect 85939 86188 86025 86193
rect 87027 86757 87113 86762
rect 87027 86705 87044 86757
rect 87096 86705 87113 86757
rect 87027 86693 87113 86705
rect 87027 86641 87044 86693
rect 87096 86641 87113 86693
rect 87027 86629 87113 86641
rect 87027 86577 87044 86629
rect 87096 86577 87113 86629
rect 87027 86565 87113 86577
rect 87027 86513 87044 86565
rect 87096 86513 87113 86565
rect 87027 86501 87113 86513
rect 87027 86449 87044 86501
rect 87096 86449 87113 86501
rect 87027 86437 87113 86449
rect 87027 86385 87044 86437
rect 87096 86385 87113 86437
rect 87027 86373 87113 86385
rect 87027 86321 87044 86373
rect 87096 86321 87113 86373
rect 87027 86309 87113 86321
rect 87027 86257 87044 86309
rect 87096 86257 87113 86309
rect 87027 86245 87113 86257
rect 87027 86193 87044 86245
rect 87096 86193 87113 86245
rect 87027 86188 87113 86193
rect 88115 86757 88201 86762
rect 88115 86705 88132 86757
rect 88184 86705 88201 86757
rect 88115 86693 88201 86705
rect 88115 86641 88132 86693
rect 88184 86641 88201 86693
rect 88115 86629 88201 86641
rect 88115 86577 88132 86629
rect 88184 86577 88201 86629
rect 88115 86565 88201 86577
rect 88115 86513 88132 86565
rect 88184 86513 88201 86565
rect 88115 86501 88201 86513
rect 88115 86449 88132 86501
rect 88184 86449 88201 86501
rect 88115 86437 88201 86449
rect 88115 86385 88132 86437
rect 88184 86385 88201 86437
rect 88115 86373 88201 86385
rect 88115 86321 88132 86373
rect 88184 86321 88201 86373
rect 88115 86309 88201 86321
rect 88115 86257 88132 86309
rect 88184 86257 88201 86309
rect 88115 86245 88201 86257
rect 88115 86193 88132 86245
rect 88184 86193 88201 86245
rect 88115 86188 88201 86193
rect 74514 84760 74600 84765
rect 74514 84708 74531 84760
rect 74583 84708 74600 84760
rect 74514 84696 74600 84708
rect 74514 84644 74531 84696
rect 74583 84644 74600 84696
rect 74514 84632 74600 84644
rect 74514 84580 74531 84632
rect 74583 84580 74600 84632
rect 74514 84568 74600 84580
rect 74514 84516 74531 84568
rect 74583 84516 74600 84568
rect 74514 84504 74600 84516
rect 74514 84452 74531 84504
rect 74583 84452 74600 84504
rect 74514 84440 74600 84452
rect 74514 84388 74531 84440
rect 74583 84388 74600 84440
rect 74514 84376 74600 84388
rect 74514 84324 74531 84376
rect 74583 84324 74600 84376
rect 74514 84312 74600 84324
rect 74514 84260 74531 84312
rect 74583 84260 74600 84312
rect 74514 84248 74600 84260
rect 74514 84196 74531 84248
rect 74583 84196 74600 84248
rect 74514 84191 74600 84196
rect 75602 84760 75688 84765
rect 75602 84708 75619 84760
rect 75671 84708 75688 84760
rect 75602 84696 75688 84708
rect 75602 84644 75619 84696
rect 75671 84644 75688 84696
rect 75602 84632 75688 84644
rect 75602 84580 75619 84632
rect 75671 84580 75688 84632
rect 75602 84568 75688 84580
rect 75602 84516 75619 84568
rect 75671 84516 75688 84568
rect 75602 84504 75688 84516
rect 75602 84452 75619 84504
rect 75671 84452 75688 84504
rect 75602 84440 75688 84452
rect 75602 84388 75619 84440
rect 75671 84388 75688 84440
rect 75602 84376 75688 84388
rect 75602 84324 75619 84376
rect 75671 84324 75688 84376
rect 75602 84312 75688 84324
rect 75602 84260 75619 84312
rect 75671 84260 75688 84312
rect 75602 84248 75688 84260
rect 75602 84196 75619 84248
rect 75671 84196 75688 84248
rect 75602 84191 75688 84196
rect 76690 84760 76776 84765
rect 76690 84708 76707 84760
rect 76759 84708 76776 84760
rect 76690 84696 76776 84708
rect 76690 84644 76707 84696
rect 76759 84644 76776 84696
rect 76690 84632 76776 84644
rect 76690 84580 76707 84632
rect 76759 84580 76776 84632
rect 76690 84568 76776 84580
rect 76690 84516 76707 84568
rect 76759 84516 76776 84568
rect 76690 84504 76776 84516
rect 76690 84452 76707 84504
rect 76759 84452 76776 84504
rect 76690 84440 76776 84452
rect 76690 84388 76707 84440
rect 76759 84388 76776 84440
rect 76690 84376 76776 84388
rect 76690 84324 76707 84376
rect 76759 84324 76776 84376
rect 76690 84312 76776 84324
rect 76690 84260 76707 84312
rect 76759 84260 76776 84312
rect 76690 84248 76776 84260
rect 76690 84196 76707 84248
rect 76759 84196 76776 84248
rect 76690 84191 76776 84196
rect 77778 84760 77864 84765
rect 77778 84708 77795 84760
rect 77847 84708 77864 84760
rect 77778 84696 77864 84708
rect 77778 84644 77795 84696
rect 77847 84644 77864 84696
rect 77778 84632 77864 84644
rect 77778 84580 77795 84632
rect 77847 84580 77864 84632
rect 77778 84568 77864 84580
rect 77778 84516 77795 84568
rect 77847 84516 77864 84568
rect 77778 84504 77864 84516
rect 77778 84452 77795 84504
rect 77847 84452 77864 84504
rect 77778 84440 77864 84452
rect 77778 84388 77795 84440
rect 77847 84388 77864 84440
rect 77778 84376 77864 84388
rect 77778 84324 77795 84376
rect 77847 84324 77864 84376
rect 77778 84312 77864 84324
rect 77778 84260 77795 84312
rect 77847 84260 77864 84312
rect 77778 84248 77864 84260
rect 77778 84196 77795 84248
rect 77847 84196 77864 84248
rect 77778 84191 77864 84196
rect 78866 84760 78952 84765
rect 78866 84708 78883 84760
rect 78935 84708 78952 84760
rect 78866 84696 78952 84708
rect 78866 84644 78883 84696
rect 78935 84644 78952 84696
rect 78866 84632 78952 84644
rect 78866 84580 78883 84632
rect 78935 84580 78952 84632
rect 78866 84568 78952 84580
rect 78866 84516 78883 84568
rect 78935 84516 78952 84568
rect 78866 84504 78952 84516
rect 78866 84452 78883 84504
rect 78935 84452 78952 84504
rect 78866 84440 78952 84452
rect 78866 84388 78883 84440
rect 78935 84388 78952 84440
rect 78866 84376 78952 84388
rect 78866 84324 78883 84376
rect 78935 84324 78952 84376
rect 78866 84312 78952 84324
rect 78866 84260 78883 84312
rect 78935 84260 78952 84312
rect 78866 84248 78952 84260
rect 78866 84196 78883 84248
rect 78935 84196 78952 84248
rect 78866 84191 78952 84196
rect 79954 84760 80040 84765
rect 79954 84708 79971 84760
rect 80023 84708 80040 84760
rect 79954 84696 80040 84708
rect 79954 84644 79971 84696
rect 80023 84644 80040 84696
rect 79954 84632 80040 84644
rect 79954 84580 79971 84632
rect 80023 84580 80040 84632
rect 79954 84568 80040 84580
rect 79954 84516 79971 84568
rect 80023 84516 80040 84568
rect 79954 84504 80040 84516
rect 79954 84452 79971 84504
rect 80023 84452 80040 84504
rect 79954 84440 80040 84452
rect 79954 84388 79971 84440
rect 80023 84388 80040 84440
rect 79954 84376 80040 84388
rect 79954 84324 79971 84376
rect 80023 84324 80040 84376
rect 79954 84312 80040 84324
rect 79954 84260 79971 84312
rect 80023 84260 80040 84312
rect 79954 84248 80040 84260
rect 79954 84196 79971 84248
rect 80023 84196 80040 84248
rect 79954 84191 80040 84196
rect 81042 84760 81128 84765
rect 81042 84708 81059 84760
rect 81111 84708 81128 84760
rect 81042 84696 81128 84708
rect 81042 84644 81059 84696
rect 81111 84644 81128 84696
rect 81042 84632 81128 84644
rect 81042 84580 81059 84632
rect 81111 84580 81128 84632
rect 81042 84568 81128 84580
rect 81042 84516 81059 84568
rect 81111 84516 81128 84568
rect 81042 84504 81128 84516
rect 81042 84452 81059 84504
rect 81111 84452 81128 84504
rect 81042 84440 81128 84452
rect 81042 84388 81059 84440
rect 81111 84388 81128 84440
rect 81042 84376 81128 84388
rect 81042 84324 81059 84376
rect 81111 84324 81128 84376
rect 81042 84312 81128 84324
rect 81042 84260 81059 84312
rect 81111 84260 81128 84312
rect 81042 84248 81128 84260
rect 81042 84196 81059 84248
rect 81111 84196 81128 84248
rect 81042 84191 81128 84196
rect 82130 84760 82216 84765
rect 82130 84708 82147 84760
rect 82199 84708 82216 84760
rect 82130 84696 82216 84708
rect 82130 84644 82147 84696
rect 82199 84644 82216 84696
rect 82130 84632 82216 84644
rect 82130 84580 82147 84632
rect 82199 84580 82216 84632
rect 82130 84568 82216 84580
rect 82130 84516 82147 84568
rect 82199 84516 82216 84568
rect 82130 84504 82216 84516
rect 82130 84452 82147 84504
rect 82199 84452 82216 84504
rect 82130 84440 82216 84452
rect 82130 84388 82147 84440
rect 82199 84388 82216 84440
rect 82130 84376 82216 84388
rect 82130 84324 82147 84376
rect 82199 84324 82216 84376
rect 82130 84312 82216 84324
rect 82130 84260 82147 84312
rect 82199 84260 82216 84312
rect 82130 84248 82216 84260
rect 82130 84196 82147 84248
rect 82199 84196 82216 84248
rect 82130 84191 82216 84196
rect 83218 84760 83304 84765
rect 83218 84708 83235 84760
rect 83287 84708 83304 84760
rect 83218 84696 83304 84708
rect 83218 84644 83235 84696
rect 83287 84644 83304 84696
rect 83218 84632 83304 84644
rect 83218 84580 83235 84632
rect 83287 84580 83304 84632
rect 83218 84568 83304 84580
rect 83218 84516 83235 84568
rect 83287 84516 83304 84568
rect 83218 84504 83304 84516
rect 83218 84452 83235 84504
rect 83287 84452 83304 84504
rect 83218 84440 83304 84452
rect 83218 84388 83235 84440
rect 83287 84388 83304 84440
rect 83218 84376 83304 84388
rect 83218 84324 83235 84376
rect 83287 84324 83304 84376
rect 83218 84312 83304 84324
rect 83218 84260 83235 84312
rect 83287 84260 83304 84312
rect 83218 84248 83304 84260
rect 83218 84196 83235 84248
rect 83287 84196 83304 84248
rect 83218 84191 83304 84196
rect 84306 84760 84392 84765
rect 84306 84708 84323 84760
rect 84375 84708 84392 84760
rect 84306 84696 84392 84708
rect 84306 84644 84323 84696
rect 84375 84644 84392 84696
rect 84306 84632 84392 84644
rect 84306 84580 84323 84632
rect 84375 84580 84392 84632
rect 84306 84568 84392 84580
rect 84306 84516 84323 84568
rect 84375 84516 84392 84568
rect 84306 84504 84392 84516
rect 84306 84452 84323 84504
rect 84375 84452 84392 84504
rect 84306 84440 84392 84452
rect 84306 84388 84323 84440
rect 84375 84388 84392 84440
rect 84306 84376 84392 84388
rect 84306 84324 84323 84376
rect 84375 84324 84392 84376
rect 84306 84312 84392 84324
rect 84306 84260 84323 84312
rect 84375 84260 84392 84312
rect 84306 84248 84392 84260
rect 84306 84196 84323 84248
rect 84375 84196 84392 84248
rect 84306 84191 84392 84196
rect 85394 84760 85480 84765
rect 85394 84708 85411 84760
rect 85463 84708 85480 84760
rect 85394 84696 85480 84708
rect 85394 84644 85411 84696
rect 85463 84644 85480 84696
rect 85394 84632 85480 84644
rect 85394 84580 85411 84632
rect 85463 84580 85480 84632
rect 85394 84568 85480 84580
rect 85394 84516 85411 84568
rect 85463 84516 85480 84568
rect 85394 84504 85480 84516
rect 85394 84452 85411 84504
rect 85463 84452 85480 84504
rect 85394 84440 85480 84452
rect 85394 84388 85411 84440
rect 85463 84388 85480 84440
rect 85394 84376 85480 84388
rect 85394 84324 85411 84376
rect 85463 84324 85480 84376
rect 85394 84312 85480 84324
rect 85394 84260 85411 84312
rect 85463 84260 85480 84312
rect 85394 84248 85480 84260
rect 85394 84196 85411 84248
rect 85463 84196 85480 84248
rect 85394 84191 85480 84196
rect 86482 84760 86568 84765
rect 86482 84708 86499 84760
rect 86551 84708 86568 84760
rect 86482 84696 86568 84708
rect 86482 84644 86499 84696
rect 86551 84644 86568 84696
rect 86482 84632 86568 84644
rect 86482 84580 86499 84632
rect 86551 84580 86568 84632
rect 86482 84568 86568 84580
rect 86482 84516 86499 84568
rect 86551 84516 86568 84568
rect 86482 84504 86568 84516
rect 86482 84452 86499 84504
rect 86551 84452 86568 84504
rect 86482 84440 86568 84452
rect 86482 84388 86499 84440
rect 86551 84388 86568 84440
rect 86482 84376 86568 84388
rect 86482 84324 86499 84376
rect 86551 84324 86568 84376
rect 86482 84312 86568 84324
rect 86482 84260 86499 84312
rect 86551 84260 86568 84312
rect 86482 84248 86568 84260
rect 86482 84196 86499 84248
rect 86551 84196 86568 84248
rect 86482 84191 86568 84196
rect 87570 84760 87656 84765
rect 87570 84708 87587 84760
rect 87639 84708 87656 84760
rect 87570 84696 87656 84708
rect 87570 84644 87587 84696
rect 87639 84644 87656 84696
rect 87570 84632 87656 84644
rect 87570 84580 87587 84632
rect 87639 84580 87656 84632
rect 87570 84568 87656 84580
rect 87570 84516 87587 84568
rect 87639 84516 87656 84568
rect 87570 84504 87656 84516
rect 87570 84452 87587 84504
rect 87639 84452 87656 84504
rect 87570 84440 87656 84452
rect 87570 84388 87587 84440
rect 87639 84388 87656 84440
rect 87570 84376 87656 84388
rect 87570 84324 87587 84376
rect 87639 84324 87656 84376
rect 87570 84312 87656 84324
rect 87570 84260 87587 84312
rect 87639 84260 87656 84312
rect 87570 84248 87656 84260
rect 87570 84196 87587 84248
rect 87639 84196 87656 84248
rect 87570 84191 87656 84196
rect 88658 84760 88744 84765
rect 88658 84708 88675 84760
rect 88727 84708 88744 84760
rect 88658 84696 88744 84708
rect 88658 84644 88675 84696
rect 88727 84644 88744 84696
rect 88658 84632 88744 84644
rect 88658 84580 88675 84632
rect 88727 84580 88744 84632
rect 88658 84568 88744 84580
rect 88658 84516 88675 84568
rect 88727 84516 88744 84568
rect 88658 84504 88744 84516
rect 88658 84452 88675 84504
rect 88727 84452 88744 84504
rect 88658 84440 88744 84452
rect 88658 84388 88675 84440
rect 88727 84388 88744 84440
rect 88658 84376 88744 84388
rect 88658 84324 88675 84376
rect 88727 84324 88744 84376
rect 88658 84312 88744 84324
rect 88658 84260 88675 84312
rect 88727 84260 88744 84312
rect 88658 84248 88744 84260
rect 88658 84196 88675 84248
rect 88727 84196 88744 84248
rect 88658 84191 88744 84196
rect 75059 82757 75145 82762
rect 75059 82705 75076 82757
rect 75128 82705 75145 82757
rect 75059 82693 75145 82705
rect 75059 82641 75076 82693
rect 75128 82641 75145 82693
rect 75059 82629 75145 82641
rect 75059 82577 75076 82629
rect 75128 82577 75145 82629
rect 75059 82565 75145 82577
rect 75059 82513 75076 82565
rect 75128 82513 75145 82565
rect 75059 82501 75145 82513
rect 75059 82449 75076 82501
rect 75128 82449 75145 82501
rect 75059 82437 75145 82449
rect 75059 82385 75076 82437
rect 75128 82385 75145 82437
rect 75059 82373 75145 82385
rect 75059 82321 75076 82373
rect 75128 82321 75145 82373
rect 75059 82309 75145 82321
rect 75059 82257 75076 82309
rect 75128 82257 75145 82309
rect 75059 82245 75145 82257
rect 75059 82193 75076 82245
rect 75128 82193 75145 82245
rect 75059 82188 75145 82193
rect 76147 82757 76233 82762
rect 76147 82705 76164 82757
rect 76216 82705 76233 82757
rect 76147 82693 76233 82705
rect 76147 82641 76164 82693
rect 76216 82641 76233 82693
rect 76147 82629 76233 82641
rect 76147 82577 76164 82629
rect 76216 82577 76233 82629
rect 76147 82565 76233 82577
rect 76147 82513 76164 82565
rect 76216 82513 76233 82565
rect 76147 82501 76233 82513
rect 76147 82449 76164 82501
rect 76216 82449 76233 82501
rect 76147 82437 76233 82449
rect 76147 82385 76164 82437
rect 76216 82385 76233 82437
rect 76147 82373 76233 82385
rect 76147 82321 76164 82373
rect 76216 82321 76233 82373
rect 76147 82309 76233 82321
rect 76147 82257 76164 82309
rect 76216 82257 76233 82309
rect 76147 82245 76233 82257
rect 76147 82193 76164 82245
rect 76216 82193 76233 82245
rect 76147 82188 76233 82193
rect 77235 82757 77321 82762
rect 77235 82705 77252 82757
rect 77304 82705 77321 82757
rect 77235 82693 77321 82705
rect 77235 82641 77252 82693
rect 77304 82641 77321 82693
rect 77235 82629 77321 82641
rect 77235 82577 77252 82629
rect 77304 82577 77321 82629
rect 77235 82565 77321 82577
rect 77235 82513 77252 82565
rect 77304 82513 77321 82565
rect 77235 82501 77321 82513
rect 77235 82449 77252 82501
rect 77304 82449 77321 82501
rect 77235 82437 77321 82449
rect 77235 82385 77252 82437
rect 77304 82385 77321 82437
rect 77235 82373 77321 82385
rect 77235 82321 77252 82373
rect 77304 82321 77321 82373
rect 77235 82309 77321 82321
rect 77235 82257 77252 82309
rect 77304 82257 77321 82309
rect 77235 82245 77321 82257
rect 77235 82193 77252 82245
rect 77304 82193 77321 82245
rect 77235 82188 77321 82193
rect 78323 82757 78409 82762
rect 78323 82705 78340 82757
rect 78392 82705 78409 82757
rect 78323 82693 78409 82705
rect 78323 82641 78340 82693
rect 78392 82641 78409 82693
rect 78323 82629 78409 82641
rect 78323 82577 78340 82629
rect 78392 82577 78409 82629
rect 78323 82565 78409 82577
rect 78323 82513 78340 82565
rect 78392 82513 78409 82565
rect 78323 82501 78409 82513
rect 78323 82449 78340 82501
rect 78392 82449 78409 82501
rect 78323 82437 78409 82449
rect 78323 82385 78340 82437
rect 78392 82385 78409 82437
rect 78323 82373 78409 82385
rect 78323 82321 78340 82373
rect 78392 82321 78409 82373
rect 78323 82309 78409 82321
rect 78323 82257 78340 82309
rect 78392 82257 78409 82309
rect 78323 82245 78409 82257
rect 78323 82193 78340 82245
rect 78392 82193 78409 82245
rect 78323 82188 78409 82193
rect 79411 82757 79497 82762
rect 79411 82705 79428 82757
rect 79480 82705 79497 82757
rect 79411 82693 79497 82705
rect 79411 82641 79428 82693
rect 79480 82641 79497 82693
rect 79411 82629 79497 82641
rect 79411 82577 79428 82629
rect 79480 82577 79497 82629
rect 79411 82565 79497 82577
rect 79411 82513 79428 82565
rect 79480 82513 79497 82565
rect 79411 82501 79497 82513
rect 79411 82449 79428 82501
rect 79480 82449 79497 82501
rect 79411 82437 79497 82449
rect 79411 82385 79428 82437
rect 79480 82385 79497 82437
rect 79411 82373 79497 82385
rect 79411 82321 79428 82373
rect 79480 82321 79497 82373
rect 79411 82309 79497 82321
rect 79411 82257 79428 82309
rect 79480 82257 79497 82309
rect 79411 82245 79497 82257
rect 79411 82193 79428 82245
rect 79480 82193 79497 82245
rect 79411 82188 79497 82193
rect 80499 82757 80585 82762
rect 80499 82705 80516 82757
rect 80568 82705 80585 82757
rect 80499 82693 80585 82705
rect 80499 82641 80516 82693
rect 80568 82641 80585 82693
rect 80499 82629 80585 82641
rect 80499 82577 80516 82629
rect 80568 82577 80585 82629
rect 80499 82565 80585 82577
rect 80499 82513 80516 82565
rect 80568 82513 80585 82565
rect 80499 82501 80585 82513
rect 80499 82449 80516 82501
rect 80568 82449 80585 82501
rect 80499 82437 80585 82449
rect 80499 82385 80516 82437
rect 80568 82385 80585 82437
rect 80499 82373 80585 82385
rect 80499 82321 80516 82373
rect 80568 82321 80585 82373
rect 80499 82309 80585 82321
rect 80499 82257 80516 82309
rect 80568 82257 80585 82309
rect 80499 82245 80585 82257
rect 80499 82193 80516 82245
rect 80568 82193 80585 82245
rect 80499 82188 80585 82193
rect 81587 82757 81673 82762
rect 81587 82705 81604 82757
rect 81656 82705 81673 82757
rect 81587 82693 81673 82705
rect 81587 82641 81604 82693
rect 81656 82641 81673 82693
rect 81587 82629 81673 82641
rect 81587 82577 81604 82629
rect 81656 82577 81673 82629
rect 81587 82565 81673 82577
rect 81587 82513 81604 82565
rect 81656 82513 81673 82565
rect 81587 82501 81673 82513
rect 81587 82449 81604 82501
rect 81656 82449 81673 82501
rect 81587 82437 81673 82449
rect 81587 82385 81604 82437
rect 81656 82385 81673 82437
rect 81587 82373 81673 82385
rect 81587 82321 81604 82373
rect 81656 82321 81673 82373
rect 81587 82309 81673 82321
rect 81587 82257 81604 82309
rect 81656 82257 81673 82309
rect 81587 82245 81673 82257
rect 81587 82193 81604 82245
rect 81656 82193 81673 82245
rect 81587 82188 81673 82193
rect 82675 82757 82761 82762
rect 82675 82705 82692 82757
rect 82744 82705 82761 82757
rect 82675 82693 82761 82705
rect 82675 82641 82692 82693
rect 82744 82641 82761 82693
rect 82675 82629 82761 82641
rect 82675 82577 82692 82629
rect 82744 82577 82761 82629
rect 82675 82565 82761 82577
rect 82675 82513 82692 82565
rect 82744 82513 82761 82565
rect 82675 82501 82761 82513
rect 82675 82449 82692 82501
rect 82744 82449 82761 82501
rect 82675 82437 82761 82449
rect 82675 82385 82692 82437
rect 82744 82385 82761 82437
rect 82675 82373 82761 82385
rect 82675 82321 82692 82373
rect 82744 82321 82761 82373
rect 82675 82309 82761 82321
rect 82675 82257 82692 82309
rect 82744 82257 82761 82309
rect 82675 82245 82761 82257
rect 82675 82193 82692 82245
rect 82744 82193 82761 82245
rect 82675 82188 82761 82193
rect 83763 82757 83849 82762
rect 83763 82705 83780 82757
rect 83832 82705 83849 82757
rect 83763 82693 83849 82705
rect 83763 82641 83780 82693
rect 83832 82641 83849 82693
rect 83763 82629 83849 82641
rect 83763 82577 83780 82629
rect 83832 82577 83849 82629
rect 83763 82565 83849 82577
rect 83763 82513 83780 82565
rect 83832 82513 83849 82565
rect 83763 82501 83849 82513
rect 83763 82449 83780 82501
rect 83832 82449 83849 82501
rect 83763 82437 83849 82449
rect 83763 82385 83780 82437
rect 83832 82385 83849 82437
rect 83763 82373 83849 82385
rect 83763 82321 83780 82373
rect 83832 82321 83849 82373
rect 83763 82309 83849 82321
rect 83763 82257 83780 82309
rect 83832 82257 83849 82309
rect 83763 82245 83849 82257
rect 83763 82193 83780 82245
rect 83832 82193 83849 82245
rect 83763 82188 83849 82193
rect 84851 82757 84937 82762
rect 84851 82705 84868 82757
rect 84920 82705 84937 82757
rect 84851 82693 84937 82705
rect 84851 82641 84868 82693
rect 84920 82641 84937 82693
rect 84851 82629 84937 82641
rect 84851 82577 84868 82629
rect 84920 82577 84937 82629
rect 84851 82565 84937 82577
rect 84851 82513 84868 82565
rect 84920 82513 84937 82565
rect 84851 82501 84937 82513
rect 84851 82449 84868 82501
rect 84920 82449 84937 82501
rect 84851 82437 84937 82449
rect 84851 82385 84868 82437
rect 84920 82385 84937 82437
rect 84851 82373 84937 82385
rect 84851 82321 84868 82373
rect 84920 82321 84937 82373
rect 84851 82309 84937 82321
rect 84851 82257 84868 82309
rect 84920 82257 84937 82309
rect 84851 82245 84937 82257
rect 84851 82193 84868 82245
rect 84920 82193 84937 82245
rect 84851 82188 84937 82193
rect 85939 82757 86025 82762
rect 85939 82705 85956 82757
rect 86008 82705 86025 82757
rect 85939 82693 86025 82705
rect 85939 82641 85956 82693
rect 86008 82641 86025 82693
rect 85939 82629 86025 82641
rect 85939 82577 85956 82629
rect 86008 82577 86025 82629
rect 85939 82565 86025 82577
rect 85939 82513 85956 82565
rect 86008 82513 86025 82565
rect 85939 82501 86025 82513
rect 85939 82449 85956 82501
rect 86008 82449 86025 82501
rect 85939 82437 86025 82449
rect 85939 82385 85956 82437
rect 86008 82385 86025 82437
rect 85939 82373 86025 82385
rect 85939 82321 85956 82373
rect 86008 82321 86025 82373
rect 85939 82309 86025 82321
rect 85939 82257 85956 82309
rect 86008 82257 86025 82309
rect 85939 82245 86025 82257
rect 85939 82193 85956 82245
rect 86008 82193 86025 82245
rect 85939 82188 86025 82193
rect 87027 82757 87113 82762
rect 87027 82705 87044 82757
rect 87096 82705 87113 82757
rect 87027 82693 87113 82705
rect 87027 82641 87044 82693
rect 87096 82641 87113 82693
rect 87027 82629 87113 82641
rect 87027 82577 87044 82629
rect 87096 82577 87113 82629
rect 87027 82565 87113 82577
rect 87027 82513 87044 82565
rect 87096 82513 87113 82565
rect 87027 82501 87113 82513
rect 87027 82449 87044 82501
rect 87096 82449 87113 82501
rect 87027 82437 87113 82449
rect 87027 82385 87044 82437
rect 87096 82385 87113 82437
rect 87027 82373 87113 82385
rect 87027 82321 87044 82373
rect 87096 82321 87113 82373
rect 87027 82309 87113 82321
rect 87027 82257 87044 82309
rect 87096 82257 87113 82309
rect 87027 82245 87113 82257
rect 87027 82193 87044 82245
rect 87096 82193 87113 82245
rect 87027 82188 87113 82193
rect 88115 82757 88201 82762
rect 88115 82705 88132 82757
rect 88184 82705 88201 82757
rect 88115 82693 88201 82705
rect 88115 82641 88132 82693
rect 88184 82641 88201 82693
rect 88115 82629 88201 82641
rect 88115 82577 88132 82629
rect 88184 82577 88201 82629
rect 88115 82565 88201 82577
rect 88115 82513 88132 82565
rect 88184 82513 88201 82565
rect 88115 82501 88201 82513
rect 88115 82449 88132 82501
rect 88184 82449 88201 82501
rect 88115 82437 88201 82449
rect 88115 82385 88132 82437
rect 88184 82385 88201 82437
rect 88115 82373 88201 82385
rect 88115 82321 88132 82373
rect 88184 82321 88201 82373
rect 88115 82309 88201 82321
rect 88115 82257 88132 82309
rect 88184 82257 88201 82309
rect 88115 82245 88201 82257
rect 88115 82193 88132 82245
rect 88184 82193 88201 82245
rect 88115 82188 88201 82193
rect 74514 80760 74600 80765
rect 74514 80708 74531 80760
rect 74583 80708 74600 80760
rect 74514 80696 74600 80708
rect 74514 80644 74531 80696
rect 74583 80644 74600 80696
rect 74514 80632 74600 80644
rect 74514 80580 74531 80632
rect 74583 80580 74600 80632
rect 74514 80568 74600 80580
rect 74514 80516 74531 80568
rect 74583 80516 74600 80568
rect 74514 80504 74600 80516
rect 74514 80452 74531 80504
rect 74583 80452 74600 80504
rect 74514 80440 74600 80452
rect 74514 80388 74531 80440
rect 74583 80388 74600 80440
rect 74514 80376 74600 80388
rect 74514 80324 74531 80376
rect 74583 80324 74600 80376
rect 74514 80312 74600 80324
rect 74514 80260 74531 80312
rect 74583 80260 74600 80312
rect 74514 80248 74600 80260
rect 74514 80196 74531 80248
rect 74583 80196 74600 80248
rect 74514 80191 74600 80196
rect 75602 80760 75688 80765
rect 75602 80708 75619 80760
rect 75671 80708 75688 80760
rect 75602 80696 75688 80708
rect 75602 80644 75619 80696
rect 75671 80644 75688 80696
rect 75602 80632 75688 80644
rect 75602 80580 75619 80632
rect 75671 80580 75688 80632
rect 75602 80568 75688 80580
rect 75602 80516 75619 80568
rect 75671 80516 75688 80568
rect 75602 80504 75688 80516
rect 75602 80452 75619 80504
rect 75671 80452 75688 80504
rect 75602 80440 75688 80452
rect 75602 80388 75619 80440
rect 75671 80388 75688 80440
rect 75602 80376 75688 80388
rect 75602 80324 75619 80376
rect 75671 80324 75688 80376
rect 75602 80312 75688 80324
rect 75602 80260 75619 80312
rect 75671 80260 75688 80312
rect 75602 80248 75688 80260
rect 75602 80196 75619 80248
rect 75671 80196 75688 80248
rect 75602 80191 75688 80196
rect 76690 80760 76776 80765
rect 76690 80708 76707 80760
rect 76759 80708 76776 80760
rect 76690 80696 76776 80708
rect 76690 80644 76707 80696
rect 76759 80644 76776 80696
rect 76690 80632 76776 80644
rect 76690 80580 76707 80632
rect 76759 80580 76776 80632
rect 76690 80568 76776 80580
rect 76690 80516 76707 80568
rect 76759 80516 76776 80568
rect 76690 80504 76776 80516
rect 76690 80452 76707 80504
rect 76759 80452 76776 80504
rect 76690 80440 76776 80452
rect 76690 80388 76707 80440
rect 76759 80388 76776 80440
rect 76690 80376 76776 80388
rect 76690 80324 76707 80376
rect 76759 80324 76776 80376
rect 76690 80312 76776 80324
rect 76690 80260 76707 80312
rect 76759 80260 76776 80312
rect 76690 80248 76776 80260
rect 76690 80196 76707 80248
rect 76759 80196 76776 80248
rect 76690 80191 76776 80196
rect 77778 80760 77864 80765
rect 77778 80708 77795 80760
rect 77847 80708 77864 80760
rect 77778 80696 77864 80708
rect 77778 80644 77795 80696
rect 77847 80644 77864 80696
rect 77778 80632 77864 80644
rect 77778 80580 77795 80632
rect 77847 80580 77864 80632
rect 77778 80568 77864 80580
rect 77778 80516 77795 80568
rect 77847 80516 77864 80568
rect 77778 80504 77864 80516
rect 77778 80452 77795 80504
rect 77847 80452 77864 80504
rect 77778 80440 77864 80452
rect 77778 80388 77795 80440
rect 77847 80388 77864 80440
rect 77778 80376 77864 80388
rect 77778 80324 77795 80376
rect 77847 80324 77864 80376
rect 77778 80312 77864 80324
rect 77778 80260 77795 80312
rect 77847 80260 77864 80312
rect 77778 80248 77864 80260
rect 77778 80196 77795 80248
rect 77847 80196 77864 80248
rect 77778 80191 77864 80196
rect 78866 80760 78952 80765
rect 78866 80708 78883 80760
rect 78935 80708 78952 80760
rect 78866 80696 78952 80708
rect 78866 80644 78883 80696
rect 78935 80644 78952 80696
rect 78866 80632 78952 80644
rect 78866 80580 78883 80632
rect 78935 80580 78952 80632
rect 78866 80568 78952 80580
rect 78866 80516 78883 80568
rect 78935 80516 78952 80568
rect 78866 80504 78952 80516
rect 78866 80452 78883 80504
rect 78935 80452 78952 80504
rect 78866 80440 78952 80452
rect 78866 80388 78883 80440
rect 78935 80388 78952 80440
rect 78866 80376 78952 80388
rect 78866 80324 78883 80376
rect 78935 80324 78952 80376
rect 78866 80312 78952 80324
rect 78866 80260 78883 80312
rect 78935 80260 78952 80312
rect 78866 80248 78952 80260
rect 78866 80196 78883 80248
rect 78935 80196 78952 80248
rect 78866 80191 78952 80196
rect 79954 80760 80040 80765
rect 79954 80708 79971 80760
rect 80023 80708 80040 80760
rect 79954 80696 80040 80708
rect 79954 80644 79971 80696
rect 80023 80644 80040 80696
rect 79954 80632 80040 80644
rect 79954 80580 79971 80632
rect 80023 80580 80040 80632
rect 79954 80568 80040 80580
rect 79954 80516 79971 80568
rect 80023 80516 80040 80568
rect 79954 80504 80040 80516
rect 79954 80452 79971 80504
rect 80023 80452 80040 80504
rect 79954 80440 80040 80452
rect 79954 80388 79971 80440
rect 80023 80388 80040 80440
rect 79954 80376 80040 80388
rect 79954 80324 79971 80376
rect 80023 80324 80040 80376
rect 79954 80312 80040 80324
rect 79954 80260 79971 80312
rect 80023 80260 80040 80312
rect 79954 80248 80040 80260
rect 79954 80196 79971 80248
rect 80023 80196 80040 80248
rect 79954 80191 80040 80196
rect 81042 80760 81128 80765
rect 81042 80708 81059 80760
rect 81111 80708 81128 80760
rect 81042 80696 81128 80708
rect 81042 80644 81059 80696
rect 81111 80644 81128 80696
rect 81042 80632 81128 80644
rect 81042 80580 81059 80632
rect 81111 80580 81128 80632
rect 81042 80568 81128 80580
rect 81042 80516 81059 80568
rect 81111 80516 81128 80568
rect 81042 80504 81128 80516
rect 81042 80452 81059 80504
rect 81111 80452 81128 80504
rect 81042 80440 81128 80452
rect 81042 80388 81059 80440
rect 81111 80388 81128 80440
rect 81042 80376 81128 80388
rect 81042 80324 81059 80376
rect 81111 80324 81128 80376
rect 81042 80312 81128 80324
rect 81042 80260 81059 80312
rect 81111 80260 81128 80312
rect 81042 80248 81128 80260
rect 81042 80196 81059 80248
rect 81111 80196 81128 80248
rect 81042 80191 81128 80196
rect 82130 80760 82216 80765
rect 82130 80708 82147 80760
rect 82199 80708 82216 80760
rect 82130 80696 82216 80708
rect 82130 80644 82147 80696
rect 82199 80644 82216 80696
rect 82130 80632 82216 80644
rect 82130 80580 82147 80632
rect 82199 80580 82216 80632
rect 82130 80568 82216 80580
rect 82130 80516 82147 80568
rect 82199 80516 82216 80568
rect 82130 80504 82216 80516
rect 82130 80452 82147 80504
rect 82199 80452 82216 80504
rect 82130 80440 82216 80452
rect 82130 80388 82147 80440
rect 82199 80388 82216 80440
rect 82130 80376 82216 80388
rect 82130 80324 82147 80376
rect 82199 80324 82216 80376
rect 82130 80312 82216 80324
rect 82130 80260 82147 80312
rect 82199 80260 82216 80312
rect 82130 80248 82216 80260
rect 82130 80196 82147 80248
rect 82199 80196 82216 80248
rect 82130 80191 82216 80196
rect 83218 80760 83304 80765
rect 83218 80708 83235 80760
rect 83287 80708 83304 80760
rect 83218 80696 83304 80708
rect 83218 80644 83235 80696
rect 83287 80644 83304 80696
rect 83218 80632 83304 80644
rect 83218 80580 83235 80632
rect 83287 80580 83304 80632
rect 83218 80568 83304 80580
rect 83218 80516 83235 80568
rect 83287 80516 83304 80568
rect 83218 80504 83304 80516
rect 83218 80452 83235 80504
rect 83287 80452 83304 80504
rect 83218 80440 83304 80452
rect 83218 80388 83235 80440
rect 83287 80388 83304 80440
rect 83218 80376 83304 80388
rect 83218 80324 83235 80376
rect 83287 80324 83304 80376
rect 83218 80312 83304 80324
rect 83218 80260 83235 80312
rect 83287 80260 83304 80312
rect 83218 80248 83304 80260
rect 83218 80196 83235 80248
rect 83287 80196 83304 80248
rect 83218 80191 83304 80196
rect 84306 80760 84392 80765
rect 84306 80708 84323 80760
rect 84375 80708 84392 80760
rect 84306 80696 84392 80708
rect 84306 80644 84323 80696
rect 84375 80644 84392 80696
rect 84306 80632 84392 80644
rect 84306 80580 84323 80632
rect 84375 80580 84392 80632
rect 84306 80568 84392 80580
rect 84306 80516 84323 80568
rect 84375 80516 84392 80568
rect 84306 80504 84392 80516
rect 84306 80452 84323 80504
rect 84375 80452 84392 80504
rect 84306 80440 84392 80452
rect 84306 80388 84323 80440
rect 84375 80388 84392 80440
rect 84306 80376 84392 80388
rect 84306 80324 84323 80376
rect 84375 80324 84392 80376
rect 84306 80312 84392 80324
rect 84306 80260 84323 80312
rect 84375 80260 84392 80312
rect 84306 80248 84392 80260
rect 84306 80196 84323 80248
rect 84375 80196 84392 80248
rect 84306 80191 84392 80196
rect 85394 80760 85480 80765
rect 85394 80708 85411 80760
rect 85463 80708 85480 80760
rect 85394 80696 85480 80708
rect 85394 80644 85411 80696
rect 85463 80644 85480 80696
rect 85394 80632 85480 80644
rect 85394 80580 85411 80632
rect 85463 80580 85480 80632
rect 85394 80568 85480 80580
rect 85394 80516 85411 80568
rect 85463 80516 85480 80568
rect 85394 80504 85480 80516
rect 85394 80452 85411 80504
rect 85463 80452 85480 80504
rect 85394 80440 85480 80452
rect 85394 80388 85411 80440
rect 85463 80388 85480 80440
rect 85394 80376 85480 80388
rect 85394 80324 85411 80376
rect 85463 80324 85480 80376
rect 85394 80312 85480 80324
rect 85394 80260 85411 80312
rect 85463 80260 85480 80312
rect 85394 80248 85480 80260
rect 85394 80196 85411 80248
rect 85463 80196 85480 80248
rect 85394 80191 85480 80196
rect 86482 80760 86568 80765
rect 86482 80708 86499 80760
rect 86551 80708 86568 80760
rect 86482 80696 86568 80708
rect 86482 80644 86499 80696
rect 86551 80644 86568 80696
rect 86482 80632 86568 80644
rect 86482 80580 86499 80632
rect 86551 80580 86568 80632
rect 86482 80568 86568 80580
rect 86482 80516 86499 80568
rect 86551 80516 86568 80568
rect 86482 80504 86568 80516
rect 86482 80452 86499 80504
rect 86551 80452 86568 80504
rect 86482 80440 86568 80452
rect 86482 80388 86499 80440
rect 86551 80388 86568 80440
rect 86482 80376 86568 80388
rect 86482 80324 86499 80376
rect 86551 80324 86568 80376
rect 86482 80312 86568 80324
rect 86482 80260 86499 80312
rect 86551 80260 86568 80312
rect 86482 80248 86568 80260
rect 86482 80196 86499 80248
rect 86551 80196 86568 80248
rect 86482 80191 86568 80196
rect 87570 80760 87656 80765
rect 87570 80708 87587 80760
rect 87639 80708 87656 80760
rect 87570 80696 87656 80708
rect 87570 80644 87587 80696
rect 87639 80644 87656 80696
rect 87570 80632 87656 80644
rect 87570 80580 87587 80632
rect 87639 80580 87656 80632
rect 87570 80568 87656 80580
rect 87570 80516 87587 80568
rect 87639 80516 87656 80568
rect 87570 80504 87656 80516
rect 87570 80452 87587 80504
rect 87639 80452 87656 80504
rect 87570 80440 87656 80452
rect 87570 80388 87587 80440
rect 87639 80388 87656 80440
rect 87570 80376 87656 80388
rect 87570 80324 87587 80376
rect 87639 80324 87656 80376
rect 87570 80312 87656 80324
rect 87570 80260 87587 80312
rect 87639 80260 87656 80312
rect 87570 80248 87656 80260
rect 87570 80196 87587 80248
rect 87639 80196 87656 80248
rect 87570 80191 87656 80196
rect 88658 80760 88744 80765
rect 88658 80708 88675 80760
rect 88727 80708 88744 80760
rect 88658 80696 88744 80708
rect 88658 80644 88675 80696
rect 88727 80644 88744 80696
rect 88658 80632 88744 80644
rect 88658 80580 88675 80632
rect 88727 80580 88744 80632
rect 88658 80568 88744 80580
rect 88658 80516 88675 80568
rect 88727 80516 88744 80568
rect 88658 80504 88744 80516
rect 88658 80452 88675 80504
rect 88727 80452 88744 80504
rect 88658 80440 88744 80452
rect 88658 80388 88675 80440
rect 88727 80388 88744 80440
rect 88658 80376 88744 80388
rect 88658 80324 88675 80376
rect 88727 80324 88744 80376
rect 88658 80312 88744 80324
rect 88658 80260 88675 80312
rect 88727 80260 88744 80312
rect 88658 80248 88744 80260
rect 88658 80196 88675 80248
rect 88727 80196 88744 80248
rect 88658 80191 88744 80196
rect 75059 78757 75145 78762
rect 75059 78705 75076 78757
rect 75128 78705 75145 78757
rect 75059 78693 75145 78705
rect 75059 78641 75076 78693
rect 75128 78641 75145 78693
rect 75059 78629 75145 78641
rect 75059 78577 75076 78629
rect 75128 78577 75145 78629
rect 75059 78565 75145 78577
rect 75059 78513 75076 78565
rect 75128 78513 75145 78565
rect 75059 78501 75145 78513
rect 75059 78449 75076 78501
rect 75128 78449 75145 78501
rect 75059 78437 75145 78449
rect 75059 78385 75076 78437
rect 75128 78385 75145 78437
rect 75059 78373 75145 78385
rect 75059 78321 75076 78373
rect 75128 78321 75145 78373
rect 75059 78309 75145 78321
rect 75059 78257 75076 78309
rect 75128 78257 75145 78309
rect 75059 78245 75145 78257
rect 75059 78193 75076 78245
rect 75128 78193 75145 78245
rect 75059 78188 75145 78193
rect 76147 78757 76233 78762
rect 76147 78705 76164 78757
rect 76216 78705 76233 78757
rect 76147 78693 76233 78705
rect 76147 78641 76164 78693
rect 76216 78641 76233 78693
rect 76147 78629 76233 78641
rect 76147 78577 76164 78629
rect 76216 78577 76233 78629
rect 76147 78565 76233 78577
rect 76147 78513 76164 78565
rect 76216 78513 76233 78565
rect 76147 78501 76233 78513
rect 76147 78449 76164 78501
rect 76216 78449 76233 78501
rect 76147 78437 76233 78449
rect 76147 78385 76164 78437
rect 76216 78385 76233 78437
rect 76147 78373 76233 78385
rect 76147 78321 76164 78373
rect 76216 78321 76233 78373
rect 76147 78309 76233 78321
rect 76147 78257 76164 78309
rect 76216 78257 76233 78309
rect 76147 78245 76233 78257
rect 76147 78193 76164 78245
rect 76216 78193 76233 78245
rect 76147 78188 76233 78193
rect 77235 78757 77321 78762
rect 77235 78705 77252 78757
rect 77304 78705 77321 78757
rect 77235 78693 77321 78705
rect 77235 78641 77252 78693
rect 77304 78641 77321 78693
rect 77235 78629 77321 78641
rect 77235 78577 77252 78629
rect 77304 78577 77321 78629
rect 77235 78565 77321 78577
rect 77235 78513 77252 78565
rect 77304 78513 77321 78565
rect 77235 78501 77321 78513
rect 77235 78449 77252 78501
rect 77304 78449 77321 78501
rect 77235 78437 77321 78449
rect 77235 78385 77252 78437
rect 77304 78385 77321 78437
rect 77235 78373 77321 78385
rect 77235 78321 77252 78373
rect 77304 78321 77321 78373
rect 77235 78309 77321 78321
rect 77235 78257 77252 78309
rect 77304 78257 77321 78309
rect 77235 78245 77321 78257
rect 77235 78193 77252 78245
rect 77304 78193 77321 78245
rect 77235 78188 77321 78193
rect 78323 78757 78409 78762
rect 78323 78705 78340 78757
rect 78392 78705 78409 78757
rect 78323 78693 78409 78705
rect 78323 78641 78340 78693
rect 78392 78641 78409 78693
rect 78323 78629 78409 78641
rect 78323 78577 78340 78629
rect 78392 78577 78409 78629
rect 78323 78565 78409 78577
rect 78323 78513 78340 78565
rect 78392 78513 78409 78565
rect 78323 78501 78409 78513
rect 78323 78449 78340 78501
rect 78392 78449 78409 78501
rect 78323 78437 78409 78449
rect 78323 78385 78340 78437
rect 78392 78385 78409 78437
rect 78323 78373 78409 78385
rect 78323 78321 78340 78373
rect 78392 78321 78409 78373
rect 78323 78309 78409 78321
rect 78323 78257 78340 78309
rect 78392 78257 78409 78309
rect 78323 78245 78409 78257
rect 78323 78193 78340 78245
rect 78392 78193 78409 78245
rect 78323 78188 78409 78193
rect 79411 78757 79497 78762
rect 79411 78705 79428 78757
rect 79480 78705 79497 78757
rect 79411 78693 79497 78705
rect 79411 78641 79428 78693
rect 79480 78641 79497 78693
rect 79411 78629 79497 78641
rect 79411 78577 79428 78629
rect 79480 78577 79497 78629
rect 79411 78565 79497 78577
rect 79411 78513 79428 78565
rect 79480 78513 79497 78565
rect 79411 78501 79497 78513
rect 79411 78449 79428 78501
rect 79480 78449 79497 78501
rect 79411 78437 79497 78449
rect 79411 78385 79428 78437
rect 79480 78385 79497 78437
rect 79411 78373 79497 78385
rect 79411 78321 79428 78373
rect 79480 78321 79497 78373
rect 79411 78309 79497 78321
rect 79411 78257 79428 78309
rect 79480 78257 79497 78309
rect 79411 78245 79497 78257
rect 79411 78193 79428 78245
rect 79480 78193 79497 78245
rect 79411 78188 79497 78193
rect 80499 78757 80585 78762
rect 80499 78705 80516 78757
rect 80568 78705 80585 78757
rect 80499 78693 80585 78705
rect 80499 78641 80516 78693
rect 80568 78641 80585 78693
rect 80499 78629 80585 78641
rect 80499 78577 80516 78629
rect 80568 78577 80585 78629
rect 80499 78565 80585 78577
rect 80499 78513 80516 78565
rect 80568 78513 80585 78565
rect 80499 78501 80585 78513
rect 80499 78449 80516 78501
rect 80568 78449 80585 78501
rect 80499 78437 80585 78449
rect 80499 78385 80516 78437
rect 80568 78385 80585 78437
rect 80499 78373 80585 78385
rect 80499 78321 80516 78373
rect 80568 78321 80585 78373
rect 80499 78309 80585 78321
rect 80499 78257 80516 78309
rect 80568 78257 80585 78309
rect 80499 78245 80585 78257
rect 80499 78193 80516 78245
rect 80568 78193 80585 78245
rect 80499 78188 80585 78193
rect 81587 78757 81673 78762
rect 81587 78705 81604 78757
rect 81656 78705 81673 78757
rect 81587 78693 81673 78705
rect 81587 78641 81604 78693
rect 81656 78641 81673 78693
rect 81587 78629 81673 78641
rect 81587 78577 81604 78629
rect 81656 78577 81673 78629
rect 81587 78565 81673 78577
rect 81587 78513 81604 78565
rect 81656 78513 81673 78565
rect 81587 78501 81673 78513
rect 81587 78449 81604 78501
rect 81656 78449 81673 78501
rect 81587 78437 81673 78449
rect 81587 78385 81604 78437
rect 81656 78385 81673 78437
rect 81587 78373 81673 78385
rect 81587 78321 81604 78373
rect 81656 78321 81673 78373
rect 81587 78309 81673 78321
rect 81587 78257 81604 78309
rect 81656 78257 81673 78309
rect 81587 78245 81673 78257
rect 81587 78193 81604 78245
rect 81656 78193 81673 78245
rect 81587 78188 81673 78193
rect 82675 78757 82761 78762
rect 82675 78705 82692 78757
rect 82744 78705 82761 78757
rect 82675 78693 82761 78705
rect 82675 78641 82692 78693
rect 82744 78641 82761 78693
rect 82675 78629 82761 78641
rect 82675 78577 82692 78629
rect 82744 78577 82761 78629
rect 82675 78565 82761 78577
rect 82675 78513 82692 78565
rect 82744 78513 82761 78565
rect 82675 78501 82761 78513
rect 82675 78449 82692 78501
rect 82744 78449 82761 78501
rect 82675 78437 82761 78449
rect 82675 78385 82692 78437
rect 82744 78385 82761 78437
rect 82675 78373 82761 78385
rect 82675 78321 82692 78373
rect 82744 78321 82761 78373
rect 82675 78309 82761 78321
rect 82675 78257 82692 78309
rect 82744 78257 82761 78309
rect 82675 78245 82761 78257
rect 82675 78193 82692 78245
rect 82744 78193 82761 78245
rect 82675 78188 82761 78193
rect 83763 78757 83849 78762
rect 83763 78705 83780 78757
rect 83832 78705 83849 78757
rect 83763 78693 83849 78705
rect 83763 78641 83780 78693
rect 83832 78641 83849 78693
rect 83763 78629 83849 78641
rect 83763 78577 83780 78629
rect 83832 78577 83849 78629
rect 83763 78565 83849 78577
rect 83763 78513 83780 78565
rect 83832 78513 83849 78565
rect 83763 78501 83849 78513
rect 83763 78449 83780 78501
rect 83832 78449 83849 78501
rect 83763 78437 83849 78449
rect 83763 78385 83780 78437
rect 83832 78385 83849 78437
rect 83763 78373 83849 78385
rect 83763 78321 83780 78373
rect 83832 78321 83849 78373
rect 83763 78309 83849 78321
rect 83763 78257 83780 78309
rect 83832 78257 83849 78309
rect 83763 78245 83849 78257
rect 83763 78193 83780 78245
rect 83832 78193 83849 78245
rect 83763 78188 83849 78193
rect 84851 78757 84937 78762
rect 84851 78705 84868 78757
rect 84920 78705 84937 78757
rect 84851 78693 84937 78705
rect 84851 78641 84868 78693
rect 84920 78641 84937 78693
rect 84851 78629 84937 78641
rect 84851 78577 84868 78629
rect 84920 78577 84937 78629
rect 84851 78565 84937 78577
rect 84851 78513 84868 78565
rect 84920 78513 84937 78565
rect 84851 78501 84937 78513
rect 84851 78449 84868 78501
rect 84920 78449 84937 78501
rect 84851 78437 84937 78449
rect 84851 78385 84868 78437
rect 84920 78385 84937 78437
rect 84851 78373 84937 78385
rect 84851 78321 84868 78373
rect 84920 78321 84937 78373
rect 84851 78309 84937 78321
rect 84851 78257 84868 78309
rect 84920 78257 84937 78309
rect 84851 78245 84937 78257
rect 84851 78193 84868 78245
rect 84920 78193 84937 78245
rect 84851 78188 84937 78193
rect 85939 78757 86025 78762
rect 85939 78705 85956 78757
rect 86008 78705 86025 78757
rect 85939 78693 86025 78705
rect 85939 78641 85956 78693
rect 86008 78641 86025 78693
rect 85939 78629 86025 78641
rect 85939 78577 85956 78629
rect 86008 78577 86025 78629
rect 85939 78565 86025 78577
rect 85939 78513 85956 78565
rect 86008 78513 86025 78565
rect 85939 78501 86025 78513
rect 85939 78449 85956 78501
rect 86008 78449 86025 78501
rect 85939 78437 86025 78449
rect 85939 78385 85956 78437
rect 86008 78385 86025 78437
rect 85939 78373 86025 78385
rect 85939 78321 85956 78373
rect 86008 78321 86025 78373
rect 85939 78309 86025 78321
rect 85939 78257 85956 78309
rect 86008 78257 86025 78309
rect 85939 78245 86025 78257
rect 85939 78193 85956 78245
rect 86008 78193 86025 78245
rect 85939 78188 86025 78193
rect 87027 78757 87113 78762
rect 87027 78705 87044 78757
rect 87096 78705 87113 78757
rect 87027 78693 87113 78705
rect 87027 78641 87044 78693
rect 87096 78641 87113 78693
rect 87027 78629 87113 78641
rect 87027 78577 87044 78629
rect 87096 78577 87113 78629
rect 87027 78565 87113 78577
rect 87027 78513 87044 78565
rect 87096 78513 87113 78565
rect 87027 78501 87113 78513
rect 87027 78449 87044 78501
rect 87096 78449 87113 78501
rect 87027 78437 87113 78449
rect 87027 78385 87044 78437
rect 87096 78385 87113 78437
rect 87027 78373 87113 78385
rect 87027 78321 87044 78373
rect 87096 78321 87113 78373
rect 87027 78309 87113 78321
rect 87027 78257 87044 78309
rect 87096 78257 87113 78309
rect 87027 78245 87113 78257
rect 87027 78193 87044 78245
rect 87096 78193 87113 78245
rect 87027 78188 87113 78193
rect 88115 78757 88201 78762
rect 88115 78705 88132 78757
rect 88184 78705 88201 78757
rect 88115 78693 88201 78705
rect 88115 78641 88132 78693
rect 88184 78641 88201 78693
rect 88115 78629 88201 78641
rect 88115 78577 88132 78629
rect 88184 78577 88201 78629
rect 88115 78565 88201 78577
rect 88115 78513 88132 78565
rect 88184 78513 88201 78565
rect 88115 78501 88201 78513
rect 88115 78449 88132 78501
rect 88184 78449 88201 78501
rect 88115 78437 88201 78449
rect 88115 78385 88132 78437
rect 88184 78385 88201 78437
rect 88115 78373 88201 78385
rect 88115 78321 88132 78373
rect 88184 78321 88201 78373
rect 88115 78309 88201 78321
rect 88115 78257 88132 78309
rect 88184 78257 88201 78309
rect 88115 78245 88201 78257
rect 88115 78193 88132 78245
rect 88184 78193 88201 78245
rect 88115 78188 88201 78193
rect 74514 76760 74600 76765
rect 74514 76708 74531 76760
rect 74583 76708 74600 76760
rect 74514 76696 74600 76708
rect 74514 76644 74531 76696
rect 74583 76644 74600 76696
rect 74514 76632 74600 76644
rect 74514 76580 74531 76632
rect 74583 76580 74600 76632
rect 74514 76568 74600 76580
rect 74514 76516 74531 76568
rect 74583 76516 74600 76568
rect 74514 76504 74600 76516
rect 74514 76452 74531 76504
rect 74583 76452 74600 76504
rect 74514 76440 74600 76452
rect 74514 76388 74531 76440
rect 74583 76388 74600 76440
rect 74514 76376 74600 76388
rect 74514 76324 74531 76376
rect 74583 76324 74600 76376
rect 74514 76312 74600 76324
rect 74514 76260 74531 76312
rect 74583 76260 74600 76312
rect 74514 76248 74600 76260
rect 74514 76196 74531 76248
rect 74583 76196 74600 76248
rect 74514 76191 74600 76196
rect 75602 76760 75688 76765
rect 75602 76708 75619 76760
rect 75671 76708 75688 76760
rect 75602 76696 75688 76708
rect 75602 76644 75619 76696
rect 75671 76644 75688 76696
rect 75602 76632 75688 76644
rect 75602 76580 75619 76632
rect 75671 76580 75688 76632
rect 75602 76568 75688 76580
rect 75602 76516 75619 76568
rect 75671 76516 75688 76568
rect 75602 76504 75688 76516
rect 75602 76452 75619 76504
rect 75671 76452 75688 76504
rect 75602 76440 75688 76452
rect 75602 76388 75619 76440
rect 75671 76388 75688 76440
rect 75602 76376 75688 76388
rect 75602 76324 75619 76376
rect 75671 76324 75688 76376
rect 75602 76312 75688 76324
rect 75602 76260 75619 76312
rect 75671 76260 75688 76312
rect 75602 76248 75688 76260
rect 75602 76196 75619 76248
rect 75671 76196 75688 76248
rect 75602 76191 75688 76196
rect 76690 76760 76776 76765
rect 76690 76708 76707 76760
rect 76759 76708 76776 76760
rect 76690 76696 76776 76708
rect 76690 76644 76707 76696
rect 76759 76644 76776 76696
rect 76690 76632 76776 76644
rect 76690 76580 76707 76632
rect 76759 76580 76776 76632
rect 76690 76568 76776 76580
rect 76690 76516 76707 76568
rect 76759 76516 76776 76568
rect 76690 76504 76776 76516
rect 76690 76452 76707 76504
rect 76759 76452 76776 76504
rect 76690 76440 76776 76452
rect 76690 76388 76707 76440
rect 76759 76388 76776 76440
rect 76690 76376 76776 76388
rect 76690 76324 76707 76376
rect 76759 76324 76776 76376
rect 76690 76312 76776 76324
rect 76690 76260 76707 76312
rect 76759 76260 76776 76312
rect 76690 76248 76776 76260
rect 76690 76196 76707 76248
rect 76759 76196 76776 76248
rect 76690 76191 76776 76196
rect 77778 76760 77864 76765
rect 77778 76708 77795 76760
rect 77847 76708 77864 76760
rect 77778 76696 77864 76708
rect 77778 76644 77795 76696
rect 77847 76644 77864 76696
rect 77778 76632 77864 76644
rect 77778 76580 77795 76632
rect 77847 76580 77864 76632
rect 77778 76568 77864 76580
rect 77778 76516 77795 76568
rect 77847 76516 77864 76568
rect 77778 76504 77864 76516
rect 77778 76452 77795 76504
rect 77847 76452 77864 76504
rect 77778 76440 77864 76452
rect 77778 76388 77795 76440
rect 77847 76388 77864 76440
rect 77778 76376 77864 76388
rect 77778 76324 77795 76376
rect 77847 76324 77864 76376
rect 77778 76312 77864 76324
rect 77778 76260 77795 76312
rect 77847 76260 77864 76312
rect 77778 76248 77864 76260
rect 77778 76196 77795 76248
rect 77847 76196 77864 76248
rect 77778 76191 77864 76196
rect 78866 76760 78952 76765
rect 78866 76708 78883 76760
rect 78935 76708 78952 76760
rect 78866 76696 78952 76708
rect 78866 76644 78883 76696
rect 78935 76644 78952 76696
rect 78866 76632 78952 76644
rect 78866 76580 78883 76632
rect 78935 76580 78952 76632
rect 78866 76568 78952 76580
rect 78866 76516 78883 76568
rect 78935 76516 78952 76568
rect 78866 76504 78952 76516
rect 78866 76452 78883 76504
rect 78935 76452 78952 76504
rect 78866 76440 78952 76452
rect 78866 76388 78883 76440
rect 78935 76388 78952 76440
rect 78866 76376 78952 76388
rect 78866 76324 78883 76376
rect 78935 76324 78952 76376
rect 78866 76312 78952 76324
rect 78866 76260 78883 76312
rect 78935 76260 78952 76312
rect 78866 76248 78952 76260
rect 78866 76196 78883 76248
rect 78935 76196 78952 76248
rect 78866 76191 78952 76196
rect 79954 76760 80040 76765
rect 79954 76708 79971 76760
rect 80023 76708 80040 76760
rect 79954 76696 80040 76708
rect 79954 76644 79971 76696
rect 80023 76644 80040 76696
rect 79954 76632 80040 76644
rect 79954 76580 79971 76632
rect 80023 76580 80040 76632
rect 79954 76568 80040 76580
rect 79954 76516 79971 76568
rect 80023 76516 80040 76568
rect 79954 76504 80040 76516
rect 79954 76452 79971 76504
rect 80023 76452 80040 76504
rect 79954 76440 80040 76452
rect 79954 76388 79971 76440
rect 80023 76388 80040 76440
rect 79954 76376 80040 76388
rect 79954 76324 79971 76376
rect 80023 76324 80040 76376
rect 79954 76312 80040 76324
rect 79954 76260 79971 76312
rect 80023 76260 80040 76312
rect 79954 76248 80040 76260
rect 79954 76196 79971 76248
rect 80023 76196 80040 76248
rect 79954 76191 80040 76196
rect 81042 76760 81128 76765
rect 81042 76708 81059 76760
rect 81111 76708 81128 76760
rect 81042 76696 81128 76708
rect 81042 76644 81059 76696
rect 81111 76644 81128 76696
rect 81042 76632 81128 76644
rect 81042 76580 81059 76632
rect 81111 76580 81128 76632
rect 81042 76568 81128 76580
rect 81042 76516 81059 76568
rect 81111 76516 81128 76568
rect 81042 76504 81128 76516
rect 81042 76452 81059 76504
rect 81111 76452 81128 76504
rect 81042 76440 81128 76452
rect 81042 76388 81059 76440
rect 81111 76388 81128 76440
rect 81042 76376 81128 76388
rect 81042 76324 81059 76376
rect 81111 76324 81128 76376
rect 81042 76312 81128 76324
rect 81042 76260 81059 76312
rect 81111 76260 81128 76312
rect 81042 76248 81128 76260
rect 81042 76196 81059 76248
rect 81111 76196 81128 76248
rect 81042 76191 81128 76196
rect 82130 76760 82216 76765
rect 82130 76708 82147 76760
rect 82199 76708 82216 76760
rect 82130 76696 82216 76708
rect 82130 76644 82147 76696
rect 82199 76644 82216 76696
rect 82130 76632 82216 76644
rect 82130 76580 82147 76632
rect 82199 76580 82216 76632
rect 82130 76568 82216 76580
rect 82130 76516 82147 76568
rect 82199 76516 82216 76568
rect 82130 76504 82216 76516
rect 82130 76452 82147 76504
rect 82199 76452 82216 76504
rect 82130 76440 82216 76452
rect 82130 76388 82147 76440
rect 82199 76388 82216 76440
rect 82130 76376 82216 76388
rect 82130 76324 82147 76376
rect 82199 76324 82216 76376
rect 82130 76312 82216 76324
rect 82130 76260 82147 76312
rect 82199 76260 82216 76312
rect 82130 76248 82216 76260
rect 82130 76196 82147 76248
rect 82199 76196 82216 76248
rect 82130 76191 82216 76196
rect 83218 76760 83304 76765
rect 83218 76708 83235 76760
rect 83287 76708 83304 76760
rect 83218 76696 83304 76708
rect 83218 76644 83235 76696
rect 83287 76644 83304 76696
rect 83218 76632 83304 76644
rect 83218 76580 83235 76632
rect 83287 76580 83304 76632
rect 83218 76568 83304 76580
rect 83218 76516 83235 76568
rect 83287 76516 83304 76568
rect 83218 76504 83304 76516
rect 83218 76452 83235 76504
rect 83287 76452 83304 76504
rect 83218 76440 83304 76452
rect 83218 76388 83235 76440
rect 83287 76388 83304 76440
rect 83218 76376 83304 76388
rect 83218 76324 83235 76376
rect 83287 76324 83304 76376
rect 83218 76312 83304 76324
rect 83218 76260 83235 76312
rect 83287 76260 83304 76312
rect 83218 76248 83304 76260
rect 83218 76196 83235 76248
rect 83287 76196 83304 76248
rect 83218 76191 83304 76196
rect 84306 76760 84392 76765
rect 84306 76708 84323 76760
rect 84375 76708 84392 76760
rect 84306 76696 84392 76708
rect 84306 76644 84323 76696
rect 84375 76644 84392 76696
rect 84306 76632 84392 76644
rect 84306 76580 84323 76632
rect 84375 76580 84392 76632
rect 84306 76568 84392 76580
rect 84306 76516 84323 76568
rect 84375 76516 84392 76568
rect 84306 76504 84392 76516
rect 84306 76452 84323 76504
rect 84375 76452 84392 76504
rect 84306 76440 84392 76452
rect 84306 76388 84323 76440
rect 84375 76388 84392 76440
rect 84306 76376 84392 76388
rect 84306 76324 84323 76376
rect 84375 76324 84392 76376
rect 84306 76312 84392 76324
rect 84306 76260 84323 76312
rect 84375 76260 84392 76312
rect 84306 76248 84392 76260
rect 84306 76196 84323 76248
rect 84375 76196 84392 76248
rect 84306 76191 84392 76196
rect 85394 76760 85480 76765
rect 85394 76708 85411 76760
rect 85463 76708 85480 76760
rect 85394 76696 85480 76708
rect 85394 76644 85411 76696
rect 85463 76644 85480 76696
rect 85394 76632 85480 76644
rect 85394 76580 85411 76632
rect 85463 76580 85480 76632
rect 85394 76568 85480 76580
rect 85394 76516 85411 76568
rect 85463 76516 85480 76568
rect 85394 76504 85480 76516
rect 85394 76452 85411 76504
rect 85463 76452 85480 76504
rect 85394 76440 85480 76452
rect 85394 76388 85411 76440
rect 85463 76388 85480 76440
rect 85394 76376 85480 76388
rect 85394 76324 85411 76376
rect 85463 76324 85480 76376
rect 85394 76312 85480 76324
rect 85394 76260 85411 76312
rect 85463 76260 85480 76312
rect 85394 76248 85480 76260
rect 85394 76196 85411 76248
rect 85463 76196 85480 76248
rect 85394 76191 85480 76196
rect 86482 76760 86568 76765
rect 86482 76708 86499 76760
rect 86551 76708 86568 76760
rect 86482 76696 86568 76708
rect 86482 76644 86499 76696
rect 86551 76644 86568 76696
rect 86482 76632 86568 76644
rect 86482 76580 86499 76632
rect 86551 76580 86568 76632
rect 86482 76568 86568 76580
rect 86482 76516 86499 76568
rect 86551 76516 86568 76568
rect 86482 76504 86568 76516
rect 86482 76452 86499 76504
rect 86551 76452 86568 76504
rect 86482 76440 86568 76452
rect 86482 76388 86499 76440
rect 86551 76388 86568 76440
rect 86482 76376 86568 76388
rect 86482 76324 86499 76376
rect 86551 76324 86568 76376
rect 86482 76312 86568 76324
rect 86482 76260 86499 76312
rect 86551 76260 86568 76312
rect 86482 76248 86568 76260
rect 86482 76196 86499 76248
rect 86551 76196 86568 76248
rect 86482 76191 86568 76196
rect 87570 76760 87656 76765
rect 87570 76708 87587 76760
rect 87639 76708 87656 76760
rect 87570 76696 87656 76708
rect 87570 76644 87587 76696
rect 87639 76644 87656 76696
rect 87570 76632 87656 76644
rect 87570 76580 87587 76632
rect 87639 76580 87656 76632
rect 87570 76568 87656 76580
rect 87570 76516 87587 76568
rect 87639 76516 87656 76568
rect 87570 76504 87656 76516
rect 87570 76452 87587 76504
rect 87639 76452 87656 76504
rect 87570 76440 87656 76452
rect 87570 76388 87587 76440
rect 87639 76388 87656 76440
rect 87570 76376 87656 76388
rect 87570 76324 87587 76376
rect 87639 76324 87656 76376
rect 87570 76312 87656 76324
rect 87570 76260 87587 76312
rect 87639 76260 87656 76312
rect 87570 76248 87656 76260
rect 87570 76196 87587 76248
rect 87639 76196 87656 76248
rect 87570 76191 87656 76196
rect 88658 76760 88744 76765
rect 88658 76708 88675 76760
rect 88727 76708 88744 76760
rect 88658 76696 88744 76708
rect 88658 76644 88675 76696
rect 88727 76644 88744 76696
rect 88658 76632 88744 76644
rect 88658 76580 88675 76632
rect 88727 76580 88744 76632
rect 88658 76568 88744 76580
rect 88658 76516 88675 76568
rect 88727 76516 88744 76568
rect 88658 76504 88744 76516
rect 88658 76452 88675 76504
rect 88727 76452 88744 76504
rect 88658 76440 88744 76452
rect 88658 76388 88675 76440
rect 88727 76388 88744 76440
rect 88658 76376 88744 76388
rect 88658 76324 88675 76376
rect 88727 76324 88744 76376
rect 88658 76312 88744 76324
rect 88658 76260 88675 76312
rect 88727 76260 88744 76312
rect 88658 76248 88744 76260
rect 88658 76196 88675 76248
rect 88727 76196 88744 76248
rect 88658 76191 88744 76196
rect 75059 74757 75145 74762
rect 75059 74705 75076 74757
rect 75128 74705 75145 74757
rect 75059 74693 75145 74705
rect 75059 74641 75076 74693
rect 75128 74641 75145 74693
rect 75059 74629 75145 74641
rect 75059 74577 75076 74629
rect 75128 74577 75145 74629
rect 75059 74565 75145 74577
rect 75059 74513 75076 74565
rect 75128 74513 75145 74565
rect 75059 74501 75145 74513
rect 75059 74449 75076 74501
rect 75128 74449 75145 74501
rect 75059 74437 75145 74449
rect 75059 74385 75076 74437
rect 75128 74385 75145 74437
rect 75059 74373 75145 74385
rect 75059 74321 75076 74373
rect 75128 74321 75145 74373
rect 75059 74309 75145 74321
rect 75059 74257 75076 74309
rect 75128 74257 75145 74309
rect 75059 74245 75145 74257
rect 75059 74193 75076 74245
rect 75128 74193 75145 74245
rect 75059 74188 75145 74193
rect 77235 74757 77321 74762
rect 77235 74705 77252 74757
rect 77304 74705 77321 74757
rect 77235 74693 77321 74705
rect 77235 74641 77252 74693
rect 77304 74641 77321 74693
rect 77235 74629 77321 74641
rect 77235 74577 77252 74629
rect 77304 74577 77321 74629
rect 77235 74565 77321 74577
rect 77235 74513 77252 74565
rect 77304 74513 77321 74565
rect 77235 74501 77321 74513
rect 77235 74449 77252 74501
rect 77304 74449 77321 74501
rect 77235 74437 77321 74449
rect 77235 74385 77252 74437
rect 77304 74385 77321 74437
rect 77235 74373 77321 74385
rect 77235 74321 77252 74373
rect 77304 74321 77321 74373
rect 77235 74309 77321 74321
rect 77235 74257 77252 74309
rect 77304 74257 77321 74309
rect 77235 74245 77321 74257
rect 77235 74193 77252 74245
rect 77304 74193 77321 74245
rect 77235 74188 77321 74193
rect 78323 74757 78409 74762
rect 78323 74705 78340 74757
rect 78392 74705 78409 74757
rect 78323 74693 78409 74705
rect 78323 74641 78340 74693
rect 78392 74641 78409 74693
rect 78323 74629 78409 74641
rect 78323 74577 78340 74629
rect 78392 74577 78409 74629
rect 78323 74565 78409 74577
rect 78323 74513 78340 74565
rect 78392 74513 78409 74565
rect 78323 74501 78409 74513
rect 78323 74449 78340 74501
rect 78392 74449 78409 74501
rect 78323 74437 78409 74449
rect 78323 74385 78340 74437
rect 78392 74385 78409 74437
rect 78323 74373 78409 74385
rect 78323 74321 78340 74373
rect 78392 74321 78409 74373
rect 78323 74309 78409 74321
rect 78323 74257 78340 74309
rect 78392 74257 78409 74309
rect 78323 74245 78409 74257
rect 78323 74193 78340 74245
rect 78392 74193 78409 74245
rect 78323 74188 78409 74193
rect 80499 74757 80585 74762
rect 80499 74705 80516 74757
rect 80568 74705 80585 74757
rect 80499 74693 80585 74705
rect 80499 74641 80516 74693
rect 80568 74641 80585 74693
rect 80499 74629 80585 74641
rect 80499 74577 80516 74629
rect 80568 74577 80585 74629
rect 80499 74565 80585 74577
rect 80499 74513 80516 74565
rect 80568 74513 80585 74565
rect 80499 74501 80585 74513
rect 80499 74449 80516 74501
rect 80568 74449 80585 74501
rect 80499 74437 80585 74449
rect 80499 74385 80516 74437
rect 80568 74385 80585 74437
rect 80499 74373 80585 74385
rect 80499 74321 80516 74373
rect 80568 74321 80585 74373
rect 80499 74309 80585 74321
rect 80499 74257 80516 74309
rect 80568 74257 80585 74309
rect 80499 74245 80585 74257
rect 80499 74193 80516 74245
rect 80568 74193 80585 74245
rect 80499 74188 80585 74193
rect 81587 74757 81673 74762
rect 81587 74705 81604 74757
rect 81656 74705 81673 74757
rect 81587 74693 81673 74705
rect 81587 74641 81604 74693
rect 81656 74641 81673 74693
rect 81587 74629 81673 74641
rect 81587 74577 81604 74629
rect 81656 74577 81673 74629
rect 81587 74565 81673 74577
rect 81587 74513 81604 74565
rect 81656 74513 81673 74565
rect 81587 74501 81673 74513
rect 81587 74449 81604 74501
rect 81656 74449 81673 74501
rect 81587 74437 81673 74449
rect 81587 74385 81604 74437
rect 81656 74385 81673 74437
rect 81587 74373 81673 74385
rect 81587 74321 81604 74373
rect 81656 74321 81673 74373
rect 81587 74309 81673 74321
rect 81587 74257 81604 74309
rect 81656 74257 81673 74309
rect 81587 74245 81673 74257
rect 81587 74193 81604 74245
rect 81656 74193 81673 74245
rect 81587 74188 81673 74193
rect 82675 74757 82761 74762
rect 82675 74705 82692 74757
rect 82744 74705 82761 74757
rect 82675 74693 82761 74705
rect 82675 74641 82692 74693
rect 82744 74641 82761 74693
rect 82675 74629 82761 74641
rect 82675 74577 82692 74629
rect 82744 74577 82761 74629
rect 82675 74565 82761 74577
rect 82675 74513 82692 74565
rect 82744 74513 82761 74565
rect 82675 74501 82761 74513
rect 82675 74449 82692 74501
rect 82744 74449 82761 74501
rect 82675 74437 82761 74449
rect 82675 74385 82692 74437
rect 82744 74385 82761 74437
rect 82675 74373 82761 74385
rect 82675 74321 82692 74373
rect 82744 74321 82761 74373
rect 82675 74309 82761 74321
rect 82675 74257 82692 74309
rect 82744 74257 82761 74309
rect 82675 74245 82761 74257
rect 82675 74193 82692 74245
rect 82744 74193 82761 74245
rect 82675 74188 82761 74193
rect 84851 74757 84937 74762
rect 84851 74705 84868 74757
rect 84920 74705 84937 74757
rect 84851 74693 84937 74705
rect 84851 74641 84868 74693
rect 84920 74641 84937 74693
rect 84851 74629 84937 74641
rect 84851 74577 84868 74629
rect 84920 74577 84937 74629
rect 84851 74565 84937 74577
rect 84851 74513 84868 74565
rect 84920 74513 84937 74565
rect 84851 74501 84937 74513
rect 84851 74449 84868 74501
rect 84920 74449 84937 74501
rect 84851 74437 84937 74449
rect 84851 74385 84868 74437
rect 84920 74385 84937 74437
rect 84851 74373 84937 74385
rect 84851 74321 84868 74373
rect 84920 74321 84937 74373
rect 84851 74309 84937 74321
rect 84851 74257 84868 74309
rect 84920 74257 84937 74309
rect 84851 74245 84937 74257
rect 84851 74193 84868 74245
rect 84920 74193 84937 74245
rect 84851 74188 84937 74193
rect 85939 74757 86025 74762
rect 85939 74705 85956 74757
rect 86008 74705 86025 74757
rect 85939 74693 86025 74705
rect 85939 74641 85956 74693
rect 86008 74641 86025 74693
rect 85939 74629 86025 74641
rect 85939 74577 85956 74629
rect 86008 74577 86025 74629
rect 85939 74565 86025 74577
rect 85939 74513 85956 74565
rect 86008 74513 86025 74565
rect 85939 74501 86025 74513
rect 85939 74449 85956 74501
rect 86008 74449 86025 74501
rect 85939 74437 86025 74449
rect 85939 74385 85956 74437
rect 86008 74385 86025 74437
rect 85939 74373 86025 74385
rect 85939 74321 85956 74373
rect 86008 74321 86025 74373
rect 85939 74309 86025 74321
rect 85939 74257 85956 74309
rect 86008 74257 86025 74309
rect 85939 74245 86025 74257
rect 85939 74193 85956 74245
rect 86008 74193 86025 74245
rect 85939 74188 86025 74193
rect 88115 74757 88201 74762
rect 88115 74705 88132 74757
rect 88184 74705 88201 74757
rect 88115 74693 88201 74705
rect 88115 74641 88132 74693
rect 88184 74641 88201 74693
rect 88115 74629 88201 74641
rect 88115 74577 88132 74629
rect 88184 74577 88201 74629
rect 88115 74565 88201 74577
rect 88115 74513 88132 74565
rect 88184 74513 88201 74565
rect 88115 74501 88201 74513
rect 88115 74449 88132 74501
rect 88184 74449 88201 74501
rect 88115 74437 88201 74449
rect 88115 74385 88132 74437
rect 88184 74385 88201 74437
rect 88115 74373 88201 74385
rect 88115 74321 88132 74373
rect 88184 74321 88201 74373
rect 88115 74309 88201 74321
rect 88115 74257 88132 74309
rect 88184 74257 88201 74309
rect 88115 74245 88201 74257
rect 88115 74193 88132 74245
rect 88184 74193 88201 74245
rect 88115 74188 88201 74193
rect 74514 72760 74600 72765
rect 74514 72708 74531 72760
rect 74583 72708 74600 72760
rect 74514 72696 74600 72708
rect 74514 72644 74531 72696
rect 74583 72644 74600 72696
rect 74514 72632 74600 72644
rect 74514 72580 74531 72632
rect 74583 72580 74600 72632
rect 74514 72568 74600 72580
rect 74514 72516 74531 72568
rect 74583 72516 74600 72568
rect 74514 72504 74600 72516
rect 74514 72452 74531 72504
rect 74583 72452 74600 72504
rect 74514 72440 74600 72452
rect 74514 72388 74531 72440
rect 74583 72388 74600 72440
rect 74514 72376 74600 72388
rect 74514 72324 74531 72376
rect 74583 72324 74600 72376
rect 74514 72312 74600 72324
rect 74514 72260 74531 72312
rect 74583 72260 74600 72312
rect 74514 72248 74600 72260
rect 74514 72196 74531 72248
rect 74583 72196 74600 72248
rect 74514 72191 74600 72196
rect 75602 72760 75688 72765
rect 75602 72708 75619 72760
rect 75671 72708 75688 72760
rect 75602 72696 75688 72708
rect 75602 72644 75619 72696
rect 75671 72644 75688 72696
rect 75602 72632 75688 72644
rect 75602 72580 75619 72632
rect 75671 72580 75688 72632
rect 75602 72568 75688 72580
rect 75602 72516 75619 72568
rect 75671 72516 75688 72568
rect 75602 72504 75688 72516
rect 75602 72452 75619 72504
rect 75671 72452 75688 72504
rect 75602 72440 75688 72452
rect 75602 72388 75619 72440
rect 75671 72388 75688 72440
rect 75602 72376 75688 72388
rect 75602 72324 75619 72376
rect 75671 72324 75688 72376
rect 75602 72312 75688 72324
rect 75602 72260 75619 72312
rect 75671 72260 75688 72312
rect 75602 72248 75688 72260
rect 75602 72196 75619 72248
rect 75671 72196 75688 72248
rect 75602 72191 75688 72196
rect 76690 72760 76776 72765
rect 76690 72708 76707 72760
rect 76759 72708 76776 72760
rect 76690 72696 76776 72708
rect 76690 72644 76707 72696
rect 76759 72644 76776 72696
rect 76690 72632 76776 72644
rect 76690 72580 76707 72632
rect 76759 72580 76776 72632
rect 76690 72568 76776 72580
rect 76690 72516 76707 72568
rect 76759 72516 76776 72568
rect 76690 72504 76776 72516
rect 76690 72452 76707 72504
rect 76759 72452 76776 72504
rect 76690 72440 76776 72452
rect 76690 72388 76707 72440
rect 76759 72388 76776 72440
rect 76690 72376 76776 72388
rect 76690 72324 76707 72376
rect 76759 72324 76776 72376
rect 76690 72312 76776 72324
rect 76690 72260 76707 72312
rect 76759 72260 76776 72312
rect 76690 72248 76776 72260
rect 76690 72196 76707 72248
rect 76759 72196 76776 72248
rect 76690 72191 76776 72196
rect 77778 72760 77864 72765
rect 77778 72708 77795 72760
rect 77847 72708 77864 72760
rect 77778 72696 77864 72708
rect 77778 72644 77795 72696
rect 77847 72644 77864 72696
rect 77778 72632 77864 72644
rect 77778 72580 77795 72632
rect 77847 72580 77864 72632
rect 77778 72568 77864 72580
rect 77778 72516 77795 72568
rect 77847 72516 77864 72568
rect 77778 72504 77864 72516
rect 77778 72452 77795 72504
rect 77847 72452 77864 72504
rect 77778 72440 77864 72452
rect 77778 72388 77795 72440
rect 77847 72388 77864 72440
rect 77778 72376 77864 72388
rect 77778 72324 77795 72376
rect 77847 72324 77864 72376
rect 77778 72312 77864 72324
rect 77778 72260 77795 72312
rect 77847 72260 77864 72312
rect 77778 72248 77864 72260
rect 77778 72196 77795 72248
rect 77847 72196 77864 72248
rect 77778 72191 77864 72196
rect 78866 72760 78952 72765
rect 78866 72708 78883 72760
rect 78935 72708 78952 72760
rect 78866 72696 78952 72708
rect 78866 72644 78883 72696
rect 78935 72644 78952 72696
rect 78866 72632 78952 72644
rect 78866 72580 78883 72632
rect 78935 72580 78952 72632
rect 78866 72568 78952 72580
rect 78866 72516 78883 72568
rect 78935 72516 78952 72568
rect 78866 72504 78952 72516
rect 78866 72452 78883 72504
rect 78935 72452 78952 72504
rect 78866 72440 78952 72452
rect 78866 72388 78883 72440
rect 78935 72388 78952 72440
rect 78866 72376 78952 72388
rect 78866 72324 78883 72376
rect 78935 72324 78952 72376
rect 78866 72312 78952 72324
rect 78866 72260 78883 72312
rect 78935 72260 78952 72312
rect 78866 72248 78952 72260
rect 78866 72196 78883 72248
rect 78935 72196 78952 72248
rect 78866 72191 78952 72196
rect 79954 72760 80040 72765
rect 79954 72708 79971 72760
rect 80023 72708 80040 72760
rect 79954 72696 80040 72708
rect 79954 72644 79971 72696
rect 80023 72644 80040 72696
rect 79954 72632 80040 72644
rect 79954 72580 79971 72632
rect 80023 72580 80040 72632
rect 79954 72568 80040 72580
rect 79954 72516 79971 72568
rect 80023 72516 80040 72568
rect 79954 72504 80040 72516
rect 79954 72452 79971 72504
rect 80023 72452 80040 72504
rect 79954 72440 80040 72452
rect 79954 72388 79971 72440
rect 80023 72388 80040 72440
rect 79954 72376 80040 72388
rect 79954 72324 79971 72376
rect 80023 72324 80040 72376
rect 79954 72312 80040 72324
rect 79954 72260 79971 72312
rect 80023 72260 80040 72312
rect 79954 72248 80040 72260
rect 79954 72196 79971 72248
rect 80023 72196 80040 72248
rect 79954 72191 80040 72196
rect 81042 72760 81128 72765
rect 81042 72708 81059 72760
rect 81111 72708 81128 72760
rect 81042 72696 81128 72708
rect 81042 72644 81059 72696
rect 81111 72644 81128 72696
rect 81042 72632 81128 72644
rect 81042 72580 81059 72632
rect 81111 72580 81128 72632
rect 81042 72568 81128 72580
rect 81042 72516 81059 72568
rect 81111 72516 81128 72568
rect 81042 72504 81128 72516
rect 81042 72452 81059 72504
rect 81111 72452 81128 72504
rect 81042 72440 81128 72452
rect 81042 72388 81059 72440
rect 81111 72388 81128 72440
rect 81042 72376 81128 72388
rect 81042 72324 81059 72376
rect 81111 72324 81128 72376
rect 81042 72312 81128 72324
rect 81042 72260 81059 72312
rect 81111 72260 81128 72312
rect 81042 72248 81128 72260
rect 81042 72196 81059 72248
rect 81111 72196 81128 72248
rect 81042 72191 81128 72196
rect 86482 72760 86568 72765
rect 86482 72708 86499 72760
rect 86551 72708 86568 72760
rect 86482 72696 86568 72708
rect 86482 72644 86499 72696
rect 86551 72644 86568 72696
rect 86482 72632 86568 72644
rect 86482 72580 86499 72632
rect 86551 72580 86568 72632
rect 86482 72568 86568 72580
rect 86482 72516 86499 72568
rect 86551 72516 86568 72568
rect 86482 72504 86568 72516
rect 86482 72452 86499 72504
rect 86551 72452 86568 72504
rect 86482 72440 86568 72452
rect 86482 72388 86499 72440
rect 86551 72388 86568 72440
rect 86482 72376 86568 72388
rect 86482 72324 86499 72376
rect 86551 72324 86568 72376
rect 86482 72312 86568 72324
rect 86482 72260 86499 72312
rect 86551 72260 86568 72312
rect 86482 72248 86568 72260
rect 86482 72196 86499 72248
rect 86551 72196 86568 72248
rect 86482 72191 86568 72196
rect 87570 72760 87656 72765
rect 87570 72708 87587 72760
rect 87639 72708 87656 72760
rect 87570 72696 87656 72708
rect 87570 72644 87587 72696
rect 87639 72644 87656 72696
rect 87570 72632 87656 72644
rect 87570 72580 87587 72632
rect 87639 72580 87656 72632
rect 87570 72568 87656 72580
rect 87570 72516 87587 72568
rect 87639 72516 87656 72568
rect 87570 72504 87656 72516
rect 87570 72452 87587 72504
rect 87639 72452 87656 72504
rect 87570 72440 87656 72452
rect 87570 72388 87587 72440
rect 87639 72388 87656 72440
rect 87570 72376 87656 72388
rect 87570 72324 87587 72376
rect 87639 72324 87656 72376
rect 87570 72312 87656 72324
rect 87570 72260 87587 72312
rect 87639 72260 87656 72312
rect 87570 72248 87656 72260
rect 87570 72196 87587 72248
rect 87639 72196 87656 72248
rect 87570 72191 87656 72196
rect 88658 72760 88744 72765
rect 88658 72708 88675 72760
rect 88727 72708 88744 72760
rect 88658 72696 88744 72708
rect 88658 72644 88675 72696
rect 88727 72644 88744 72696
rect 88658 72632 88744 72644
rect 88658 72580 88675 72632
rect 88727 72580 88744 72632
rect 88658 72568 88744 72580
rect 88658 72516 88675 72568
rect 88727 72516 88744 72568
rect 88658 72504 88744 72516
rect 88658 72452 88675 72504
rect 88727 72452 88744 72504
rect 88658 72440 88744 72452
rect 88658 72388 88675 72440
rect 88727 72388 88744 72440
rect 88658 72376 88744 72388
rect 88658 72324 88675 72376
rect 88727 72324 88744 72376
rect 88658 72312 88744 72324
rect 88658 72260 88675 72312
rect 88727 72260 88744 72312
rect 88658 72248 88744 72260
rect 88658 72196 88675 72248
rect 88727 72196 88744 72248
rect 88658 72191 88744 72196
rect 75059 70757 75145 70762
rect 75059 70705 75076 70757
rect 75128 70705 75145 70757
rect 75059 70693 75145 70705
rect 75059 70641 75076 70693
rect 75128 70641 75145 70693
rect 75059 70629 75145 70641
rect 75059 70577 75076 70629
rect 75128 70577 75145 70629
rect 75059 70565 75145 70577
rect 75059 70513 75076 70565
rect 75128 70513 75145 70565
rect 75059 70501 75145 70513
rect 75059 70449 75076 70501
rect 75128 70449 75145 70501
rect 75059 70437 75145 70449
rect 75059 70385 75076 70437
rect 75128 70385 75145 70437
rect 75059 70373 75145 70385
rect 75059 70321 75076 70373
rect 75128 70321 75145 70373
rect 75059 70309 75145 70321
rect 75059 70257 75076 70309
rect 75128 70257 75145 70309
rect 75059 70245 75145 70257
rect 75059 70193 75076 70245
rect 75128 70193 75145 70245
rect 75059 70188 75145 70193
rect 76147 70757 76233 70762
rect 76147 70705 76164 70757
rect 76216 70705 76233 70757
rect 76147 70693 76233 70705
rect 76147 70641 76164 70693
rect 76216 70641 76233 70693
rect 76147 70629 76233 70641
rect 76147 70577 76164 70629
rect 76216 70577 76233 70629
rect 76147 70565 76233 70577
rect 76147 70513 76164 70565
rect 76216 70513 76233 70565
rect 76147 70501 76233 70513
rect 76147 70449 76164 70501
rect 76216 70449 76233 70501
rect 76147 70437 76233 70449
rect 76147 70385 76164 70437
rect 76216 70385 76233 70437
rect 76147 70373 76233 70385
rect 76147 70321 76164 70373
rect 76216 70321 76233 70373
rect 76147 70309 76233 70321
rect 76147 70257 76164 70309
rect 76216 70257 76233 70309
rect 76147 70245 76233 70257
rect 76147 70193 76164 70245
rect 76216 70193 76233 70245
rect 76147 70188 76233 70193
rect 77235 70757 77321 70762
rect 77235 70705 77252 70757
rect 77304 70705 77321 70757
rect 77235 70693 77321 70705
rect 77235 70641 77252 70693
rect 77304 70641 77321 70693
rect 77235 70629 77321 70641
rect 77235 70577 77252 70629
rect 77304 70577 77321 70629
rect 77235 70565 77321 70577
rect 77235 70513 77252 70565
rect 77304 70513 77321 70565
rect 77235 70501 77321 70513
rect 77235 70449 77252 70501
rect 77304 70449 77321 70501
rect 77235 70437 77321 70449
rect 77235 70385 77252 70437
rect 77304 70385 77321 70437
rect 77235 70373 77321 70385
rect 77235 70321 77252 70373
rect 77304 70321 77321 70373
rect 77235 70309 77321 70321
rect 77235 70257 77252 70309
rect 77304 70257 77321 70309
rect 77235 70245 77321 70257
rect 77235 70193 77252 70245
rect 77304 70193 77321 70245
rect 77235 70188 77321 70193
rect 78323 70757 78409 70762
rect 78323 70705 78340 70757
rect 78392 70705 78409 70757
rect 78323 70693 78409 70705
rect 78323 70641 78340 70693
rect 78392 70641 78409 70693
rect 78323 70629 78409 70641
rect 78323 70577 78340 70629
rect 78392 70577 78409 70629
rect 78323 70565 78409 70577
rect 78323 70513 78340 70565
rect 78392 70513 78409 70565
rect 78323 70501 78409 70513
rect 78323 70449 78340 70501
rect 78392 70449 78409 70501
rect 78323 70437 78409 70449
rect 78323 70385 78340 70437
rect 78392 70385 78409 70437
rect 78323 70373 78409 70385
rect 78323 70321 78340 70373
rect 78392 70321 78409 70373
rect 78323 70309 78409 70321
rect 78323 70257 78340 70309
rect 78392 70257 78409 70309
rect 78323 70245 78409 70257
rect 78323 70193 78340 70245
rect 78392 70193 78409 70245
rect 78323 70188 78409 70193
rect 79411 70757 79497 70762
rect 79411 70705 79428 70757
rect 79480 70705 79497 70757
rect 79411 70693 79497 70705
rect 79411 70641 79428 70693
rect 79480 70641 79497 70693
rect 79411 70629 79497 70641
rect 79411 70577 79428 70629
rect 79480 70577 79497 70629
rect 79411 70565 79497 70577
rect 79411 70513 79428 70565
rect 79480 70513 79497 70565
rect 79411 70501 79497 70513
rect 79411 70449 79428 70501
rect 79480 70449 79497 70501
rect 79411 70437 79497 70449
rect 79411 70385 79428 70437
rect 79480 70385 79497 70437
rect 79411 70373 79497 70385
rect 79411 70321 79428 70373
rect 79480 70321 79497 70373
rect 79411 70309 79497 70321
rect 79411 70257 79428 70309
rect 79480 70257 79497 70309
rect 79411 70245 79497 70257
rect 79411 70193 79428 70245
rect 79480 70193 79497 70245
rect 79411 70188 79497 70193
rect 81587 70757 81673 70762
rect 81587 70705 81604 70757
rect 81656 70705 81673 70757
rect 81587 70693 81673 70705
rect 81587 70641 81604 70693
rect 81656 70641 81673 70693
rect 81587 70629 81673 70641
rect 81587 70577 81604 70629
rect 81656 70577 81673 70629
rect 81587 70565 81673 70577
rect 81587 70513 81604 70565
rect 81656 70513 81673 70565
rect 81587 70501 81673 70513
rect 81587 70449 81604 70501
rect 81656 70449 81673 70501
rect 81587 70437 81673 70449
rect 81587 70385 81604 70437
rect 81656 70385 81673 70437
rect 81587 70373 81673 70385
rect 81587 70321 81604 70373
rect 81656 70321 81673 70373
rect 81587 70309 81673 70321
rect 81587 70257 81604 70309
rect 81656 70257 81673 70309
rect 81587 70245 81673 70257
rect 81587 70193 81604 70245
rect 81656 70193 81673 70245
rect 81587 70188 81673 70193
rect 82675 70757 82761 70762
rect 82675 70705 82692 70757
rect 82744 70705 82761 70757
rect 82675 70693 82761 70705
rect 82675 70641 82692 70693
rect 82744 70641 82761 70693
rect 82675 70629 82761 70641
rect 82675 70577 82692 70629
rect 82744 70577 82761 70629
rect 82675 70565 82761 70577
rect 82675 70513 82692 70565
rect 82744 70513 82761 70565
rect 82675 70501 82761 70513
rect 82675 70449 82692 70501
rect 82744 70449 82761 70501
rect 82675 70437 82761 70449
rect 82675 70385 82692 70437
rect 82744 70385 82761 70437
rect 82675 70373 82761 70385
rect 82675 70321 82692 70373
rect 82744 70321 82761 70373
rect 82675 70309 82761 70321
rect 82675 70257 82692 70309
rect 82744 70257 82761 70309
rect 82675 70245 82761 70257
rect 82675 70193 82692 70245
rect 82744 70193 82761 70245
rect 82675 70188 82761 70193
rect 83763 70757 83849 70762
rect 83763 70705 83780 70757
rect 83832 70705 83849 70757
rect 83763 70693 83849 70705
rect 83763 70641 83780 70693
rect 83832 70641 83849 70693
rect 83763 70629 83849 70641
rect 83763 70577 83780 70629
rect 83832 70577 83849 70629
rect 83763 70565 83849 70577
rect 83763 70513 83780 70565
rect 83832 70513 83849 70565
rect 83763 70501 83849 70513
rect 83763 70449 83780 70501
rect 83832 70449 83849 70501
rect 83763 70437 83849 70449
rect 83763 70385 83780 70437
rect 83832 70385 83849 70437
rect 83763 70373 83849 70385
rect 83763 70321 83780 70373
rect 83832 70321 83849 70373
rect 83763 70309 83849 70321
rect 83763 70257 83780 70309
rect 83832 70257 83849 70309
rect 83763 70245 83849 70257
rect 83763 70193 83780 70245
rect 83832 70193 83849 70245
rect 83763 70188 83849 70193
rect 84851 70757 84937 70762
rect 84851 70705 84868 70757
rect 84920 70705 84937 70757
rect 84851 70693 84937 70705
rect 84851 70641 84868 70693
rect 84920 70641 84937 70693
rect 84851 70629 84937 70641
rect 84851 70577 84868 70629
rect 84920 70577 84937 70629
rect 84851 70565 84937 70577
rect 84851 70513 84868 70565
rect 84920 70513 84937 70565
rect 84851 70501 84937 70513
rect 84851 70449 84868 70501
rect 84920 70449 84937 70501
rect 84851 70437 84937 70449
rect 84851 70385 84868 70437
rect 84920 70385 84937 70437
rect 84851 70373 84937 70385
rect 84851 70321 84868 70373
rect 84920 70321 84937 70373
rect 84851 70309 84937 70321
rect 84851 70257 84868 70309
rect 84920 70257 84937 70309
rect 84851 70245 84937 70257
rect 84851 70193 84868 70245
rect 84920 70193 84937 70245
rect 84851 70188 84937 70193
rect 85939 70757 86025 70762
rect 85939 70705 85956 70757
rect 86008 70705 86025 70757
rect 85939 70693 86025 70705
rect 85939 70641 85956 70693
rect 86008 70641 86025 70693
rect 85939 70629 86025 70641
rect 85939 70577 85956 70629
rect 86008 70577 86025 70629
rect 85939 70565 86025 70577
rect 85939 70513 85956 70565
rect 86008 70513 86025 70565
rect 85939 70501 86025 70513
rect 85939 70449 85956 70501
rect 86008 70449 86025 70501
rect 85939 70437 86025 70449
rect 85939 70385 85956 70437
rect 86008 70385 86025 70437
rect 85939 70373 86025 70385
rect 85939 70321 85956 70373
rect 86008 70321 86025 70373
rect 85939 70309 86025 70321
rect 85939 70257 85956 70309
rect 86008 70257 86025 70309
rect 85939 70245 86025 70257
rect 85939 70193 85956 70245
rect 86008 70193 86025 70245
rect 85939 70188 86025 70193
rect 87027 70757 87113 70762
rect 87027 70705 87044 70757
rect 87096 70705 87113 70757
rect 87027 70693 87113 70705
rect 87027 70641 87044 70693
rect 87096 70641 87113 70693
rect 87027 70629 87113 70641
rect 87027 70577 87044 70629
rect 87096 70577 87113 70629
rect 87027 70565 87113 70577
rect 87027 70513 87044 70565
rect 87096 70513 87113 70565
rect 87027 70501 87113 70513
rect 87027 70449 87044 70501
rect 87096 70449 87113 70501
rect 87027 70437 87113 70449
rect 87027 70385 87044 70437
rect 87096 70385 87113 70437
rect 87027 70373 87113 70385
rect 87027 70321 87044 70373
rect 87096 70321 87113 70373
rect 87027 70309 87113 70321
rect 87027 70257 87044 70309
rect 87096 70257 87113 70309
rect 87027 70245 87113 70257
rect 87027 70193 87044 70245
rect 87096 70193 87113 70245
rect 87027 70188 87113 70193
rect 88115 70757 88201 70762
rect 88115 70705 88132 70757
rect 88184 70705 88201 70757
rect 88115 70693 88201 70705
rect 88115 70641 88132 70693
rect 88184 70641 88201 70693
rect 88115 70629 88201 70641
rect 88115 70577 88132 70629
rect 88184 70577 88201 70629
rect 88115 70565 88201 70577
rect 88115 70513 88132 70565
rect 88184 70513 88201 70565
rect 88115 70501 88201 70513
rect 88115 70449 88132 70501
rect 88184 70449 88201 70501
rect 88115 70437 88201 70449
rect 88115 70385 88132 70437
rect 88184 70385 88201 70437
rect 88115 70373 88201 70385
rect 88115 70321 88132 70373
rect 88184 70321 88201 70373
rect 88115 70309 88201 70321
rect 88115 70257 88132 70309
rect 88184 70257 88201 70309
rect 88115 70245 88201 70257
rect 88115 70193 88132 70245
rect 88184 70193 88201 70245
rect 88115 70188 88201 70193
rect 75329 69764 75413 69770
rect 75329 69712 75345 69764
rect 75397 69712 75413 69764
rect 75329 69706 75413 69712
rect 75875 69764 75959 69770
rect 75875 69712 75891 69764
rect 75943 69712 75959 69764
rect 75875 69706 75959 69712
rect 76421 69755 76505 69761
rect 76421 69703 76437 69755
rect 76489 69703 76505 69755
rect 76421 69697 76505 69703
rect 76966 69754 77050 69760
rect 76966 69702 76982 69754
rect 77034 69702 77050 69754
rect 82947 69754 83031 69760
rect 76966 69696 77050 69702
rect 78597 69742 78681 69748
rect 78597 69690 78613 69742
rect 78665 69690 78681 69742
rect 78597 69684 78681 69690
rect 79140 69739 79224 69745
rect 79140 69687 79156 69739
rect 79208 69687 79224 69739
rect 79140 69681 79224 69687
rect 79682 69738 79766 69744
rect 79682 69686 79698 69738
rect 79750 69686 79766 69738
rect 79682 69680 79766 69686
rect 80229 69743 80313 69749
rect 80229 69691 80245 69743
rect 80297 69691 80313 69743
rect 82947 69702 82963 69754
rect 83015 69702 83031 69754
rect 82947 69696 83031 69702
rect 83490 69758 83574 69764
rect 83490 69706 83506 69758
rect 83558 69706 83574 69758
rect 83490 69700 83574 69706
rect 84032 69752 84116 69758
rect 84032 69700 84048 69752
rect 84100 69700 84116 69752
rect 86213 69754 86297 69760
rect 84032 69694 84116 69700
rect 84589 69743 84673 69749
rect 80229 69685 80313 69691
rect 84589 69691 84605 69743
rect 84657 69691 84673 69743
rect 86213 69702 86229 69754
rect 86281 69702 86297 69754
rect 86213 69696 86297 69702
rect 86757 69747 86841 69753
rect 84589 69685 84673 69691
rect 86757 69695 86773 69747
rect 86825 69695 86841 69747
rect 86757 69689 86841 69695
rect 87307 69751 87391 69757
rect 87307 69699 87323 69751
rect 87375 69699 87391 69751
rect 87307 69693 87391 69699
rect 87840 69751 87924 69757
rect 87840 69699 87856 69751
rect 87908 69699 87924 69751
rect 87840 69693 87924 69699
rect 101838 69088 102410 69096
rect 101838 69036 101874 69088
rect 101926 69036 101938 69088
rect 101990 69036 102002 69088
rect 102054 69036 102066 69088
rect 102118 69036 102130 69088
rect 102182 69036 102194 69088
rect 102246 69036 102258 69088
rect 102310 69036 102322 69088
rect 102374 69036 102410 69088
rect 101838 69029 102410 69036
rect 98896 68949 98942 68970
rect 98896 68915 98902 68949
rect 98936 68915 98942 68949
rect 96641 68907 96725 68913
rect 96641 68855 96657 68907
rect 96709 68883 96725 68907
rect 96709 68855 97112 68883
rect 96641 68849 97112 68855
rect 98896 68877 98942 68915
rect 97066 68845 97112 68849
rect 97066 68839 97124 68845
rect 97066 68805 97078 68839
rect 97112 68805 97124 68839
rect 97066 68799 97124 68805
rect 97679 68800 97689 68852
rect 97741 68800 97751 68852
rect 97685 68798 97743 68800
rect 98079 68789 98089 68841
rect 98141 68789 98151 68841
rect 98236 68793 98246 68845
rect 98298 68793 98308 68845
rect 98896 68843 98902 68877
rect 98936 68843 98942 68877
rect 103378 68933 103634 68961
rect 103378 68875 103416 68933
rect 100363 68858 100421 68864
rect 100535 68858 100593 68864
rect 100707 68858 100765 68864
rect 100879 68858 100937 68864
rect 101051 68858 101109 68864
rect 101256 68858 101314 68864
rect 101433 68858 101491 68864
rect 101605 68858 101663 68864
rect 101777 68858 101835 68864
rect 101949 68858 102007 68864
rect 102121 68858 102179 68864
rect 102293 68858 102351 68864
rect 102958 68858 103416 68875
rect 98896 68805 98942 68843
rect 97210 68758 97268 68764
rect 97210 68724 97222 68758
rect 97256 68724 97268 68758
rect 97978 68732 97988 68784
rect 98040 68732 98050 68784
rect 98896 68771 98902 68805
rect 98936 68775 98942 68805
rect 100091 68808 100138 68852
rect 100363 68824 100375 68858
rect 100409 68824 100547 68858
rect 100581 68824 100719 68858
rect 100753 68824 100891 68858
rect 100925 68824 101063 68858
rect 101097 68824 101268 68858
rect 101302 68824 101445 68858
rect 101479 68824 101617 68858
rect 101651 68824 101789 68858
rect 101823 68824 101961 68858
rect 101995 68824 102133 68858
rect 102167 68824 102305 68858
rect 102339 68824 103416 68858
rect 100363 68818 100421 68824
rect 100535 68818 100593 68824
rect 100707 68818 100765 68824
rect 100879 68818 100937 68824
rect 101051 68818 101109 68824
rect 101256 68818 101314 68824
rect 101433 68818 101491 68824
rect 101605 68818 101663 68824
rect 101777 68818 101835 68824
rect 101949 68818 102007 68824
rect 102121 68818 102179 68824
rect 102293 68818 102351 68824
rect 102958 68811 103416 68824
rect 98936 68771 100042 68775
rect 98896 68769 100042 68771
rect 98896 68735 99633 68769
rect 99667 68735 99705 68769
rect 99739 68735 99777 68769
rect 99811 68735 99849 68769
rect 99883 68735 99921 68769
rect 99955 68735 99993 68769
rect 100027 68735 100042 68769
rect 98896 68733 100042 68735
rect 97210 68723 97268 68724
rect 96641 68718 97268 68723
rect 96641 68717 97256 68718
rect 96641 68665 96657 68717
rect 96709 68689 97256 68717
rect 98896 68699 98902 68733
rect 98936 68730 100042 68733
rect 98936 68699 98942 68730
rect 99619 68729 100042 68730
rect 100091 68774 100097 68808
rect 100131 68778 100138 68808
rect 100131 68774 100601 68778
rect 100091 68772 100601 68774
rect 100091 68738 100371 68772
rect 100405 68738 100443 68772
rect 100477 68738 100601 68772
rect 100091 68736 100601 68738
rect 96709 68665 96725 68689
rect 96641 68659 96725 68665
rect 98896 68661 98942 68699
rect 98896 68627 98902 68661
rect 98936 68627 98942 68661
rect 100091 68702 100097 68736
rect 100131 68732 100601 68736
rect 103378 68753 103416 68811
rect 103596 68753 103634 68933
rect 100131 68702 100138 68732
rect 103378 68725 103634 68753
rect 100091 68658 100138 68702
rect 98896 68606 98942 68627
rect 98600 68542 98978 68549
rect 98600 68490 98635 68542
rect 98687 68490 98699 68542
rect 98751 68490 98763 68542
rect 98815 68490 98827 68542
rect 98879 68490 98891 68542
rect 98943 68490 98978 68542
rect 98600 68484 98978 68490
rect 101850 67937 102397 67947
rect 101850 67885 101873 67937
rect 101925 67885 101937 67937
rect 101989 67885 102001 67937
rect 102053 67885 102065 67937
rect 102117 67885 102129 67937
rect 102181 67885 102193 67937
rect 102245 67885 102257 67937
rect 102309 67885 102321 67937
rect 102373 67885 102397 67937
rect 101850 67876 102397 67885
rect 98896 67799 98942 67820
rect 98896 67765 98902 67799
rect 98936 67765 98942 67799
rect 96641 67757 96725 67763
rect 96641 67705 96657 67757
rect 96709 67733 96725 67757
rect 96709 67705 97112 67733
rect 96641 67699 97112 67705
rect 98896 67727 98942 67765
rect 97066 67695 97112 67699
rect 97066 67689 97124 67695
rect 97066 67655 97078 67689
rect 97112 67655 97124 67689
rect 97066 67649 97124 67655
rect 97679 67650 97689 67702
rect 97741 67650 97751 67702
rect 97685 67648 97743 67650
rect 98079 67639 98089 67691
rect 98141 67639 98151 67691
rect 98236 67643 98246 67695
rect 98298 67643 98308 67695
rect 98896 67693 98902 67727
rect 98936 67693 98942 67727
rect 103366 67782 103622 67810
rect 103366 67725 103404 67782
rect 100363 67708 100421 67714
rect 100535 67708 100593 67714
rect 100707 67708 100765 67714
rect 100879 67708 100937 67714
rect 101051 67708 101109 67714
rect 101256 67708 101314 67714
rect 101433 67708 101491 67714
rect 101605 67708 101663 67714
rect 101777 67708 101835 67714
rect 101949 67708 102007 67714
rect 102121 67708 102179 67714
rect 102293 67708 102351 67714
rect 102958 67708 103404 67725
rect 98896 67655 98942 67693
rect 97210 67608 97268 67614
rect 97210 67574 97222 67608
rect 97256 67574 97268 67608
rect 97978 67582 97988 67634
rect 98040 67582 98050 67634
rect 98896 67621 98902 67655
rect 98936 67625 98942 67655
rect 100091 67658 100138 67702
rect 100363 67674 100375 67708
rect 100409 67674 100547 67708
rect 100581 67674 100719 67708
rect 100753 67674 100891 67708
rect 100925 67674 101063 67708
rect 101097 67674 101268 67708
rect 101302 67674 101445 67708
rect 101479 67674 101617 67708
rect 101651 67674 101789 67708
rect 101823 67674 101961 67708
rect 101995 67674 102133 67708
rect 102167 67674 102305 67708
rect 102339 67674 103404 67708
rect 100363 67668 100421 67674
rect 100535 67668 100593 67674
rect 100707 67668 100765 67674
rect 100879 67668 100937 67674
rect 101051 67668 101109 67674
rect 101256 67668 101314 67674
rect 101433 67668 101491 67674
rect 101605 67668 101663 67674
rect 101777 67668 101835 67674
rect 101949 67668 102007 67674
rect 102121 67668 102179 67674
rect 102293 67668 102351 67674
rect 102958 67661 103404 67674
rect 98936 67621 100042 67625
rect 98896 67619 100042 67621
rect 98896 67585 99633 67619
rect 99667 67585 99705 67619
rect 99739 67585 99777 67619
rect 99811 67585 99849 67619
rect 99883 67585 99921 67619
rect 99955 67585 99993 67619
rect 100027 67585 100042 67619
rect 98896 67583 100042 67585
rect 97210 67573 97268 67574
rect 96641 67568 97268 67573
rect 96641 67567 97256 67568
rect 96641 67515 96657 67567
rect 96709 67539 97256 67567
rect 98896 67549 98902 67583
rect 98936 67580 100042 67583
rect 98936 67549 98942 67580
rect 99619 67579 100042 67580
rect 100091 67624 100097 67658
rect 100131 67628 100138 67658
rect 100131 67624 100601 67628
rect 100091 67622 100601 67624
rect 100091 67588 100371 67622
rect 100405 67588 100443 67622
rect 100477 67588 100601 67622
rect 100091 67586 100601 67588
rect 96709 67515 96725 67539
rect 96641 67509 96725 67515
rect 98896 67511 98942 67549
rect 98896 67477 98902 67511
rect 98936 67477 98942 67511
rect 100091 67552 100097 67586
rect 100131 67582 100601 67586
rect 103366 67602 103404 67661
rect 103584 67602 103622 67782
rect 100131 67552 100138 67582
rect 103366 67574 103622 67602
rect 100091 67508 100138 67552
rect 98896 67456 98942 67477
rect 98598 67392 98976 67399
rect 98598 67340 98633 67392
rect 98685 67340 98697 67392
rect 98749 67340 98761 67392
rect 98813 67340 98825 67392
rect 98877 67340 98889 67392
rect 98941 67340 98976 67392
rect 98598 67334 98976 67340
rect 101840 65395 102387 65405
rect 101840 65343 101863 65395
rect 101915 65343 101927 65395
rect 101979 65343 101991 65395
rect 102043 65343 102055 65395
rect 102107 65343 102119 65395
rect 102171 65343 102183 65395
rect 102235 65343 102247 65395
rect 102299 65343 102311 65395
rect 102363 65343 102387 65395
rect 101840 65334 102387 65343
rect 98896 65259 98942 65280
rect 98896 65225 98902 65259
rect 98936 65225 98942 65259
rect 96641 65217 96725 65223
rect 96641 65165 96657 65217
rect 96709 65193 96725 65217
rect 96709 65165 97112 65193
rect 96641 65159 97112 65165
rect 98896 65187 98942 65225
rect 97066 65155 97112 65159
rect 97066 65149 97124 65155
rect 97066 65115 97078 65149
rect 97112 65115 97124 65149
rect 97066 65109 97124 65115
rect 97679 65110 97689 65162
rect 97741 65110 97751 65162
rect 97685 65108 97743 65110
rect 98079 65099 98089 65151
rect 98141 65099 98151 65151
rect 98236 65103 98246 65155
rect 98298 65103 98308 65155
rect 98896 65153 98902 65187
rect 98936 65153 98942 65187
rect 103224 65250 103480 65278
rect 103224 65184 103262 65250
rect 100363 65168 100421 65174
rect 100535 65168 100593 65174
rect 100707 65168 100765 65174
rect 100879 65168 100937 65174
rect 101051 65168 101109 65174
rect 101256 65168 101314 65174
rect 101433 65168 101491 65174
rect 101605 65168 101663 65174
rect 101777 65168 101835 65174
rect 101949 65168 102007 65174
rect 102121 65168 102179 65174
rect 102293 65168 102351 65174
rect 102958 65168 103262 65184
rect 98896 65115 98942 65153
rect 97210 65068 97268 65074
rect 97210 65034 97222 65068
rect 97256 65034 97268 65068
rect 97978 65042 97988 65094
rect 98040 65042 98050 65094
rect 98896 65081 98902 65115
rect 98936 65085 98942 65115
rect 100091 65118 100138 65162
rect 100363 65134 100375 65168
rect 100409 65134 100547 65168
rect 100581 65134 100719 65168
rect 100753 65134 100891 65168
rect 100925 65134 101063 65168
rect 101097 65134 101268 65168
rect 101302 65134 101445 65168
rect 101479 65134 101617 65168
rect 101651 65134 101789 65168
rect 101823 65134 101961 65168
rect 101995 65134 102133 65168
rect 102167 65134 102305 65168
rect 102339 65134 103262 65168
rect 100363 65128 100421 65134
rect 100535 65128 100593 65134
rect 100707 65128 100765 65134
rect 100879 65128 100937 65134
rect 101051 65128 101109 65134
rect 101256 65128 101314 65134
rect 101433 65128 101491 65134
rect 101605 65128 101663 65134
rect 101777 65128 101835 65134
rect 101949 65128 102007 65134
rect 102121 65128 102179 65134
rect 102293 65128 102351 65134
rect 102958 65120 103262 65134
rect 98936 65081 100042 65085
rect 98896 65079 100042 65081
rect 98896 65045 99633 65079
rect 99667 65045 99705 65079
rect 99739 65045 99777 65079
rect 99811 65045 99849 65079
rect 99883 65045 99921 65079
rect 99955 65045 99993 65079
rect 100027 65045 100042 65079
rect 98896 65043 100042 65045
rect 97210 65033 97268 65034
rect 96641 65028 97268 65033
rect 96641 65027 97256 65028
rect 96641 64975 96657 65027
rect 96709 64999 97256 65027
rect 98896 65009 98902 65043
rect 98936 65040 100042 65043
rect 98936 65009 98942 65040
rect 99619 65039 100042 65040
rect 100091 65084 100097 65118
rect 100131 65088 100138 65118
rect 100131 65084 100601 65088
rect 100091 65082 100601 65084
rect 100091 65048 100371 65082
rect 100405 65048 100443 65082
rect 100477 65048 100601 65082
rect 100091 65046 100601 65048
rect 96709 64975 96725 64999
rect 96641 64969 96725 64975
rect 98896 64971 98942 65009
rect 98896 64937 98902 64971
rect 98936 64937 98942 64971
rect 100091 65012 100097 65046
rect 100131 65042 100601 65046
rect 103224 65070 103262 65120
rect 103442 65070 103480 65250
rect 103224 65042 103480 65070
rect 100131 65012 100138 65042
rect 100091 64968 100138 65012
rect 98896 64916 98942 64937
rect 98516 64851 98894 64858
rect 98516 64799 98551 64851
rect 98603 64799 98615 64851
rect 98667 64799 98679 64851
rect 98731 64799 98743 64851
rect 98795 64799 98807 64851
rect 98859 64799 98894 64851
rect 98516 64793 98894 64799
rect 101840 64125 102387 64135
rect 101840 64073 101863 64125
rect 101915 64073 101927 64125
rect 101979 64073 101991 64125
rect 102043 64073 102055 64125
rect 102107 64073 102119 64125
rect 102171 64073 102183 64125
rect 102235 64073 102247 64125
rect 102299 64073 102311 64125
rect 102363 64073 102387 64125
rect 101840 64064 102387 64073
rect 98896 63989 98942 64010
rect 98896 63955 98902 63989
rect 98936 63955 98942 63989
rect 96641 63947 96725 63953
rect 96641 63895 96657 63947
rect 96709 63923 96725 63947
rect 96709 63895 97112 63923
rect 96641 63889 97112 63895
rect 98896 63917 98942 63955
rect 97066 63885 97112 63889
rect 97066 63879 97124 63885
rect 97066 63845 97078 63879
rect 97112 63845 97124 63879
rect 97066 63839 97124 63845
rect 97679 63840 97689 63892
rect 97741 63840 97751 63892
rect 97685 63838 97743 63840
rect 98079 63829 98089 63881
rect 98141 63829 98151 63881
rect 98236 63833 98246 63885
rect 98298 63833 98308 63885
rect 98896 63883 98902 63917
rect 98936 63883 98942 63917
rect 103195 63960 103451 63988
rect 103195 63914 103233 63960
rect 100363 63898 100421 63904
rect 100535 63898 100593 63904
rect 100707 63898 100765 63904
rect 100879 63898 100937 63904
rect 101051 63898 101109 63904
rect 101256 63898 101314 63904
rect 101433 63898 101491 63904
rect 101605 63898 101663 63904
rect 101777 63898 101835 63904
rect 101949 63898 102007 63904
rect 102121 63898 102179 63904
rect 102293 63898 102351 63904
rect 102958 63898 103233 63914
rect 98896 63845 98942 63883
rect 97210 63798 97268 63804
rect 97210 63764 97222 63798
rect 97256 63764 97268 63798
rect 97978 63772 97988 63824
rect 98040 63772 98050 63824
rect 98896 63811 98902 63845
rect 98936 63815 98942 63845
rect 100091 63848 100138 63892
rect 100363 63864 100375 63898
rect 100409 63864 100547 63898
rect 100581 63864 100719 63898
rect 100753 63864 100891 63898
rect 100925 63864 101063 63898
rect 101097 63864 101268 63898
rect 101302 63864 101445 63898
rect 101479 63864 101617 63898
rect 101651 63864 101789 63898
rect 101823 63864 101961 63898
rect 101995 63864 102133 63898
rect 102167 63864 102305 63898
rect 102339 63864 103233 63898
rect 100363 63858 100421 63864
rect 100535 63858 100593 63864
rect 100707 63858 100765 63864
rect 100879 63858 100937 63864
rect 101051 63858 101109 63864
rect 101256 63858 101314 63864
rect 101433 63858 101491 63864
rect 101605 63858 101663 63864
rect 101777 63858 101835 63864
rect 101949 63858 102007 63864
rect 102121 63858 102179 63864
rect 102293 63858 102351 63864
rect 102958 63850 103233 63864
rect 98936 63811 100042 63815
rect 98896 63809 100042 63811
rect 98896 63775 99633 63809
rect 99667 63775 99705 63809
rect 99739 63775 99777 63809
rect 99811 63775 99849 63809
rect 99883 63775 99921 63809
rect 99955 63775 99993 63809
rect 100027 63775 100042 63809
rect 98896 63773 100042 63775
rect 97210 63763 97268 63764
rect 96641 63758 97268 63763
rect 96641 63757 97256 63758
rect 96641 63705 96657 63757
rect 96709 63729 97256 63757
rect 98896 63739 98902 63773
rect 98936 63770 100042 63773
rect 98936 63739 98942 63770
rect 99619 63769 100042 63770
rect 100091 63814 100097 63848
rect 100131 63818 100138 63848
rect 100131 63814 100601 63818
rect 100091 63812 100601 63814
rect 100091 63778 100371 63812
rect 100405 63778 100443 63812
rect 100477 63778 100601 63812
rect 100091 63776 100601 63778
rect 96709 63705 96725 63729
rect 96641 63699 96725 63705
rect 98896 63701 98942 63739
rect 98896 63667 98902 63701
rect 98936 63667 98942 63701
rect 100091 63742 100097 63776
rect 100131 63772 100601 63776
rect 103195 63780 103233 63850
rect 103413 63780 103451 63960
rect 100131 63742 100138 63772
rect 103195 63752 103451 63780
rect 100091 63698 100138 63742
rect 98896 63646 98942 63667
rect 98514 63582 98892 63589
rect 98514 63530 98549 63582
rect 98601 63530 98613 63582
rect 98665 63530 98677 63582
rect 98729 63530 98741 63582
rect 98793 63530 98805 63582
rect 98857 63530 98892 63582
rect 98514 63524 98892 63530
rect 64166 63204 64422 63232
rect 64166 63024 64204 63204
rect 64384 63024 64422 63204
rect 64166 62996 64422 63024
rect 69626 63204 69882 63232
rect 69626 63024 69664 63204
rect 69844 63024 69882 63204
rect 69626 62996 69882 63024
rect 69754 62986 69872 62996
rect 64330 62177 64394 62190
rect 64320 62171 64404 62177
rect 64320 62119 64336 62171
rect 64388 62119 64404 62171
rect 64320 62113 64404 62119
rect 62513 61223 62597 61229
rect 62513 61171 62529 61223
rect 62581 61171 62597 61223
rect 62513 61165 62597 61171
rect 63785 61223 63869 61229
rect 63785 61171 63801 61223
rect 63853 61171 63869 61223
rect 63785 61165 63869 61171
rect 60666 60110 60915 60116
rect 60666 60058 60700 60110
rect 60752 60058 60764 60110
rect 60816 60058 60828 60110
rect 60880 60058 60915 60110
rect 60666 60052 60915 60058
rect 62139 60109 62455 60126
rect 62139 60057 62175 60109
rect 62227 60057 62239 60109
rect 62291 60057 62303 60109
rect 62355 60057 62367 60109
rect 62419 60057 62455 60109
rect 62139 60040 62455 60057
rect 62523 59967 62587 61165
rect 64330 60129 64394 62113
rect 66512 61667 66596 61673
rect 66512 61615 66528 61667
rect 66580 61615 66596 61667
rect 66512 61609 66596 61615
rect 62658 60110 62905 60119
rect 62658 60058 62691 60110
rect 62743 60058 62755 60110
rect 62807 60058 62819 60110
rect 62871 60058 62905 60110
rect 62658 60049 62905 60058
rect 64020 60102 64261 60111
rect 64020 60050 64050 60102
rect 64102 60050 64114 60102
rect 64166 60050 64178 60102
rect 64230 60050 64261 60102
rect 64467 60109 64785 60116
rect 64467 60057 64504 60109
rect 64556 60057 64568 60109
rect 64620 60057 64632 60109
rect 64684 60057 64696 60109
rect 64748 60057 64785 60109
rect 64467 60050 64785 60057
rect 66005 60108 66452 60115
rect 66005 60056 66042 60108
rect 66094 60056 66106 60108
rect 66158 60056 66170 60108
rect 66222 60056 66234 60108
rect 66286 60056 66298 60108
rect 66350 60056 66362 60108
rect 66414 60056 66452 60108
rect 66005 60050 66452 60056
rect 64020 60042 64261 60050
rect 66522 59962 66586 61609
rect 66659 60105 66906 60113
rect 66659 60053 66692 60105
rect 66744 60053 66756 60105
rect 66808 60053 66820 60105
rect 66872 60053 66906 60105
rect 66659 60045 66906 60053
rect 62514 59036 62598 59042
rect 62514 58984 62530 59036
rect 62582 58984 62598 59036
rect 62514 58978 62598 58984
rect 64326 59034 64410 59040
rect 64326 58982 64342 59034
rect 64394 58982 64410 59034
rect 64326 58976 64410 58982
rect 60960 58802 61972 58866
rect 64948 58803 65967 58867
rect 60839 57872 60891 58676
rect 60829 57820 60839 57872
rect 60891 57820 60901 57872
rect 50105 57143 50152 57195
rect 50204 57143 50233 57195
rect 50105 55833 50233 57143
rect 50095 55827 50243 55833
rect 50095 55775 50111 55827
rect 50163 55775 50175 55827
rect 50227 55775 50243 55827
rect 50095 55769 50243 55775
rect 50105 55734 50233 55769
rect 61448 54454 61512 58802
rect 62514 58441 62598 58447
rect 62514 58389 62530 58441
rect 62582 58389 62598 58441
rect 62514 58383 62598 58389
rect 64326 58441 64410 58447
rect 64326 58389 64342 58441
rect 64394 58389 64410 58441
rect 64326 58383 64410 58389
rect 62524 57583 62588 58383
rect 64336 58350 64400 58383
rect 64336 58286 64586 58350
rect 64522 57591 64586 58286
rect 64512 57585 64596 57591
rect 62514 57577 62598 57583
rect 62514 57525 62530 57577
rect 62582 57525 62598 57577
rect 64512 57533 64528 57585
rect 64580 57533 64596 57585
rect 64512 57527 64596 57533
rect 62514 57519 62598 57525
rect 62524 57502 62588 57519
rect 65422 54459 65486 58803
rect 66839 57872 66891 58684
rect 66829 57820 66839 57872
rect 66891 57820 66901 57872
rect 66839 57817 66891 57820
rect 61438 54448 61522 54454
rect 61438 54396 61454 54448
rect 61506 54396 61522 54448
rect 61438 54390 61522 54396
rect 65412 54453 65496 54459
rect 65412 54401 65428 54453
rect 65480 54401 65496 54453
rect 65412 54395 65496 54401
rect 47687 54321 47835 54327
rect 47687 54269 47703 54321
rect 47755 54269 47767 54321
rect 47819 54269 47835 54321
rect 47687 54263 47835 54269
rect 47696 54223 47824 54263
rect 44391 53768 44475 53774
rect 44391 53716 44407 53768
rect 44459 53716 44475 53768
rect 44391 53710 44475 53716
rect 43615 53345 43699 53351
rect 26885 53303 38710 53310
rect 26885 53187 26901 53303
rect 27017 53187 38577 53303
rect 38693 53187 38710 53303
rect 43615 53293 43631 53345
rect 43683 53293 43699 53345
rect 43615 53287 43699 53293
rect 26885 53181 38710 53187
rect 65044 52862 65128 52868
rect 59035 52824 59183 52830
rect 59035 52772 59051 52824
rect 59103 52772 59115 52824
rect 59167 52772 59183 52824
rect 65044 52810 65060 52862
rect 65112 52810 65128 52862
rect 65044 52804 65128 52810
rect 59035 52766 59183 52772
rect 59045 52666 59173 52766
rect 45206 52624 59173 52666
rect 45206 52572 51014 52624
rect 51066 52572 51078 52624
rect 51130 52572 59173 52624
rect 45206 52538 59173 52572
rect 60462 52611 60590 52649
rect 60462 52559 60499 52611
rect 60551 52559 60590 52611
rect 41372 52111 41491 52120
rect 41372 52059 41405 52111
rect 41457 52059 41491 52111
rect 41372 52047 41491 52059
rect 41372 51995 41405 52047
rect 41457 51995 41491 52047
rect 43101 52036 43111 52088
rect 43163 52036 43400 52088
rect 44695 52081 44788 52098
rect 41372 51983 41491 51995
rect 26054 51945 37850 51952
rect 26054 51829 26070 51945
rect 26186 51829 37717 51945
rect 37833 51829 37850 51945
rect 26054 51823 37850 51829
rect 41372 51931 41405 51983
rect 41457 51931 41491 51983
rect 41372 51919 41491 51931
rect 41372 51867 41405 51919
rect 41457 51867 41491 51919
rect 41372 51855 41491 51867
rect 41372 51803 41405 51855
rect 41457 51803 41491 51855
rect 41372 51791 41491 51803
rect 41372 51739 41405 51791
rect 41457 51739 41491 51791
rect 41372 51727 41491 51739
rect 41372 51675 41405 51727
rect 41457 51675 41491 51727
rect 44695 52029 44715 52081
rect 44767 52029 44788 52081
rect 44695 52017 44788 52029
rect 44695 51965 44715 52017
rect 44767 51965 44788 52017
rect 44695 51953 44788 51965
rect 44695 51901 44715 51953
rect 44767 51901 44788 51953
rect 44695 51889 44788 51901
rect 44695 51837 44715 51889
rect 44767 51837 44788 51889
rect 44695 51825 44788 51837
rect 44695 51773 44715 51825
rect 44767 51773 44788 51825
rect 44695 51761 44788 51773
rect 44695 51709 44715 51761
rect 44767 51709 44788 51761
rect 44695 51692 44788 51709
rect 41372 51667 41491 51675
rect 39449 51660 39597 51666
rect 38768 51597 38832 51622
rect 38758 51591 38842 51597
rect 38758 51539 38774 51591
rect 38826 51539 38842 51591
rect 38758 51533 38842 51539
rect 39449 51544 39465 51660
rect 39581 51590 39597 51660
rect 45206 51656 45334 52538
rect 44888 51601 45334 51656
rect 39581 51544 39760 51590
rect 39449 51538 39760 51544
rect 42178 51541 42188 51593
rect 42240 51541 43475 51593
rect 44603 51537 45334 51601
rect 38768 51120 38832 51533
rect 44888 51528 45334 51537
rect 44690 51424 44807 51449
rect 44690 51372 44722 51424
rect 44774 51372 44807 51424
rect 44690 51360 44807 51372
rect 44690 51308 44722 51360
rect 44774 51308 44807 51360
rect 44690 51296 44807 51308
rect 42680 51229 42690 51281
rect 42742 51229 43366 51281
rect 44690 51244 44722 51296
rect 44774 51244 44807 51296
rect 44690 51220 44807 51244
rect 38758 51114 38842 51120
rect 38758 51062 38774 51114
rect 38826 51062 38842 51114
rect 41855 51104 42188 51105
rect 38758 51056 38842 51062
rect 38203 50776 38287 50782
rect 38203 50724 38219 50776
rect 38271 50724 38287 50776
rect 38203 50718 38287 50724
rect 18894 50610 22248 50633
rect 18894 50558 18913 50610
rect 18965 50558 18977 50610
rect 19029 50558 19041 50610
rect 19093 50558 19105 50610
rect 19157 50558 19169 50610
rect 19221 50558 19233 50610
rect 19285 50558 19297 50610
rect 19349 50558 19361 50610
rect 19413 50558 19425 50610
rect 19477 50558 19489 50610
rect 19541 50558 19553 50610
rect 19605 50558 19617 50610
rect 19669 50558 19681 50610
rect 19733 50558 19745 50610
rect 19797 50558 19809 50610
rect 19861 50558 19873 50610
rect 19925 50558 19937 50610
rect 19989 50558 20001 50610
rect 20053 50558 20065 50610
rect 20117 50558 20129 50610
rect 20181 50558 20193 50610
rect 20245 50558 20257 50610
rect 20309 50558 20321 50610
rect 20373 50558 20385 50610
rect 20437 50558 20449 50610
rect 20501 50558 20513 50610
rect 20565 50558 20577 50610
rect 20629 50558 20641 50610
rect 20693 50558 20705 50610
rect 20757 50558 20769 50610
rect 20821 50558 20833 50610
rect 20885 50558 20897 50610
rect 20949 50558 20961 50610
rect 21013 50558 21025 50610
rect 21077 50558 21089 50610
rect 21141 50558 21153 50610
rect 21205 50558 21217 50610
rect 21269 50558 21281 50610
rect 21333 50558 21345 50610
rect 21397 50558 21409 50610
rect 21461 50558 21473 50610
rect 21525 50558 21537 50610
rect 21589 50558 21601 50610
rect 21653 50558 21665 50610
rect 21717 50558 21729 50610
rect 21781 50558 21793 50610
rect 21845 50558 21857 50610
rect 21909 50558 21921 50610
rect 21973 50558 21985 50610
rect 22037 50558 22049 50610
rect 22101 50558 22113 50610
rect 22165 50558 22177 50610
rect 22229 50558 22248 50610
rect 18894 50536 22248 50558
rect 38213 49999 38277 50718
rect 38202 49993 38286 49999
rect 38202 49941 38218 49993
rect 38270 49941 38286 49993
rect 38202 49935 38286 49941
rect 31635 49472 31735 49504
rect 31635 49420 31659 49472
rect 31711 49420 31735 49472
rect 31635 49408 31735 49420
rect 31635 49356 31659 49408
rect 31711 49356 31735 49408
rect 31635 49344 31735 49356
rect 31635 49292 31659 49344
rect 31711 49292 31735 49344
rect 31635 49280 31735 49292
rect 31635 49228 31659 49280
rect 31711 49228 31735 49280
rect 31635 49197 31735 49228
rect 16491 49165 16747 49193
rect 16491 48985 16529 49165
rect 16709 49134 16747 49165
rect 16709 49128 30411 49134
rect 16709 49012 24109 49128
rect 24225 49012 30411 49128
rect 16709 49006 30411 49012
rect 31759 49006 32972 49134
rect 16709 48985 16747 49006
rect 16491 48957 16747 48985
rect 31632 48941 31739 48967
rect 31632 48889 31659 48941
rect 31711 48889 31739 48941
rect 31632 48877 31739 48889
rect 31632 48825 31659 48877
rect 31711 48825 31739 48877
rect 31632 48813 31739 48825
rect 31632 48761 31659 48813
rect 31711 48761 31739 48813
rect 31632 48736 31739 48761
rect 18902 47602 22252 47627
rect 18902 47550 18919 47602
rect 18971 47550 18983 47602
rect 19035 47550 19047 47602
rect 19099 47550 19111 47602
rect 19163 47550 19175 47602
rect 19227 47550 19239 47602
rect 19291 47550 19303 47602
rect 19355 47550 19367 47602
rect 19419 47550 19431 47602
rect 19483 47550 19495 47602
rect 19547 47550 19559 47602
rect 19611 47550 19623 47602
rect 19675 47550 19687 47602
rect 19739 47550 19751 47602
rect 19803 47550 19815 47602
rect 19867 47550 19879 47602
rect 19931 47550 19943 47602
rect 19995 47550 20007 47602
rect 20059 47550 20071 47602
rect 20123 47550 20135 47602
rect 20187 47550 20199 47602
rect 20251 47550 20263 47602
rect 20315 47550 20327 47602
rect 20379 47550 20391 47602
rect 20443 47550 20455 47602
rect 20507 47550 20519 47602
rect 20571 47550 20583 47602
rect 20635 47550 20647 47602
rect 20699 47550 20711 47602
rect 20763 47550 20775 47602
rect 20827 47550 20839 47602
rect 20891 47550 20903 47602
rect 20955 47550 20967 47602
rect 21019 47550 21031 47602
rect 21083 47550 21095 47602
rect 21147 47550 21159 47602
rect 21211 47550 21223 47602
rect 21275 47550 21287 47602
rect 21339 47550 21351 47602
rect 21403 47550 21415 47602
rect 21467 47550 21479 47602
rect 21531 47550 21543 47602
rect 21595 47550 21607 47602
rect 21659 47550 21671 47602
rect 21723 47550 21735 47602
rect 21787 47550 21799 47602
rect 21851 47550 21863 47602
rect 21915 47550 21927 47602
rect 21979 47550 21991 47602
rect 22043 47550 22055 47602
rect 22107 47550 22119 47602
rect 22171 47550 22183 47602
rect 22235 47550 22252 47602
rect 18902 47525 22252 47550
rect 32844 45724 32972 49006
rect 38213 48140 38277 49935
rect 38768 48479 38832 51056
rect 41852 51053 42188 51104
rect 42240 51053 42250 51105
rect 39828 50776 39912 50782
rect 39828 50724 39844 50776
rect 39896 50724 39912 50776
rect 39828 50718 39912 50724
rect 45182 50604 47216 50610
rect 45182 50552 47084 50604
rect 47136 50552 47148 50604
rect 47200 50552 47216 50604
rect 45182 50546 47216 50552
rect 39449 50431 39760 50437
rect 43101 50436 43111 50488
rect 43163 50436 43372 50488
rect 44688 50479 44803 50508
rect 39449 50315 39465 50431
rect 39581 50385 39760 50431
rect 44688 50427 44719 50479
rect 44771 50427 44803 50479
rect 44688 50415 44803 50427
rect 39581 50315 39597 50385
rect 39449 50309 39597 50315
rect 44688 50363 44719 50415
rect 44771 50363 44803 50415
rect 44688 50351 44803 50363
rect 41359 50274 41468 50303
rect 41359 50222 41387 50274
rect 41439 50222 41468 50274
rect 41359 50210 41468 50222
rect 41359 50158 41387 50210
rect 41439 50158 41468 50210
rect 41359 50146 41468 50158
rect 41359 50094 41387 50146
rect 41439 50094 41468 50146
rect 41359 50066 41468 50094
rect 44688 50299 44719 50351
rect 44771 50299 44803 50351
rect 44688 50287 44803 50299
rect 44688 50235 44719 50287
rect 44771 50235 44803 50287
rect 44688 50223 44803 50235
rect 44688 50171 44719 50223
rect 44771 50171 44803 50223
rect 44688 50159 44803 50171
rect 44688 50107 44719 50159
rect 44771 50107 44803 50159
rect 44688 50079 44803 50107
rect 45182 50000 45246 50546
rect 42178 49937 42188 49989
rect 42240 49937 43470 49989
rect 44616 49936 45246 50000
rect 44700 49825 44783 49845
rect 59046 49842 59174 49847
rect 44700 49773 44715 49825
rect 44767 49773 44783 49825
rect 59036 49836 59184 49842
rect 59036 49784 59052 49836
rect 59104 49784 59116 49836
rect 59168 49784 59184 49836
rect 59036 49778 59184 49784
rect 44700 49761 44783 49773
rect 44700 49709 44715 49761
rect 44767 49709 44783 49761
rect 44700 49697 44783 49709
rect 42680 49629 42690 49681
rect 42742 49629 43353 49681
rect 44700 49645 44715 49697
rect 44767 49645 44783 49697
rect 44700 49626 44783 49645
rect 59046 49470 59174 49778
rect 41357 49440 41472 49469
rect 41357 49388 41388 49440
rect 41440 49388 41472 49440
rect 41357 49376 41472 49388
rect 41357 49324 41388 49376
rect 41440 49324 41472 49376
rect 41357 49312 41472 49324
rect 41357 49260 41388 49312
rect 41440 49260 41472 49312
rect 41357 49248 41472 49260
rect 41357 49196 41388 49248
rect 41440 49196 41472 49248
rect 41357 49184 41472 49196
rect 41357 49132 41388 49184
rect 41440 49132 41472 49184
rect 41357 49120 41472 49132
rect 41357 49068 41388 49120
rect 41440 49068 41472 49120
rect 41357 49040 41472 49068
rect 45208 49430 59174 49470
rect 45208 49378 53599 49430
rect 53651 49378 53663 49430
rect 53715 49378 59174 49430
rect 45208 49342 59174 49378
rect 39449 49018 39597 49024
rect 39449 48902 39465 49018
rect 39581 48948 39597 49018
rect 39581 48902 39755 48948
rect 39449 48896 39755 48902
rect 43101 48836 43111 48888
rect 43163 48836 43345 48888
rect 44691 48729 44776 48734
rect 44691 48677 44707 48729
rect 44759 48677 44776 48729
rect 44691 48665 44776 48677
rect 44691 48613 44707 48665
rect 44759 48613 44776 48665
rect 44691 48601 44776 48613
rect 44691 48549 44707 48601
rect 44759 48549 44776 48601
rect 44691 48537 44776 48549
rect 44691 48485 44707 48537
rect 44759 48485 44776 48537
rect 44691 48480 44776 48485
rect 38758 48473 38842 48479
rect 38758 48421 38774 48473
rect 38826 48421 38842 48473
rect 38758 48415 38842 48421
rect 41892 48411 42186 48463
rect 42238 48411 42244 48463
rect 45208 48430 45336 49342
rect 42186 48391 42244 48411
rect 44896 48398 45336 48430
rect 42186 48339 43474 48391
rect 44625 48334 45336 48398
rect 44896 48302 45336 48334
rect 44686 48233 44788 48261
rect 44686 48181 44711 48233
rect 44763 48181 44788 48233
rect 44686 48169 44788 48181
rect 38203 48134 38287 48140
rect 38203 48082 38219 48134
rect 38271 48082 38287 48134
rect 38203 48076 38287 48082
rect 39821 48134 39905 48140
rect 39821 48082 39837 48134
rect 39889 48082 39905 48134
rect 39821 48076 39905 48082
rect 44686 48117 44711 48169
rect 44763 48117 44788 48169
rect 44686 48105 44788 48117
rect 42680 48029 42690 48081
rect 42742 48029 43361 48081
rect 44686 48053 44711 48105
rect 44763 48053 44788 48105
rect 44686 48025 44788 48053
rect 60462 48117 60590 52559
rect 65054 49842 65118 52804
rect 66460 52608 66588 52654
rect 66460 52556 66499 52608
rect 66551 52556 66588 52608
rect 65044 49836 65128 49842
rect 65044 49784 65060 49836
rect 65112 49784 65128 49836
rect 65044 49778 65128 49784
rect 62799 48598 62887 48616
rect 62799 48546 62817 48598
rect 62869 48546 62887 48598
rect 62799 48534 62887 48546
rect 62799 48482 62817 48534
rect 62869 48482 62887 48534
rect 62799 48470 62887 48482
rect 62799 48418 62817 48470
rect 62869 48418 62887 48470
rect 62799 48406 62887 48418
rect 62799 48354 62817 48406
rect 62869 48354 62887 48406
rect 62799 48342 62887 48354
rect 62799 48290 62817 48342
rect 62869 48290 62887 48342
rect 62799 48278 62887 48290
rect 62799 48226 62817 48278
rect 62869 48226 62887 48278
rect 62799 48208 62887 48226
rect 60462 48065 60499 48117
rect 60551 48065 60590 48117
rect 39449 47789 39756 47795
rect 39449 47673 39465 47789
rect 39581 47743 39756 47789
rect 39581 47673 39597 47743
rect 39449 47667 39597 47673
rect 41359 47633 41446 47659
rect 41359 47581 41376 47633
rect 41428 47581 41446 47633
rect 41359 47569 41446 47581
rect 41359 47517 41376 47569
rect 41428 47517 41446 47569
rect 41359 47505 41446 47517
rect 41359 47453 41376 47505
rect 41428 47453 41446 47505
rect 41359 47427 41446 47453
rect 60462 47437 60590 48065
rect 62727 48113 62811 48119
rect 62727 48061 62743 48113
rect 62795 48061 62811 48113
rect 62727 48055 62811 48061
rect 64101 48117 64185 48123
rect 64101 48065 64117 48117
rect 64169 48065 64185 48117
rect 64101 48059 64185 48065
rect 66460 48117 66588 52556
rect 66460 48065 66499 48117
rect 66551 48065 66588 48117
rect 99940 48167 103294 48196
rect 99940 48115 99959 48167
rect 100011 48115 100023 48167
rect 100075 48115 100087 48167
rect 100139 48115 100151 48167
rect 100203 48115 100215 48167
rect 100267 48115 100279 48167
rect 100331 48115 100343 48167
rect 100395 48115 100407 48167
rect 100459 48115 100471 48167
rect 100523 48115 100535 48167
rect 100587 48115 100599 48167
rect 100651 48115 100663 48167
rect 100715 48115 100727 48167
rect 100779 48115 100791 48167
rect 100843 48115 100855 48167
rect 100907 48115 100919 48167
rect 100971 48115 100983 48167
rect 101035 48115 101047 48167
rect 101099 48115 101111 48167
rect 101163 48115 101175 48167
rect 101227 48115 101239 48167
rect 101291 48115 101303 48167
rect 101355 48115 101367 48167
rect 101419 48115 101431 48167
rect 101483 48115 101495 48167
rect 101547 48115 101559 48167
rect 101611 48115 101623 48167
rect 101675 48115 101687 48167
rect 101739 48115 101751 48167
rect 101803 48115 101815 48167
rect 101867 48115 101879 48167
rect 101931 48115 101943 48167
rect 101995 48115 102007 48167
rect 102059 48115 102071 48167
rect 102123 48115 102135 48167
rect 102187 48115 102199 48167
rect 102251 48115 102263 48167
rect 102315 48115 102327 48167
rect 102379 48115 102391 48167
rect 102443 48115 102455 48167
rect 102507 48115 102519 48167
rect 102571 48115 102583 48167
rect 102635 48115 102647 48167
rect 102699 48115 102711 48167
rect 102763 48115 102775 48167
rect 102827 48115 102839 48167
rect 102891 48115 102903 48167
rect 102955 48115 102967 48167
rect 103019 48115 103031 48167
rect 103083 48115 103095 48167
rect 103147 48115 103159 48167
rect 103211 48115 103223 48167
rect 103275 48115 103294 48167
rect 99940 48087 103294 48115
rect 62818 47417 62882 47683
rect 66460 47445 66588 48065
rect 92236 47882 92320 47888
rect 92236 47830 92252 47882
rect 92304 47830 92320 47882
rect 92236 47824 92320 47830
rect 96430 47715 96524 47736
rect 96430 47663 96451 47715
rect 96503 47663 96524 47715
rect 96430 47651 96524 47663
rect 94903 47631 94996 47633
rect 94903 47579 94923 47631
rect 94975 47579 94996 47631
rect 94903 47567 94996 47579
rect 94903 47515 94923 47567
rect 94975 47515 94996 47567
rect 96430 47599 96451 47651
rect 96503 47599 96524 47651
rect 96430 47587 96524 47599
rect 96430 47535 96451 47587
rect 96503 47535 96524 47587
rect 96430 47515 96524 47535
rect 94903 47514 94996 47515
rect 59644 47350 59944 47414
rect 60954 47353 66096 47417
rect 43101 47236 43111 47288
rect 43163 47236 43385 47288
rect 44695 47275 44785 47299
rect 44695 47223 44714 47275
rect 44766 47223 44785 47275
rect 44695 47211 44785 47223
rect 44695 47159 44714 47211
rect 44766 47159 44785 47211
rect 44695 47147 44785 47159
rect 44695 47095 44714 47147
rect 44766 47095 44785 47147
rect 44695 47083 44785 47095
rect 59644 47085 59708 47350
rect 65871 47349 66047 47353
rect 65871 47297 65901 47349
rect 65953 47297 65965 47349
rect 66017 47297 66047 47349
rect 67162 47348 67360 47412
rect 65871 47268 66047 47297
rect 67296 47085 67360 47348
rect 68390 47317 91029 47445
rect 96540 47325 96776 47453
rect 44695 47031 44714 47083
rect 44766 47031 44785 47083
rect 44695 47019 44785 47031
rect 59634 47079 59718 47085
rect 59634 47027 59650 47079
rect 59702 47027 59718 47079
rect 59634 47021 59718 47027
rect 67286 47079 67370 47085
rect 67286 47027 67302 47079
rect 67354 47027 67370 47079
rect 67286 47021 67370 47027
rect 44695 46967 44714 47019
rect 44766 46967 44785 47019
rect 44695 46955 44785 46967
rect 44695 46903 44714 46955
rect 44766 46903 44785 46955
rect 44695 46879 44785 46903
rect 44629 46795 45631 46798
rect 42176 46741 42186 46793
rect 42238 46741 43480 46793
rect 44634 46792 45631 46795
rect 44634 46740 45499 46792
rect 45551 46740 45563 46792
rect 45615 46740 45631 46792
rect 44634 46734 45631 46740
rect 44693 46623 44781 46646
rect 44693 46571 44711 46623
rect 44763 46571 44781 46623
rect 44693 46559 44781 46571
rect 44693 46507 44711 46559
rect 44763 46507 44781 46559
rect 44693 46495 44781 46507
rect 42680 46429 42690 46481
rect 42742 46429 43354 46481
rect 44693 46443 44711 46495
rect 44763 46443 44781 46495
rect 44693 46421 44781 46443
rect 60489 46123 60553 46128
rect 32844 45687 51163 45724
rect 32844 45635 51014 45687
rect 51066 45635 51078 45687
rect 51130 45635 51163 45687
rect 32844 45596 51163 45635
rect 32810 44825 53755 44864
rect 32810 44773 53599 44825
rect 53651 44773 53663 44825
rect 53715 44773 53755 44825
rect 32810 44736 53755 44773
rect 18916 43074 22243 43087
rect 18916 43022 18953 43074
rect 19005 43022 19017 43074
rect 19069 43022 19081 43074
rect 19133 43022 19145 43074
rect 19197 43022 19209 43074
rect 19261 43022 19273 43074
rect 19325 43022 19337 43074
rect 19389 43022 19401 43074
rect 19453 43022 19465 43074
rect 19517 43022 19529 43074
rect 19581 43022 19593 43074
rect 19645 43022 19657 43074
rect 19709 43022 19721 43074
rect 19773 43022 19785 43074
rect 19837 43022 19849 43074
rect 19901 43022 19913 43074
rect 19965 43022 19977 43074
rect 20029 43022 20041 43074
rect 20093 43022 20105 43074
rect 20157 43022 20169 43074
rect 20221 43022 20233 43074
rect 20285 43022 20297 43074
rect 20349 43022 20361 43074
rect 20413 43022 20425 43074
rect 20477 43022 20489 43074
rect 20541 43022 20553 43074
rect 20605 43022 20617 43074
rect 20669 43022 20681 43074
rect 20733 43022 20745 43074
rect 20797 43022 20809 43074
rect 20861 43022 20873 43074
rect 20925 43022 20937 43074
rect 20989 43022 21001 43074
rect 21053 43022 21065 43074
rect 21117 43022 21129 43074
rect 21181 43022 21193 43074
rect 21245 43022 21257 43074
rect 21309 43022 21321 43074
rect 21373 43022 21385 43074
rect 21437 43022 21449 43074
rect 21501 43022 21513 43074
rect 21565 43022 21577 43074
rect 21629 43022 21641 43074
rect 21693 43022 21705 43074
rect 21757 43022 21769 43074
rect 21821 43022 21833 43074
rect 21885 43022 21897 43074
rect 21949 43022 21961 43074
rect 22013 43022 22025 43074
rect 22077 43022 22089 43074
rect 22141 43022 22153 43074
rect 22205 43022 22243 43074
rect 18916 43009 22243 43022
rect 31632 41918 31717 41944
rect 31632 41866 31648 41918
rect 31700 41866 31717 41918
rect 31632 41854 31717 41866
rect 31632 41802 31648 41854
rect 31700 41802 31717 41854
rect 31632 41790 31717 41802
rect 31632 41738 31648 41790
rect 31700 41738 31717 41790
rect 31632 41726 31717 41738
rect 31632 41674 31648 41726
rect 31700 41674 31717 41726
rect 16488 41624 16744 41652
rect 31632 41649 31717 41674
rect 16488 41444 16526 41624
rect 16706 41604 16744 41624
rect 16706 41598 30419 41604
rect 32810 41601 32938 44736
rect 56640 44125 56724 44131
rect 56640 44073 56656 44125
rect 56708 44073 56724 44125
rect 56640 44061 56724 44073
rect 56640 44009 56656 44061
rect 56708 44009 56724 44061
rect 56640 44003 56724 44009
rect 56650 43015 56714 44003
rect 58768 43426 58906 43432
rect 58768 43374 58784 43426
rect 58836 43374 58906 43426
rect 58768 43362 58906 43374
rect 58768 43310 58784 43362
rect 58836 43310 58906 43362
rect 58768 43304 58906 43310
rect 57317 41788 57401 41794
rect 16706 41482 25970 41598
rect 26086 41482 30419 41598
rect 16706 41476 30419 41482
rect 16706 41444 16744 41476
rect 31737 41473 32938 41601
rect 56273 41547 56337 41757
rect 57317 41736 57333 41788
rect 57385 41736 57401 41788
rect 57317 41730 57401 41736
rect 56263 41541 56347 41547
rect 56263 41489 56279 41541
rect 56331 41489 56347 41541
rect 56263 41483 56347 41489
rect 16488 41416 16744 41444
rect 31634 41398 31726 41426
rect 31634 41346 31654 41398
rect 31706 41346 31726 41398
rect 31634 41334 31726 41346
rect 31634 41282 31654 41334
rect 31706 41282 31726 41334
rect 31634 41270 31726 41282
rect 31634 41218 31654 41270
rect 31706 41218 31726 41270
rect 56649 41243 56713 41712
rect 58778 41243 58906 43304
rect 60455 43362 60583 46123
rect 61481 46007 61491 46059
rect 61543 46007 61553 46059
rect 65312 46007 65322 46059
rect 65374 46007 65384 46059
rect 61491 44967 61543 46007
rect 65322 44967 65374 46007
rect 61481 44915 61491 44967
rect 61543 44915 61553 44967
rect 65312 44915 65322 44967
rect 65374 44915 65384 44967
rect 65322 44905 65374 44915
rect 62478 44125 62562 44131
rect 62478 44073 62494 44125
rect 62546 44073 62562 44125
rect 62478 44061 62562 44073
rect 62478 44009 62494 44061
rect 62546 44009 62562 44061
rect 62478 44003 62562 44009
rect 66457 44125 66585 46127
rect 66457 44073 66494 44125
rect 66546 44073 66585 44125
rect 66457 44061 66585 44073
rect 66457 44009 66494 44061
rect 66546 44009 66585 44061
rect 60455 43310 60495 43362
rect 60547 43310 60583 43362
rect 60145 43122 60229 43128
rect 60145 43070 60161 43122
rect 60213 43070 60229 43122
rect 60455 43094 60583 43310
rect 61941 43180 62298 43195
rect 60145 43064 60229 43070
rect 60977 43009 61453 43073
rect 61941 43064 61965 43180
rect 62273 43064 62298 43180
rect 62488 43120 62552 44003
rect 64478 43426 64562 43432
rect 64478 43374 64494 43426
rect 64546 43374 64562 43426
rect 64478 43362 64562 43374
rect 64478 43310 64494 43362
rect 64546 43310 64562 43362
rect 64478 43304 64562 43310
rect 64169 43122 64253 43128
rect 64488 43125 64552 43304
rect 61941 43049 62298 43064
rect 62976 43013 63385 43077
rect 64169 43070 64185 43122
rect 64237 43070 64253 43122
rect 66065 43122 66149 43128
rect 64169 43064 64253 43070
rect 31634 41191 31726 41218
rect 56639 41237 56723 41243
rect 56639 41185 56655 41237
rect 56707 41185 56723 41237
rect 56639 41173 56723 41185
rect 56639 41121 56655 41173
rect 56707 41121 56723 41173
rect 56639 41115 56723 41121
rect 58768 41237 58906 41243
rect 58768 41185 58784 41237
rect 58836 41185 58906 41237
rect 58768 41173 58906 41185
rect 58768 41121 58784 41173
rect 58836 41121 58906 41173
rect 58768 41115 58906 41121
rect 60487 40888 60551 41791
rect 61389 41311 61453 43009
rect 61379 41305 61463 41311
rect 61379 41253 61395 41305
rect 61447 41253 61463 41305
rect 61379 41247 61463 41253
rect 62487 40888 62551 41790
rect 63321 41311 63385 43013
rect 64971 43011 65438 43075
rect 66065 43070 66081 43122
rect 66133 43070 66149 43122
rect 66457 43096 66585 44009
rect 68390 43434 68518 47317
rect 96419 47220 96525 47222
rect 94903 47214 95009 47216
rect 94903 47162 94930 47214
rect 94982 47162 95009 47214
rect 94903 47150 95009 47162
rect 94903 47098 94930 47150
rect 94982 47098 95009 47150
rect 94903 47086 95009 47098
rect 94903 47034 94930 47086
rect 94982 47034 95009 47086
rect 94903 47022 95009 47034
rect 94903 46970 94930 47022
rect 94982 46970 95009 47022
rect 96419 47168 96446 47220
rect 96498 47168 96525 47220
rect 96419 47156 96525 47168
rect 96419 47104 96446 47156
rect 96498 47104 96525 47156
rect 96419 47092 96525 47104
rect 96419 47040 96446 47092
rect 96498 47040 96525 47092
rect 96419 47028 96525 47040
rect 96419 46976 96446 47028
rect 96498 46976 96525 47028
rect 96419 46974 96525 46976
rect 94903 46968 95009 46970
rect 92184 46632 92194 46812
rect 92374 46632 92384 46812
rect 92844 46747 93125 46752
rect 92844 46695 92862 46747
rect 92914 46695 92926 46747
rect 92978 46695 92990 46747
rect 93042 46695 93054 46747
rect 93106 46695 93125 46747
rect 92844 46690 93125 46695
rect 96648 46699 96776 47325
rect 104640 46728 104896 46756
rect 104640 46699 104678 46728
rect 96648 46571 104678 46699
rect 96430 46389 96524 46410
rect 96430 46337 96451 46389
rect 96503 46337 96524 46389
rect 96430 46325 96524 46337
rect 94910 46295 95000 46302
rect 94910 46243 94929 46295
rect 94981 46243 95000 46295
rect 94910 46231 95000 46243
rect 94910 46179 94929 46231
rect 94981 46179 95000 46231
rect 96430 46273 96451 46325
rect 96503 46273 96524 46325
rect 96430 46261 96524 46273
rect 96430 46209 96451 46261
rect 96503 46209 96524 46261
rect 96430 46189 96524 46209
rect 94910 46173 95000 46179
rect 69467 46018 91009 46146
rect 96650 46129 96778 46571
rect 104640 46548 104678 46571
rect 104858 46548 104896 46728
rect 104640 46520 104896 46548
rect 69467 44133 69595 46018
rect 96558 46001 96778 46129
rect 96425 45854 96531 45856
rect 94898 45834 95003 45845
rect 94898 45782 94924 45834
rect 94976 45782 95003 45834
rect 94898 45770 95003 45782
rect 94898 45718 94924 45770
rect 94976 45718 95003 45770
rect 94898 45706 95003 45718
rect 94898 45654 94924 45706
rect 94976 45654 95003 45706
rect 94898 45643 95003 45654
rect 96425 45802 96452 45854
rect 96504 45802 96531 45854
rect 96425 45790 96531 45802
rect 96425 45738 96452 45790
rect 96504 45738 96531 45790
rect 96425 45726 96531 45738
rect 96425 45674 96452 45726
rect 96504 45674 96531 45726
rect 96425 45662 96531 45674
rect 96425 45610 96452 45662
rect 96504 45610 96531 45662
rect 96425 45608 96531 45610
rect 92236 45601 92320 45607
rect 92236 45549 92252 45601
rect 92304 45549 92320 45601
rect 92236 45543 92320 45549
rect 99938 45171 103292 45200
rect 99938 45119 99957 45171
rect 100009 45119 100021 45171
rect 100073 45119 100085 45171
rect 100137 45119 100149 45171
rect 100201 45119 100213 45171
rect 100265 45119 100277 45171
rect 100329 45119 100341 45171
rect 100393 45119 100405 45171
rect 100457 45119 100469 45171
rect 100521 45119 100533 45171
rect 100585 45119 100597 45171
rect 100649 45119 100661 45171
rect 100713 45119 100725 45171
rect 100777 45119 100789 45171
rect 100841 45119 100853 45171
rect 100905 45119 100917 45171
rect 100969 45119 100981 45171
rect 101033 45119 101045 45171
rect 101097 45119 101109 45171
rect 101161 45119 101173 45171
rect 101225 45119 101237 45171
rect 101289 45119 101301 45171
rect 101353 45119 101365 45171
rect 101417 45119 101429 45171
rect 101481 45119 101493 45171
rect 101545 45119 101557 45171
rect 101609 45119 101621 45171
rect 101673 45119 101685 45171
rect 101737 45119 101749 45171
rect 101801 45119 101813 45171
rect 101865 45119 101877 45171
rect 101929 45119 101941 45171
rect 101993 45119 102005 45171
rect 102057 45119 102069 45171
rect 102121 45119 102133 45171
rect 102185 45119 102197 45171
rect 102249 45119 102261 45171
rect 102313 45119 102325 45171
rect 102377 45119 102389 45171
rect 102441 45119 102453 45171
rect 102505 45119 102517 45171
rect 102569 45119 102581 45171
rect 102633 45119 102645 45171
rect 102697 45119 102709 45171
rect 102761 45119 102773 45171
rect 102825 45119 102837 45171
rect 102889 45119 102901 45171
rect 102953 45119 102965 45171
rect 103017 45119 103029 45171
rect 103081 45119 103093 45171
rect 103145 45119 103157 45171
rect 103209 45119 103221 45171
rect 103273 45119 103292 45171
rect 99938 45091 103292 45119
rect 71772 45043 71856 45049
rect 71772 44991 71788 45043
rect 71840 44991 71856 45043
rect 71772 44985 71856 44991
rect 71782 44519 71846 44985
rect 80754 44232 80838 44238
rect 80754 44180 80770 44232
rect 80822 44180 80838 44232
rect 80754 44174 80838 44180
rect 69457 44127 69605 44133
rect 69457 44011 69473 44127
rect 69589 44011 69605 44127
rect 69457 44005 69605 44011
rect 68379 43428 68527 43434
rect 68379 43312 68395 43428
rect 68511 43312 68527 43428
rect 80773 43398 80857 43404
rect 80773 43346 80789 43398
rect 80841 43346 80857 43398
rect 80773 43340 80857 43346
rect 68379 43306 68527 43312
rect 68390 43283 68518 43306
rect 66065 43064 66149 43070
rect 66971 43074 67400 43080
rect 66971 43022 67332 43074
rect 67384 43022 67400 43074
rect 66971 43016 67400 43022
rect 65374 42740 65438 43011
rect 65364 42734 65448 42740
rect 65364 42682 65380 42734
rect 65432 42682 65448 42734
rect 71761 42710 71795 42765
rect 65364 42676 65448 42682
rect 70658 42704 71822 42710
rect 70658 42652 70674 42704
rect 70726 42652 71822 42704
rect 70658 42646 71822 42652
rect 80742 42444 80826 42450
rect 80742 42392 80758 42444
rect 80810 42392 80826 42444
rect 80742 42386 80826 42392
rect 70971 42005 71055 42069
rect 64487 41381 64551 41797
rect 66490 41381 66554 41796
rect 80773 41568 80857 41574
rect 80773 41516 80789 41568
rect 80841 41516 80857 41568
rect 80773 41510 80857 41516
rect 64477 41375 64561 41381
rect 64477 41323 64493 41375
rect 64545 41323 64561 41375
rect 64477 41311 64561 41323
rect 63311 41305 63395 41311
rect 63311 41253 63327 41305
rect 63379 41253 63395 41305
rect 64477 41259 64493 41311
rect 64545 41259 64561 41311
rect 64477 41253 64561 41259
rect 66480 41375 66564 41381
rect 66480 41323 66496 41375
rect 66548 41323 66564 41375
rect 66480 41311 66564 41323
rect 66480 41259 66496 41311
rect 66548 41259 66564 41311
rect 66480 41253 66564 41259
rect 70969 41375 71053 41381
rect 70969 41323 70985 41375
rect 71037 41323 71053 41375
rect 70969 41311 71053 41323
rect 70969 41259 70985 41311
rect 71037 41259 71053 41311
rect 70969 41253 71053 41259
rect 63311 41247 63395 41253
rect 71774 41099 71858 41105
rect 71774 41047 71790 41099
rect 71842 41047 71858 41099
rect 71774 41041 71858 41047
rect 71784 40916 71848 41041
rect 60477 40882 60561 40888
rect 60477 40830 60493 40882
rect 60545 40830 60561 40882
rect 60477 40818 60561 40830
rect 60477 40766 60493 40818
rect 60545 40766 60561 40818
rect 60477 40760 60561 40766
rect 62477 40882 62561 40888
rect 62477 40830 62493 40882
rect 62545 40830 62561 40882
rect 62477 40818 62561 40830
rect 62477 40766 62493 40818
rect 62545 40766 62561 40818
rect 62477 40760 62561 40766
rect 70361 40882 70445 40888
rect 70361 40830 70377 40882
rect 70429 40830 70445 40882
rect 70361 40818 70445 40830
rect 70361 40766 70377 40818
rect 70429 40766 70445 40818
rect 70361 40760 70445 40766
rect 80156 40678 80821 40742
rect 57335 40454 68243 40468
rect 53168 40310 53232 40319
rect 53158 40304 53242 40310
rect 53158 40252 53174 40304
rect 53226 40252 53242 40304
rect 57335 40274 57355 40454
rect 68223 40274 68243 40454
rect 57335 40260 68243 40274
rect 53158 40246 53242 40252
rect 57112 40182 57291 40211
rect 18910 40079 22252 40097
rect 18910 40027 18923 40079
rect 18975 40027 18987 40079
rect 19039 40027 19051 40079
rect 19103 40027 19115 40079
rect 19167 40027 19179 40079
rect 19231 40027 19243 40079
rect 19295 40027 19307 40079
rect 19359 40027 19371 40079
rect 19423 40027 19435 40079
rect 19487 40027 19499 40079
rect 19551 40027 19563 40079
rect 19615 40027 19627 40079
rect 19679 40027 19691 40079
rect 19743 40027 19755 40079
rect 19807 40027 19819 40079
rect 19871 40027 19883 40079
rect 19935 40027 19947 40079
rect 19999 40027 20011 40079
rect 20063 40027 20075 40079
rect 20127 40027 20139 40079
rect 20191 40027 20203 40079
rect 20255 40027 20267 40079
rect 20319 40027 20331 40079
rect 20383 40027 20395 40079
rect 20447 40027 20459 40079
rect 20511 40027 20523 40079
rect 20575 40027 20587 40079
rect 20639 40027 20651 40079
rect 20703 40027 20715 40079
rect 20767 40027 20779 40079
rect 20831 40027 20843 40079
rect 20895 40027 20907 40079
rect 20959 40027 20971 40079
rect 21023 40027 21035 40079
rect 21087 40027 21099 40079
rect 21151 40027 21163 40079
rect 21215 40027 21227 40079
rect 21279 40027 21291 40079
rect 21343 40027 21355 40079
rect 21407 40027 21419 40079
rect 21471 40027 21483 40079
rect 21535 40027 21547 40079
rect 21599 40027 21611 40079
rect 21663 40027 21675 40079
rect 21727 40027 21739 40079
rect 21791 40027 21803 40079
rect 21855 40027 21867 40079
rect 21919 40027 21931 40079
rect 21983 40027 21995 40079
rect 22047 40027 22059 40079
rect 22111 40027 22123 40079
rect 22175 40027 22187 40079
rect 22239 40027 22252 40079
rect 18910 40009 22252 40027
rect 51307 39730 54045 39731
rect 51298 39724 54045 39730
rect 51298 39672 51314 39724
rect 51366 39672 54045 39724
rect 51298 39667 54045 39672
rect 51298 39666 51382 39667
rect 53981 39565 54045 39667
rect 53167 39105 53180 39157
rect 53232 39105 54123 39157
rect 55270 39106 56416 39158
rect 56468 39106 56478 39158
rect 53940 39002 54043 39020
rect 53940 38950 53965 39002
rect 54017 38950 54043 39002
rect 53940 38938 54043 38950
rect 53940 38886 53965 38938
rect 54017 38886 54043 38938
rect 53940 38874 54043 38886
rect 53940 38822 53965 38874
rect 54017 38822 54043 38874
rect 53940 38810 54043 38822
rect 53940 38758 53965 38810
rect 54017 38758 54043 38810
rect 53940 38741 54043 38758
rect 31567 38445 31660 38468
rect 31567 38393 31587 38445
rect 31639 38393 31660 38445
rect 31567 38381 31660 38393
rect 31567 38329 31587 38381
rect 31639 38329 31660 38381
rect 31567 38317 31660 38329
rect 31567 38265 31587 38317
rect 31639 38265 31660 38317
rect 31567 38253 31660 38265
rect 52182 38453 52272 38468
rect 52182 38401 52201 38453
rect 52253 38401 52272 38453
rect 52182 38389 52272 38401
rect 52182 38337 52201 38389
rect 52253 38337 52272 38389
rect 52182 38325 52272 38337
rect 52182 38273 52201 38325
rect 52253 38273 52272 38325
rect 52182 38258 52272 38273
rect 31567 38201 31587 38253
rect 31639 38201 31660 38253
rect 31567 38179 31660 38201
rect 44020 38157 50807 38163
rect 24093 38118 30339 38124
rect 24093 38002 24109 38118
rect 24225 38002 30339 38118
rect 31733 38095 38954 38127
rect 44020 38105 44036 38157
rect 44088 38105 50556 38157
rect 50608 38105 50807 38157
rect 52278 38109 53180 38161
rect 53232 38109 53242 38161
rect 44020 38099 50807 38105
rect 31502 38089 38954 38095
rect 31502 38037 38877 38089
rect 38929 38037 38954 38089
rect 31502 38031 38954 38037
rect 24093 37996 30339 38002
rect 31733 37999 38954 38031
rect 52167 37996 52271 38020
rect 31566 37919 31658 37947
rect 31566 37867 31586 37919
rect 31638 37867 31658 37919
rect 31566 37855 31658 37867
rect 31566 37803 31586 37855
rect 31638 37803 31658 37855
rect 31566 37791 31658 37803
rect 31566 37739 31586 37791
rect 31638 37739 31658 37791
rect 31566 37712 31658 37739
rect 52167 37944 52193 37996
rect 52245 37944 52271 37996
rect 52167 37932 52271 37944
rect 52167 37880 52193 37932
rect 52245 37880 52271 37932
rect 52167 37868 52271 37880
rect 52167 37816 52193 37868
rect 52245 37816 52271 37868
rect 52167 37804 52271 37816
rect 52167 37752 52193 37804
rect 52245 37752 52271 37804
rect 52167 37728 52271 37752
rect 55276 37137 55379 37155
rect 55276 37085 55301 37137
rect 55353 37085 55379 37137
rect 55276 37073 55379 37085
rect 55276 37021 55301 37073
rect 55353 37021 55379 37073
rect 55276 37009 55379 37021
rect 55276 36957 55301 37009
rect 55353 36957 55379 37009
rect 55276 36945 55379 36957
rect 50540 36908 51317 36914
rect 50540 36856 50556 36908
rect 50608 36856 51249 36908
rect 51301 36856 51317 36908
rect 50540 36850 51317 36856
rect 55276 36893 55301 36945
rect 55353 36893 55379 36945
rect 55276 36881 55379 36893
rect 55276 36829 55301 36881
rect 55353 36829 55379 36881
rect 55276 36817 55379 36829
rect 55276 36765 55301 36817
rect 55353 36765 55379 36817
rect 55276 36748 55379 36765
rect 53180 36657 54067 36658
rect 53170 36605 53180 36657
rect 53232 36605 54067 36657
rect 55369 36607 56815 36659
rect 56867 36607 56877 36659
rect 55309 36425 55670 36431
rect 55309 36373 55602 36425
rect 55654 36373 55670 36425
rect 55309 36367 55670 36373
rect 51233 36235 51317 36241
rect 51233 36183 51249 36235
rect 51301 36183 51317 36235
rect 51233 36177 51317 36183
rect 55296 35551 55391 35552
rect 55296 35542 55411 35551
rect 55296 35490 55342 35542
rect 55394 35490 55411 35542
rect 55296 35478 55411 35490
rect 55296 35426 55342 35478
rect 55394 35426 55411 35478
rect 55296 35414 55411 35426
rect 55296 35362 55342 35414
rect 55394 35362 55411 35414
rect 55296 35350 55411 35362
rect 55296 35298 55342 35350
rect 55394 35298 55411 35350
rect 55296 35286 55411 35298
rect 55296 35234 55342 35286
rect 55394 35234 55411 35286
rect 55296 35222 55411 35234
rect 55296 35170 55342 35222
rect 55394 35170 55411 35222
rect 55296 35162 55411 35170
rect 55296 35161 55391 35162
rect 53669 35004 53679 35056
rect 53731 35004 54062 35056
rect 55370 35005 56815 35057
rect 56867 35005 56877 35057
rect 51239 34913 51249 34965
rect 51301 34913 51311 34965
rect 50922 34843 51167 34855
rect 50922 34791 50954 34843
rect 51006 34791 51018 34843
rect 51070 34791 51082 34843
rect 51134 34791 51167 34843
rect 50922 34780 51167 34791
rect 51377 34842 51703 34860
rect 51377 34790 51418 34842
rect 51470 34790 51482 34842
rect 51534 34790 51546 34842
rect 51598 34790 51610 34842
rect 51662 34790 51703 34842
rect 51377 34773 51703 34790
rect 55291 34799 55670 34805
rect 55291 34747 55602 34799
rect 55654 34747 55670 34799
rect 55291 34741 55670 34747
rect 57112 34690 57143 40182
rect 57259 34690 57291 40182
rect 68323 40185 68503 40206
rect 68323 38469 68355 40185
rect 68471 38469 68503 40185
rect 80156 39518 80220 40678
rect 80770 39804 80854 39810
rect 80770 39752 80786 39804
rect 80838 39752 80854 39804
rect 80770 39746 80854 39752
rect 78012 39512 80857 39518
rect 78012 39460 78028 39512
rect 78080 39460 80857 39512
rect 78012 39454 80857 39460
rect 71774 39244 71858 39250
rect 71774 39192 71790 39244
rect 71842 39192 71858 39244
rect 71774 39186 71858 39192
rect 71784 39152 71848 39186
rect 80793 39114 80857 39454
rect 68323 38454 68397 38469
rect 68431 38454 68503 38469
rect 68323 38448 68503 38454
rect 68362 38442 68467 38448
rect 80770 38013 80854 38019
rect 68362 37976 68467 37987
rect 71769 37981 71853 37987
rect 68341 37968 68488 37976
rect 68341 37020 68356 37968
rect 68472 37020 68488 37968
rect 71769 37929 71785 37981
rect 71837 37929 71853 37981
rect 80770 37961 80786 38013
rect 80838 37961 80854 38013
rect 80770 37955 80854 37961
rect 71769 37923 71853 37929
rect 71774 37544 71858 37550
rect 71774 37492 71790 37544
rect 71842 37492 71858 37544
rect 71774 37486 71858 37492
rect 71784 37349 71848 37486
rect 68341 37012 68488 37020
rect 80769 37022 80853 37028
rect 68362 36999 68467 37012
rect 80769 36970 80785 37022
rect 80837 36970 80853 37022
rect 80769 36964 80853 36970
rect 80775 36206 80859 36212
rect 71786 36196 71870 36202
rect 68327 36122 68502 36151
rect 71786 36144 71802 36196
rect 71854 36144 71870 36196
rect 80775 36154 80791 36206
rect 80843 36154 80859 36206
rect 80775 36148 80859 36154
rect 71786 36138 71870 36144
rect 68327 35366 68356 36122
rect 68472 35366 68502 36122
rect 71776 35692 71860 35698
rect 71776 35640 71792 35692
rect 71844 35640 71860 35692
rect 71776 35634 71860 35640
rect 71786 35542 71850 35634
rect 80773 35535 80857 35541
rect 80773 35483 80789 35535
rect 80841 35483 80857 35535
rect 80773 35477 80857 35483
rect 68327 35359 68397 35366
rect 68431 35359 68502 35366
rect 68327 35338 68502 35359
rect 68362 35333 68467 35338
rect 57112 34662 57291 34690
rect 62756 34424 62808 35052
rect 51239 34423 56416 34424
rect 51239 34371 51249 34423
rect 51301 34372 56416 34423
rect 56468 34372 62808 34424
rect 63578 34494 68312 34558
rect 63578 34460 63666 34494
rect 63700 34460 63738 34494
rect 63772 34460 63810 34494
rect 63844 34460 63882 34494
rect 63916 34460 63954 34494
rect 63988 34460 64026 34494
rect 64060 34460 64098 34494
rect 64132 34460 64170 34494
rect 64204 34460 64242 34494
rect 64276 34460 64314 34494
rect 64348 34460 64386 34494
rect 64420 34460 64458 34494
rect 64492 34460 64530 34494
rect 64564 34460 64602 34494
rect 64636 34460 64674 34494
rect 64708 34460 64746 34494
rect 64780 34460 64818 34494
rect 64852 34460 64890 34494
rect 64924 34460 64962 34494
rect 64996 34460 65034 34494
rect 65068 34460 65106 34494
rect 65140 34460 65178 34494
rect 65212 34460 65250 34494
rect 65284 34460 65322 34494
rect 65356 34460 65394 34494
rect 65428 34460 65466 34494
rect 65500 34460 65538 34494
rect 65572 34460 65610 34494
rect 65644 34460 65682 34494
rect 65716 34460 65754 34494
rect 65788 34460 65826 34494
rect 65860 34460 65898 34494
rect 65932 34460 65970 34494
rect 66004 34460 66042 34494
rect 66076 34460 66114 34494
rect 66148 34460 66186 34494
rect 66220 34460 66258 34494
rect 66292 34460 66330 34494
rect 66364 34460 66402 34494
rect 66436 34460 66474 34494
rect 66508 34460 66546 34494
rect 66580 34460 66618 34494
rect 66652 34460 66690 34494
rect 66724 34460 66762 34494
rect 66796 34460 66834 34494
rect 66868 34460 66906 34494
rect 66940 34460 66978 34494
rect 67012 34460 67050 34494
rect 67084 34460 67122 34494
rect 67156 34460 67194 34494
rect 67228 34460 67266 34494
rect 67300 34460 67338 34494
rect 67372 34460 67410 34494
rect 67444 34460 67482 34494
rect 67516 34460 67554 34494
rect 67588 34460 67626 34494
rect 67660 34460 67698 34494
rect 67732 34460 67770 34494
rect 67804 34460 67842 34494
rect 67876 34460 67914 34494
rect 67948 34460 67986 34494
rect 68020 34460 68058 34494
rect 68092 34460 68130 34494
rect 68164 34460 68312 34494
rect 63578 34379 68312 34460
rect 71775 34399 71859 34405
rect 51301 34371 62808 34372
rect 71775 34347 71791 34399
rect 71843 34347 71859 34399
rect 71775 34341 71859 34347
rect 80775 34396 80859 34402
rect 80775 34344 80791 34396
rect 80843 34344 80859 34396
rect 80775 34338 80859 34344
rect 55325 33939 55409 33952
rect 55325 33887 55341 33939
rect 55393 33887 55409 33939
rect 60842 33933 62361 33967
rect 55325 33875 55409 33887
rect 55325 33823 55341 33875
rect 55393 33823 55409 33875
rect 55325 33811 55409 33823
rect 55325 33759 55341 33811
rect 55393 33759 55409 33811
rect 62327 33778 62361 33933
rect 55325 33747 55409 33759
rect 55325 33695 55341 33747
rect 55393 33695 55409 33747
rect 55325 33683 55409 33695
rect 55325 33631 55341 33683
rect 55393 33631 55409 33683
rect 55325 33619 55409 33631
rect 50917 33600 51175 33614
rect 50917 33548 50956 33600
rect 51008 33548 51020 33600
rect 51072 33548 51084 33600
rect 51136 33548 51175 33600
rect 50917 33535 51175 33548
rect 51376 33600 51705 33617
rect 51376 33548 51386 33600
rect 51438 33548 51450 33600
rect 51502 33548 51514 33600
rect 51566 33548 51578 33600
rect 51630 33548 51642 33600
rect 51694 33548 51705 33600
rect 55325 33567 55341 33619
rect 55393 33567 55409 33619
rect 55325 33554 55409 33567
rect 62325 33691 62361 33778
rect 51376 33531 51705 33548
rect 51239 33422 51249 33474
rect 51301 33422 51311 33474
rect 53170 33407 53180 33459
rect 53232 33407 54054 33459
rect 55368 33405 55945 33457
rect 55997 33405 56007 33457
rect 62325 33440 62359 33691
rect 81628 33440 81712 33446
rect 62307 33439 62380 33440
rect 62307 33387 62317 33439
rect 62369 33387 62380 33439
rect 81628 33388 81644 33440
rect 81696 33388 81712 33440
rect 81628 33382 81712 33388
rect 55315 33141 55670 33147
rect 55315 33089 55602 33141
rect 55654 33089 55670 33141
rect 55315 33083 55670 33089
rect 55326 32338 55414 32352
rect 55326 32286 55344 32338
rect 55396 32286 55414 32338
rect 55326 32274 55414 32286
rect 55326 32222 55344 32274
rect 55396 32222 55414 32274
rect 55326 32210 55414 32222
rect 51231 32190 51315 32196
rect 51231 32138 51247 32190
rect 51299 32138 51315 32190
rect 51231 32132 51315 32138
rect 55326 32158 55344 32210
rect 55396 32158 55414 32210
rect 55326 32146 55414 32158
rect 55326 32094 55344 32146
rect 55396 32094 55414 32146
rect 55326 32082 55414 32094
rect 55326 32030 55344 32082
rect 55396 32030 55414 32082
rect 55326 32018 55414 32030
rect 55326 31966 55344 32018
rect 55396 31966 55414 32018
rect 55326 31952 55414 31966
rect 80292 31866 80365 31867
rect 53669 31805 53679 31857
rect 53731 31805 54065 31857
rect 55368 31805 55945 31857
rect 55997 31805 56007 31857
rect 80292 31814 80302 31866
rect 80354 31814 80365 31866
rect 50522 31613 51315 31617
rect 50519 31611 51315 31613
rect 50519 31607 51247 31611
rect 50519 31555 50535 31607
rect 50587 31559 51247 31607
rect 51299 31559 51315 31611
rect 50587 31555 51315 31559
rect 50519 31553 51315 31555
rect 55298 31602 55670 31608
rect 50519 31549 50603 31553
rect 55298 31550 55602 31602
rect 55654 31550 55670 31602
rect 55298 31544 55670 31550
rect 49870 31235 50353 31265
rect 49870 31055 49893 31235
rect 50329 31197 50353 31235
rect 55586 31260 55670 31280
rect 55586 31208 55602 31260
rect 55654 31208 55670 31260
rect 55586 31197 55670 31208
rect 50329 31196 55670 31197
rect 50329 31144 55602 31196
rect 55654 31144 55670 31196
rect 50329 31132 55670 31144
rect 50329 31088 55602 31132
rect 50329 31055 50353 31088
rect 49870 31025 50353 31055
rect 55586 31080 55602 31088
rect 55654 31080 55670 31132
rect 55586 31068 55670 31080
rect 55586 31016 55602 31068
rect 55654 31016 55670 31068
rect 55586 30996 55670 31016
rect 31563 30682 31658 30691
rect 31563 30630 31584 30682
rect 31636 30630 31658 30682
rect 31563 30618 31658 30630
rect 31563 30566 31584 30618
rect 31636 30566 31658 30618
rect 31563 30554 31658 30566
rect 31563 30502 31584 30554
rect 31636 30502 31658 30554
rect 31563 30490 31658 30502
rect 31563 30438 31584 30490
rect 31636 30438 31658 30490
rect 31563 30430 31658 30438
rect 52167 30687 52268 30717
rect 52167 30635 52191 30687
rect 52243 30635 52268 30687
rect 52167 30623 52268 30635
rect 52167 30571 52191 30623
rect 52243 30571 52268 30623
rect 52167 30559 52268 30571
rect 52167 30507 52191 30559
rect 52243 30507 52268 30559
rect 52167 30495 52268 30507
rect 52167 30443 52191 30495
rect 52243 30443 52268 30495
rect 52167 30414 52268 30443
rect 53980 30467 55670 30473
rect 53980 30415 55602 30467
rect 55654 30415 55670 30467
rect 53980 30409 55670 30415
rect 25954 30353 30350 30359
rect 25954 30237 25970 30353
rect 26086 30237 30350 30353
rect 31720 30325 38945 30358
rect 31491 30319 38945 30325
rect 31491 30267 38849 30319
rect 38901 30267 38945 30319
rect 44009 30329 50833 30335
rect 44009 30277 44025 30329
rect 44077 30277 50535 30329
rect 50587 30277 50833 30329
rect 52288 30280 53679 30332
rect 53731 30280 53741 30332
rect 44009 30271 50833 30277
rect 31491 30261 38945 30267
rect 25954 30231 30350 30237
rect 31720 30230 38945 30261
rect 31562 30195 31657 30196
rect 31562 30143 31583 30195
rect 31635 30143 31657 30195
rect 31562 30131 31657 30143
rect 31562 30079 31583 30131
rect 31635 30079 31657 30131
rect 31562 30067 31657 30079
rect 31562 30015 31583 30067
rect 31635 30015 31657 30067
rect 31562 30003 31657 30015
rect 31562 29951 31583 30003
rect 31635 29951 31657 30003
rect 52177 30168 52263 30185
rect 53980 30183 54044 30409
rect 52177 30116 52194 30168
rect 52246 30116 52263 30168
rect 52177 30104 52263 30116
rect 52177 30052 52194 30104
rect 52246 30052 52263 30104
rect 52177 30040 52263 30052
rect 52177 29988 52194 30040
rect 52246 29988 52263 30040
rect 52177 29972 52263 29988
rect 53669 29693 53679 29745
rect 53731 29693 54124 29745
rect 55262 29693 56416 29745
rect 56468 29693 56478 29745
rect 53891 29580 54025 29599
rect 53891 29528 53916 29580
rect 53968 29528 54025 29580
rect 53891 29516 54025 29528
rect 53891 29464 53916 29516
rect 53968 29464 54025 29516
rect 53891 29452 54025 29464
rect 53891 29400 53916 29452
rect 53968 29400 54025 29452
rect 53891 29388 54025 29400
rect 53891 29336 53916 29388
rect 53968 29336 54025 29388
rect 53891 29318 54025 29336
rect 55945 29151 57993 29152
rect 55935 29099 55945 29151
rect 55997 29099 57993 29151
rect 53657 29063 53741 29069
rect 53657 29011 53673 29063
rect 53725 29011 53741 29063
rect 53657 29005 53741 29011
rect 53667 28995 53731 29005
rect 80302 28938 80355 31814
rect 81638 30334 81702 33382
rect 92108 32299 92192 32305
rect 92108 32247 92124 32299
rect 92176 32247 92192 32299
rect 92108 32241 92192 32247
rect 97184 32139 97285 32143
rect 97184 32087 97208 32139
rect 97260 32087 97285 32139
rect 97184 32075 97285 32087
rect 95659 32045 95749 32060
rect 95659 31993 95678 32045
rect 95730 31993 95749 32045
rect 95659 31981 95749 31993
rect 95659 31929 95678 31981
rect 95730 31929 95749 31981
rect 97184 32023 97208 32075
rect 97260 32023 97285 32075
rect 97184 32011 97285 32023
rect 97184 31959 97208 32011
rect 97260 31959 97285 32011
rect 97184 31955 97285 31959
rect 95659 31914 95749 31929
rect 93385 31895 93636 31903
rect 93385 31843 93420 31895
rect 93472 31843 93484 31895
rect 93536 31843 93548 31895
rect 93600 31843 93636 31895
rect 93385 31836 93636 31843
rect 90830 31667 90914 31673
rect 90830 31615 90846 31667
rect 90898 31615 90914 31667
rect 90830 31609 90914 31615
rect 97171 31594 97272 31598
rect 95652 31581 95753 31585
rect 95652 31529 95676 31581
rect 95728 31529 95753 31581
rect 95652 31517 95753 31529
rect 95652 31465 95676 31517
rect 95728 31465 95753 31517
rect 95652 31453 95753 31465
rect 95652 31401 95676 31453
rect 95728 31401 95753 31453
rect 97171 31542 97195 31594
rect 97247 31542 97272 31594
rect 97171 31530 97272 31542
rect 97171 31478 97195 31530
rect 97247 31478 97272 31530
rect 97171 31466 97272 31478
rect 97171 31414 97195 31466
rect 97247 31414 97272 31466
rect 97171 31410 97272 31414
rect 95652 31397 95753 31401
rect 93446 31354 93635 31359
rect 93446 31302 93482 31354
rect 93534 31302 93546 31354
rect 93598 31302 93635 31354
rect 93446 31297 93635 31302
rect 92112 31239 92196 31245
rect 92112 31187 92128 31239
rect 92180 31187 92196 31239
rect 92112 31181 92196 31187
rect 99686 31235 103027 31254
rect 99686 31183 99698 31235
rect 99750 31183 99762 31235
rect 99814 31183 99826 31235
rect 99878 31183 99890 31235
rect 99942 31183 99954 31235
rect 100006 31183 100018 31235
rect 100070 31183 100082 31235
rect 100134 31183 100146 31235
rect 100198 31183 100210 31235
rect 100262 31183 100274 31235
rect 100326 31183 100338 31235
rect 100390 31183 100402 31235
rect 100454 31183 100466 31235
rect 100518 31183 100530 31235
rect 100582 31183 100594 31235
rect 100646 31183 100658 31235
rect 100710 31183 100722 31235
rect 100774 31183 100786 31235
rect 100838 31183 100850 31235
rect 100902 31183 100914 31235
rect 100966 31183 100978 31235
rect 101030 31183 101042 31235
rect 101094 31183 101106 31235
rect 101158 31183 101170 31235
rect 101222 31183 101234 31235
rect 101286 31183 101298 31235
rect 101350 31183 101362 31235
rect 101414 31183 101426 31235
rect 101478 31183 101490 31235
rect 101542 31183 101554 31235
rect 101606 31183 101618 31235
rect 101670 31183 101682 31235
rect 101734 31183 101746 31235
rect 101798 31183 101810 31235
rect 101862 31183 101874 31235
rect 101926 31183 101938 31235
rect 101990 31183 102002 31235
rect 102054 31183 102066 31235
rect 102118 31183 102130 31235
rect 102182 31183 102194 31235
rect 102246 31183 102258 31235
rect 102310 31183 102322 31235
rect 102374 31183 102386 31235
rect 102438 31183 102450 31235
rect 102502 31183 102514 31235
rect 102566 31183 102578 31235
rect 102630 31183 102642 31235
rect 102694 31183 102706 31235
rect 102758 31183 102770 31235
rect 102822 31183 102834 31235
rect 102886 31183 102898 31235
rect 102950 31183 102962 31235
rect 103014 31183 103027 31235
rect 99686 31165 103027 31183
rect 92111 30970 92195 30976
rect 92111 30918 92127 30970
rect 92179 30918 92195 30970
rect 92111 30912 92195 30918
rect 93436 30806 93541 30817
rect 93436 30754 93462 30806
rect 93514 30754 93541 30806
rect 93436 30743 93541 30754
rect 97176 30803 97277 30807
rect 97176 30751 97200 30803
rect 97252 30751 97277 30803
rect 97176 30739 97277 30751
rect 95655 30724 95753 30729
rect 95655 30672 95678 30724
rect 95730 30672 95753 30724
rect 95655 30660 95753 30672
rect 95655 30608 95678 30660
rect 95730 30608 95753 30660
rect 97176 30687 97200 30739
rect 97252 30687 97277 30739
rect 97176 30675 97277 30687
rect 97176 30623 97200 30675
rect 97252 30623 97277 30675
rect 97176 30619 97277 30623
rect 95655 30604 95753 30608
rect 81628 30328 81712 30334
rect 81628 30276 81644 30328
rect 81696 30276 81712 30328
rect 81628 30270 81712 30276
rect 90818 30328 90902 30334
rect 90818 30276 90834 30328
rect 90886 30276 90902 30328
rect 90818 30270 90902 30276
rect 92851 30265 94171 30287
rect 92851 30213 94087 30265
rect 94139 30213 94171 30265
rect 92851 30191 94171 30213
rect 95647 30250 95748 30254
rect 95647 30198 95671 30250
rect 95723 30198 95748 30250
rect 95647 30186 95748 30198
rect 95647 30134 95671 30186
rect 95723 30134 95748 30186
rect 95647 30122 95748 30134
rect 95647 30070 95671 30122
rect 95723 30070 95748 30122
rect 95647 30066 95748 30070
rect 97176 30247 97277 30251
rect 97176 30195 97200 30247
rect 97252 30195 97277 30247
rect 97176 30183 97277 30195
rect 97176 30131 97200 30183
rect 97252 30131 97277 30183
rect 97176 30119 97277 30131
rect 97176 30067 97200 30119
rect 97252 30067 97277 30119
rect 97176 30063 97277 30067
rect 92111 29901 92195 29907
rect 92111 29849 92127 29901
rect 92179 29849 92195 29901
rect 92111 29843 92195 29849
rect 104557 29794 104813 29822
rect 104557 29766 104595 29794
rect 93054 29723 93253 29729
rect 93054 29671 93095 29723
rect 93147 29671 93159 29723
rect 93211 29671 93253 29723
rect 93054 29666 93253 29671
rect 97450 29638 104595 29766
rect 104557 29614 104595 29638
rect 104775 29614 104813 29794
rect 104557 29586 104813 29614
rect 92108 29578 92192 29584
rect 92108 29526 92124 29578
rect 92176 29526 92192 29578
rect 92108 29520 92192 29526
rect 97193 29423 97294 29427
rect 97193 29371 97217 29423
rect 97269 29371 97294 29423
rect 97193 29359 97294 29371
rect 95658 29334 95752 29344
rect 95658 29282 95679 29334
rect 95731 29282 95752 29334
rect 95658 29270 95752 29282
rect 95658 29218 95679 29270
rect 95731 29218 95752 29270
rect 97193 29307 97217 29359
rect 97269 29307 97294 29359
rect 97193 29295 97294 29307
rect 97193 29243 97217 29295
rect 97269 29243 97294 29295
rect 97193 29239 97294 29243
rect 95658 29209 95752 29218
rect 93598 29175 93838 29184
rect 93598 29123 93628 29175
rect 93680 29123 93692 29175
rect 93744 29123 93756 29175
rect 93808 29123 93838 29175
rect 93598 29114 93838 29123
rect 80292 28937 80365 28938
rect 80292 28885 80302 28937
rect 80354 28885 80365 28937
rect 90826 28937 90899 28938
rect 90826 28885 90836 28937
rect 90888 28885 90899 28937
rect 95646 28897 95747 28901
rect 95646 28845 95670 28897
rect 95722 28845 95747 28897
rect 95646 28833 95747 28845
rect 95646 28781 95670 28833
rect 95722 28781 95747 28833
rect 95646 28769 95747 28781
rect 95646 28717 95670 28769
rect 95722 28717 95747 28769
rect 95646 28713 95747 28717
rect 97176 28875 97277 28879
rect 97176 28823 97200 28875
rect 97252 28823 97277 28875
rect 97176 28811 97277 28823
rect 97176 28759 97200 28811
rect 97252 28759 97277 28811
rect 97176 28747 97277 28759
rect 97176 28695 97200 28747
rect 97252 28695 97277 28747
rect 97176 28691 97277 28695
rect 93448 28632 93613 28635
rect 93448 28580 93472 28632
rect 93524 28580 93536 28632
rect 93588 28580 93613 28632
rect 93448 28577 93613 28580
rect 92119 28508 92203 28514
rect 92119 28456 92135 28508
rect 92187 28456 92203 28508
rect 92119 28450 92203 28456
rect 56841 27811 57961 27812
rect 56805 27759 56815 27811
rect 56867 27759 57961 27811
rect 54973 27320 60455 27438
rect 54973 27202 58755 27320
rect 54973 17437 55209 27202
rect 80516 26428 80589 26429
rect 80516 26376 80526 26428
rect 80578 26376 80589 26428
rect 79673 25118 79746 25119
rect 79673 25066 79683 25118
rect 79735 25066 79746 25118
rect 57324 24314 78478 24413
rect 57153 24229 78478 24314
rect 57153 24205 57446 24229
rect 57406 24113 57446 24205
rect 78170 24205 78478 24229
rect 78170 24113 78211 24205
rect 57406 24089 78211 24113
rect 79683 22005 79736 25066
rect 80526 23382 80579 26376
rect 83095 24738 83170 28419
rect 99683 28236 103063 28255
rect 92108 28203 92192 28209
rect 92108 28151 92124 28203
rect 92176 28151 92192 28203
rect 99683 28184 99715 28236
rect 99767 28184 99779 28236
rect 99831 28184 99843 28236
rect 99895 28184 99907 28236
rect 99959 28184 99971 28236
rect 100023 28184 100035 28236
rect 100087 28184 100099 28236
rect 100151 28184 100163 28236
rect 100215 28184 100227 28236
rect 100279 28184 100291 28236
rect 100343 28184 100355 28236
rect 100407 28184 100419 28236
rect 100471 28184 100483 28236
rect 100535 28184 100547 28236
rect 100599 28184 100611 28236
rect 100663 28184 100675 28236
rect 100727 28184 100739 28236
rect 100791 28184 100803 28236
rect 100855 28184 100867 28236
rect 100919 28184 100931 28236
rect 100983 28184 100995 28236
rect 101047 28184 101059 28236
rect 101111 28184 101123 28236
rect 101175 28184 101187 28236
rect 101239 28184 101251 28236
rect 101303 28184 101315 28236
rect 101367 28184 101379 28236
rect 101431 28184 101443 28236
rect 101495 28184 101507 28236
rect 101559 28184 101571 28236
rect 101623 28184 101635 28236
rect 101687 28184 101699 28236
rect 101751 28184 101763 28236
rect 101815 28184 101827 28236
rect 101879 28184 101891 28236
rect 101943 28184 101955 28236
rect 102007 28184 102019 28236
rect 102071 28184 102083 28236
rect 102135 28184 102147 28236
rect 102199 28184 102211 28236
rect 102263 28184 102275 28236
rect 102327 28184 102339 28236
rect 102391 28184 102403 28236
rect 102455 28184 102467 28236
rect 102519 28184 102531 28236
rect 102583 28184 102595 28236
rect 102647 28184 102659 28236
rect 102711 28184 102723 28236
rect 102775 28184 102787 28236
rect 102839 28184 102851 28236
rect 102903 28184 102915 28236
rect 102967 28184 102979 28236
rect 103031 28184 103063 28236
rect 99683 28166 103063 28184
rect 92108 28145 92192 28151
rect 93393 28089 94172 28111
rect 93393 28037 94088 28089
rect 94140 28037 94172 28089
rect 93393 28015 94172 28037
rect 97183 28044 97284 28048
rect 97183 27992 97207 28044
rect 97259 27992 97284 28044
rect 97183 27980 97284 27992
rect 95656 27937 95755 27956
rect 95656 27885 95679 27937
rect 95731 27885 95755 27937
rect 95656 27873 95755 27885
rect 95656 27821 95679 27873
rect 95731 27821 95755 27873
rect 97183 27928 97207 27980
rect 97259 27928 97284 27980
rect 97183 27916 97284 27928
rect 97183 27864 97207 27916
rect 97259 27864 97284 27916
rect 97183 27860 97284 27864
rect 95656 27803 95755 27821
rect 93443 27543 93590 27553
rect 93443 27491 93458 27543
rect 93510 27491 93522 27543
rect 93574 27491 93590 27543
rect 93443 27481 93590 27491
rect 95649 27497 95750 27501
rect 95649 27445 95673 27497
rect 95725 27445 95750 27497
rect 95649 27433 95750 27445
rect 95649 27381 95673 27433
rect 95725 27381 95750 27433
rect 95649 27369 95750 27381
rect 95649 27317 95673 27369
rect 95725 27317 95750 27369
rect 95649 27313 95750 27317
rect 97173 27491 97274 27495
rect 97173 27439 97197 27491
rect 97249 27439 97274 27491
rect 97173 27427 97274 27439
rect 97173 27375 97197 27427
rect 97249 27375 97274 27427
rect 97173 27363 97274 27375
rect 97173 27311 97197 27363
rect 97249 27311 97274 27363
rect 97173 27307 97274 27311
rect 92115 27138 92199 27144
rect 92115 27086 92131 27138
rect 92183 27086 92199 27138
rect 92115 27080 92199 27086
rect 92108 25359 92192 25365
rect 92108 25307 92124 25359
rect 92176 25307 92192 25359
rect 92108 25301 92192 25307
rect 97184 25199 97285 25203
rect 97184 25147 97208 25199
rect 97260 25147 97285 25199
rect 97184 25135 97285 25147
rect 95659 25105 95749 25120
rect 95659 25053 95678 25105
rect 95730 25053 95749 25105
rect 95659 25041 95749 25053
rect 95659 24989 95678 25041
rect 95730 24989 95749 25041
rect 97184 25083 97208 25135
rect 97260 25083 97285 25135
rect 97184 25071 97285 25083
rect 97184 25019 97208 25071
rect 97260 25019 97285 25071
rect 97184 25015 97285 25019
rect 95659 24974 95749 24989
rect 93385 24955 93636 24963
rect 93385 24903 93420 24955
rect 93472 24903 93484 24955
rect 93536 24903 93548 24955
rect 93600 24903 93636 24955
rect 93385 24896 93636 24903
rect 83085 24726 83180 24738
rect 83085 24674 83106 24726
rect 83158 24674 83180 24726
rect 83085 24663 83180 24674
rect 90814 24733 90909 24738
rect 90814 24726 90914 24733
rect 90814 24674 90835 24726
rect 90887 24674 90914 24726
rect 90814 24669 90914 24674
rect 90814 24663 90909 24669
rect 97171 24654 97272 24658
rect 95652 24641 95753 24645
rect 95652 24589 95676 24641
rect 95728 24589 95753 24641
rect 95652 24577 95753 24589
rect 95652 24525 95676 24577
rect 95728 24525 95753 24577
rect 95652 24513 95753 24525
rect 95652 24461 95676 24513
rect 95728 24461 95753 24513
rect 97171 24602 97195 24654
rect 97247 24602 97272 24654
rect 97171 24590 97272 24602
rect 97171 24538 97195 24590
rect 97247 24538 97272 24590
rect 97171 24526 97272 24538
rect 97171 24474 97195 24526
rect 97247 24474 97272 24526
rect 97171 24470 97272 24474
rect 95652 24457 95753 24461
rect 93446 24414 93635 24419
rect 93446 24362 93482 24414
rect 93534 24362 93546 24414
rect 93598 24362 93635 24414
rect 93446 24357 93635 24362
rect 92112 24299 92196 24305
rect 92112 24247 92128 24299
rect 92180 24247 92196 24299
rect 92112 24241 92196 24247
rect 99683 24302 103034 24331
rect 99683 24250 99700 24302
rect 99752 24250 99764 24302
rect 99816 24250 99828 24302
rect 99880 24250 99892 24302
rect 99944 24250 99956 24302
rect 100008 24250 100020 24302
rect 100072 24250 100084 24302
rect 100136 24250 100148 24302
rect 100200 24250 100212 24302
rect 100264 24250 100276 24302
rect 100328 24250 100340 24302
rect 100392 24250 100404 24302
rect 100456 24250 100468 24302
rect 100520 24250 100532 24302
rect 100584 24250 100596 24302
rect 100648 24250 100660 24302
rect 100712 24250 100724 24302
rect 100776 24250 100788 24302
rect 100840 24250 100852 24302
rect 100904 24250 100916 24302
rect 100968 24250 100980 24302
rect 101032 24250 101044 24302
rect 101096 24250 101108 24302
rect 101160 24250 101172 24302
rect 101224 24250 101236 24302
rect 101288 24250 101300 24302
rect 101352 24250 101364 24302
rect 101416 24250 101428 24302
rect 101480 24250 101492 24302
rect 101544 24250 101556 24302
rect 101608 24250 101620 24302
rect 101672 24250 101684 24302
rect 101736 24250 101748 24302
rect 101800 24250 101812 24302
rect 101864 24250 101876 24302
rect 101928 24250 101940 24302
rect 101992 24250 102004 24302
rect 102056 24250 102068 24302
rect 102120 24250 102132 24302
rect 102184 24250 102196 24302
rect 102248 24250 102260 24302
rect 102312 24250 102324 24302
rect 102376 24250 102388 24302
rect 102440 24250 102452 24302
rect 102504 24250 102516 24302
rect 102568 24250 102580 24302
rect 102632 24250 102644 24302
rect 102696 24250 102708 24302
rect 102760 24250 102772 24302
rect 102824 24250 102836 24302
rect 102888 24250 102900 24302
rect 102952 24250 102964 24302
rect 103016 24250 103034 24302
rect 99683 24221 103034 24250
rect 92111 24030 92195 24036
rect 92111 23978 92127 24030
rect 92179 23978 92195 24030
rect 92111 23972 92195 23978
rect 93436 23866 93541 23877
rect 93436 23814 93462 23866
rect 93514 23814 93541 23866
rect 93436 23803 93541 23814
rect 97176 23863 97277 23867
rect 97176 23811 97200 23863
rect 97252 23811 97277 23863
rect 97176 23799 97277 23811
rect 95655 23784 95753 23789
rect 95655 23732 95678 23784
rect 95730 23732 95753 23784
rect 95655 23720 95753 23732
rect 95655 23668 95678 23720
rect 95730 23668 95753 23720
rect 97176 23747 97200 23799
rect 97252 23747 97277 23799
rect 97176 23735 97277 23747
rect 97176 23683 97200 23735
rect 97252 23683 97277 23735
rect 97176 23679 97277 23683
rect 95655 23664 95753 23668
rect 90818 23387 90902 23394
rect 80516 23381 80589 23382
rect 80516 23329 80526 23381
rect 80578 23329 80589 23381
rect 90818 23335 90835 23387
rect 90887 23335 90902 23387
rect 90818 23330 90902 23335
rect 90825 23329 90898 23330
rect 92851 23325 94171 23347
rect 92851 23273 94087 23325
rect 94139 23273 94171 23325
rect 92851 23251 94171 23273
rect 95647 23310 95748 23314
rect 95647 23258 95671 23310
rect 95723 23258 95748 23310
rect 95647 23246 95748 23258
rect 95647 23194 95671 23246
rect 95723 23194 95748 23246
rect 95647 23182 95748 23194
rect 95647 23130 95671 23182
rect 95723 23130 95748 23182
rect 95647 23126 95748 23130
rect 97176 23307 97277 23311
rect 97176 23255 97200 23307
rect 97252 23255 97277 23307
rect 97176 23243 97277 23255
rect 97176 23191 97200 23243
rect 97252 23191 97277 23243
rect 97176 23179 97277 23191
rect 97176 23127 97200 23179
rect 97252 23127 97277 23179
rect 97176 23123 97277 23127
rect 92111 22961 92195 22967
rect 92111 22909 92127 22961
rect 92179 22909 92195 22961
rect 92111 22903 92195 22909
rect 104573 22854 104829 22882
rect 104573 22826 104611 22854
rect 93054 22783 93253 22789
rect 93054 22731 93095 22783
rect 93147 22731 93159 22783
rect 93211 22731 93253 22783
rect 93054 22726 93253 22731
rect 97450 22698 104611 22826
rect 104573 22674 104611 22698
rect 104791 22674 104829 22854
rect 104573 22646 104829 22674
rect 92108 22638 92192 22644
rect 92108 22586 92124 22638
rect 92176 22586 92192 22638
rect 92108 22580 92192 22586
rect 97193 22483 97294 22487
rect 97193 22431 97217 22483
rect 97269 22431 97294 22483
rect 97193 22419 97294 22431
rect 95658 22394 95752 22404
rect 95658 22342 95679 22394
rect 95731 22342 95752 22394
rect 95658 22330 95752 22342
rect 95658 22278 95679 22330
rect 95731 22278 95752 22330
rect 97193 22367 97217 22419
rect 97269 22367 97294 22419
rect 97193 22355 97294 22367
rect 97193 22303 97217 22355
rect 97269 22303 97294 22355
rect 97193 22299 97294 22303
rect 95658 22269 95752 22278
rect 93598 22235 93838 22244
rect 93598 22183 93628 22235
rect 93680 22183 93692 22235
rect 93744 22183 93756 22235
rect 93808 22183 93838 22235
rect 93598 22174 93838 22183
rect 79673 22004 79747 22005
rect 79673 21952 79684 22004
rect 79736 21952 79747 22004
rect 90830 22001 90910 22005
rect 79683 21949 79736 21952
rect 90830 21949 90844 22001
rect 90896 21949 90910 22001
rect 90830 21945 90910 21949
rect 95646 21957 95747 21961
rect 95646 21905 95670 21957
rect 95722 21905 95747 21957
rect 95646 21893 95747 21905
rect 95646 21841 95670 21893
rect 95722 21841 95747 21893
rect 95646 21829 95747 21841
rect 95646 21777 95670 21829
rect 95722 21777 95747 21829
rect 95646 21773 95747 21777
rect 97176 21935 97277 21939
rect 97176 21883 97200 21935
rect 97252 21883 97277 21935
rect 97176 21871 97277 21883
rect 97176 21819 97200 21871
rect 97252 21819 97277 21871
rect 97176 21807 97277 21819
rect 97176 21755 97200 21807
rect 97252 21755 97277 21807
rect 97176 21751 97277 21755
rect 93448 21692 93613 21695
rect 93448 21640 93472 21692
rect 93524 21640 93536 21692
rect 93588 21640 93613 21692
rect 93448 21637 93613 21640
rect 92119 21568 92203 21574
rect 92119 21516 92135 21568
rect 92187 21516 92203 21568
rect 92119 21510 92203 21516
rect 99671 21296 103037 21314
rect 92108 21263 92192 21269
rect 92108 21211 92124 21263
rect 92176 21211 92192 21263
rect 99671 21244 99696 21296
rect 99748 21244 99760 21296
rect 99812 21244 99824 21296
rect 99876 21244 99888 21296
rect 99940 21244 99952 21296
rect 100004 21244 100016 21296
rect 100068 21244 100080 21296
rect 100132 21244 100144 21296
rect 100196 21244 100208 21296
rect 100260 21244 100272 21296
rect 100324 21244 100336 21296
rect 100388 21244 100400 21296
rect 100452 21244 100464 21296
rect 100516 21244 100528 21296
rect 100580 21244 100592 21296
rect 100644 21244 100656 21296
rect 100708 21244 100720 21296
rect 100772 21244 100784 21296
rect 100836 21244 100848 21296
rect 100900 21244 100912 21296
rect 100964 21244 100976 21296
rect 101028 21244 101040 21296
rect 101092 21244 101104 21296
rect 101156 21244 101168 21296
rect 101220 21244 101232 21296
rect 101284 21244 101296 21296
rect 101348 21244 101360 21296
rect 101412 21244 101424 21296
rect 101476 21244 101488 21296
rect 101540 21244 101552 21296
rect 101604 21244 101616 21296
rect 101668 21244 101680 21296
rect 101732 21244 101744 21296
rect 101796 21244 101808 21296
rect 101860 21244 101872 21296
rect 101924 21244 101936 21296
rect 101988 21244 102000 21296
rect 102052 21244 102064 21296
rect 102116 21244 102128 21296
rect 102180 21244 102192 21296
rect 102244 21244 102256 21296
rect 102308 21244 102320 21296
rect 102372 21244 102384 21296
rect 102436 21244 102448 21296
rect 102500 21244 102512 21296
rect 102564 21244 102576 21296
rect 102628 21244 102640 21296
rect 102692 21244 102704 21296
rect 102756 21244 102768 21296
rect 102820 21244 102832 21296
rect 102884 21244 102896 21296
rect 102948 21244 102960 21296
rect 103012 21244 103037 21296
rect 99671 21226 103037 21244
rect 92108 21205 92192 21211
rect 93393 21149 94172 21171
rect 93393 21097 94088 21149
rect 94140 21097 94172 21149
rect 93393 21075 94172 21097
rect 97183 21104 97284 21108
rect 97183 21052 97207 21104
rect 97259 21052 97284 21104
rect 97183 21040 97284 21052
rect 95656 20997 95755 21016
rect 95656 20945 95679 20997
rect 95731 20945 95755 20997
rect 95656 20933 95755 20945
rect 95656 20881 95679 20933
rect 95731 20881 95755 20933
rect 97183 20988 97207 21040
rect 97259 20988 97284 21040
rect 97183 20976 97284 20988
rect 97183 20924 97207 20976
rect 97259 20924 97284 20976
rect 97183 20920 97284 20924
rect 95656 20863 95755 20881
rect 93443 20603 93590 20613
rect 93443 20551 93458 20603
rect 93510 20551 93522 20603
rect 93574 20551 93590 20603
rect 93443 20541 93590 20551
rect 95649 20557 95750 20561
rect 95649 20505 95673 20557
rect 95725 20505 95750 20557
rect 95649 20493 95750 20505
rect 95649 20441 95673 20493
rect 95725 20441 95750 20493
rect 95649 20429 95750 20441
rect 95649 20377 95673 20429
rect 95725 20377 95750 20429
rect 95649 20373 95750 20377
rect 97173 20551 97274 20555
rect 97173 20499 97197 20551
rect 97249 20499 97274 20551
rect 97173 20487 97274 20499
rect 97173 20435 97197 20487
rect 97249 20435 97274 20487
rect 97173 20423 97274 20435
rect 97173 20371 97197 20423
rect 97249 20371 97274 20423
rect 97173 20367 97274 20371
rect 92115 20198 92199 20204
rect 92115 20146 92131 20198
rect 92183 20146 92199 20198
rect 92115 20140 92199 20146
rect 54973 17223 55101 17437
rect 53489 17172 53601 17200
rect 53489 17120 53519 17172
rect 53571 17120 53601 17172
rect 53489 17108 53601 17120
rect 53489 17056 53519 17108
rect 53571 17056 53601 17108
rect 53489 17044 53601 17056
rect 53489 16992 53519 17044
rect 53571 16992 53601 17044
rect 53489 16980 53601 16992
rect 53489 16928 53519 16980
rect 53571 16928 53601 16980
rect 53489 16916 53601 16928
rect 53489 16864 53519 16916
rect 53571 16864 53601 16916
rect 53489 16852 53601 16864
rect 53489 16800 53519 16852
rect 53571 16800 53601 16852
rect 53489 16788 53601 16800
rect 53489 16736 53519 16788
rect 53571 16736 53601 16788
rect 53489 16724 53601 16736
rect 53489 16672 53519 16724
rect 53571 16672 53601 16724
rect 53489 16660 53601 16672
rect 53489 16608 53519 16660
rect 53571 16608 53601 16660
rect 53489 16596 53601 16608
rect 53489 16544 53519 16596
rect 53571 16544 53601 16596
rect 53489 16532 53601 16544
rect 53489 16480 53519 16532
rect 53571 16480 53601 16532
rect 53489 16468 53601 16480
rect 53489 16416 53519 16468
rect 53571 16416 53601 16468
rect 53489 16404 53601 16416
rect 53489 16352 53519 16404
rect 53571 16352 53601 16404
rect 53489 16340 53601 16352
rect 53489 16288 53519 16340
rect 53571 16288 53601 16340
rect 53489 16276 53601 16288
rect 53489 16224 53519 16276
rect 53571 16224 53601 16276
rect 53489 16212 53601 16224
rect 53489 16160 53519 16212
rect 53571 16160 53601 16212
rect 53489 16148 53601 16160
rect 53489 16096 53519 16148
rect 53571 16096 53601 16148
rect 53489 16084 53601 16096
rect 53489 16032 53519 16084
rect 53571 16032 53601 16084
rect 53489 16020 53601 16032
rect 53489 15968 53519 16020
rect 53571 15968 53601 16020
rect 53489 15956 53601 15968
rect 53489 15904 53519 15956
rect 53571 15904 53601 15956
rect 53489 15892 53601 15904
rect 53489 15840 53519 15892
rect 53571 15840 53601 15892
rect 53489 15828 53601 15840
rect 53489 15776 53519 15828
rect 53571 15776 53601 15828
rect 53489 15764 53601 15776
rect 53489 15712 53519 15764
rect 53571 15712 53601 15764
rect 53489 15700 53601 15712
rect 53489 15648 53519 15700
rect 53571 15648 53601 15700
rect 53489 15636 53601 15648
rect 53489 15584 53519 15636
rect 53571 15584 53601 15636
rect 53489 15572 53601 15584
rect 53489 15520 53519 15572
rect 53571 15520 53601 15572
rect 53489 15508 53601 15520
rect 53489 15456 53519 15508
rect 53571 15456 53601 15508
rect 53489 15444 53601 15456
rect 53489 15392 53519 15444
rect 53571 15392 53601 15444
rect 53489 15380 53601 15392
rect 53489 15328 53519 15380
rect 53571 15328 53601 15380
rect 53489 15316 53601 15328
rect 53489 15264 53519 15316
rect 53571 15264 53601 15316
rect 53489 15252 53601 15264
rect 53489 15200 53519 15252
rect 53571 15200 53601 15252
rect 53489 15188 53601 15200
rect 53489 15136 53519 15188
rect 53571 15136 53601 15188
rect 53489 15124 53601 15136
rect 53489 15072 53519 15124
rect 53571 15072 53601 15124
rect 53489 15060 53601 15072
rect 53489 15008 53519 15060
rect 53571 15008 53601 15060
rect 53489 14996 53601 15008
rect 53489 14944 53519 14996
rect 53571 14944 53601 14996
rect 53489 14932 53601 14944
rect 53489 14880 53519 14932
rect 53571 14880 53601 14932
rect 53489 14868 53601 14880
rect 53489 14816 53519 14868
rect 53571 14816 53601 14868
rect 53489 14804 53601 14816
rect 53489 14752 53519 14804
rect 53571 14752 53601 14804
rect 53489 14740 53601 14752
rect 53489 14688 53519 14740
rect 53571 14688 53601 14740
rect 53489 14676 53601 14688
rect 53489 14624 53519 14676
rect 53571 14624 53601 14676
rect 53489 14612 53601 14624
rect 53489 14560 53519 14612
rect 53571 14560 53601 14612
rect 53489 14548 53601 14560
rect 53489 14496 53519 14548
rect 53571 14496 53601 14548
rect 53489 14484 53601 14496
rect 53489 14432 53519 14484
rect 53571 14432 53601 14484
rect 53489 14420 53601 14432
rect 53489 14368 53519 14420
rect 53571 14368 53601 14420
rect 53489 14356 53601 14368
rect 53489 14304 53519 14356
rect 53571 14304 53601 14356
rect 53489 14292 53601 14304
rect 53489 14240 53519 14292
rect 53571 14240 53601 14292
rect 53489 14228 53601 14240
rect 53489 14176 53519 14228
rect 53571 14176 53601 14228
rect 53489 14164 53601 14176
rect 53489 14112 53519 14164
rect 53571 14112 53601 14164
rect 53489 14100 53601 14112
rect 53489 14048 53519 14100
rect 53571 14048 53601 14100
rect 53489 14036 53601 14048
rect 53489 13984 53519 14036
rect 53571 13984 53601 14036
rect 53489 13972 53601 13984
rect 53489 13920 53519 13972
rect 53571 13920 53601 13972
rect 53489 13892 53601 13920
rect 54973 13657 55091 17223
rect 56484 17165 56618 17197
rect 56484 17113 56525 17165
rect 56577 17113 56618 17165
rect 56484 17101 56618 17113
rect 56484 17049 56525 17101
rect 56577 17049 56618 17101
rect 56484 17037 56618 17049
rect 56484 16985 56525 17037
rect 56577 16985 56618 17037
rect 56484 16973 56618 16985
rect 56484 16921 56525 16973
rect 56577 16921 56618 16973
rect 56484 16909 56618 16921
rect 56484 16857 56525 16909
rect 56577 16857 56618 16909
rect 56484 16845 56618 16857
rect 56484 16793 56525 16845
rect 56577 16793 56618 16845
rect 56484 16781 56618 16793
rect 56484 16729 56525 16781
rect 56577 16729 56618 16781
rect 56484 16717 56618 16729
rect 56484 16665 56525 16717
rect 56577 16665 56618 16717
rect 56484 16653 56618 16665
rect 56484 16601 56525 16653
rect 56577 16601 56618 16653
rect 56484 16589 56618 16601
rect 56484 16537 56525 16589
rect 56577 16537 56618 16589
rect 56484 16525 56618 16537
rect 56484 16473 56525 16525
rect 56577 16473 56618 16525
rect 56484 16461 56618 16473
rect 56484 16409 56525 16461
rect 56577 16409 56618 16461
rect 56484 16397 56618 16409
rect 56484 16345 56525 16397
rect 56577 16345 56618 16397
rect 56484 16333 56618 16345
rect 56484 16281 56525 16333
rect 56577 16281 56618 16333
rect 56484 16269 56618 16281
rect 56484 16217 56525 16269
rect 56577 16217 56618 16269
rect 56484 16205 56618 16217
rect 56484 16153 56525 16205
rect 56577 16153 56618 16205
rect 56484 16141 56618 16153
rect 56484 16089 56525 16141
rect 56577 16089 56618 16141
rect 56484 16077 56618 16089
rect 56484 16025 56525 16077
rect 56577 16025 56618 16077
rect 56484 16013 56618 16025
rect 56484 15961 56525 16013
rect 56577 15961 56618 16013
rect 56484 15949 56618 15961
rect 56484 15897 56525 15949
rect 56577 15897 56618 15949
rect 56484 15885 56618 15897
rect 56484 15833 56525 15885
rect 56577 15833 56618 15885
rect 56484 15821 56618 15833
rect 56484 15769 56525 15821
rect 56577 15769 56618 15821
rect 56484 15757 56618 15769
rect 56484 15705 56525 15757
rect 56577 15705 56618 15757
rect 56484 15693 56618 15705
rect 56484 15641 56525 15693
rect 56577 15641 56618 15693
rect 56484 15629 56618 15641
rect 56484 15577 56525 15629
rect 56577 15577 56618 15629
rect 56484 15565 56618 15577
rect 56484 15513 56525 15565
rect 56577 15513 56618 15565
rect 56484 15501 56618 15513
rect 56484 15449 56525 15501
rect 56577 15449 56618 15501
rect 56484 15437 56618 15449
rect 56484 15385 56525 15437
rect 56577 15385 56618 15437
rect 56484 15373 56618 15385
rect 56484 15321 56525 15373
rect 56577 15321 56618 15373
rect 56484 15309 56618 15321
rect 56484 15257 56525 15309
rect 56577 15257 56618 15309
rect 56484 15245 56618 15257
rect 56484 15193 56525 15245
rect 56577 15193 56618 15245
rect 56484 15181 56618 15193
rect 56484 15129 56525 15181
rect 56577 15129 56618 15181
rect 56484 15117 56618 15129
rect 56484 15065 56525 15117
rect 56577 15065 56618 15117
rect 56484 15053 56618 15065
rect 56484 15001 56525 15053
rect 56577 15001 56618 15053
rect 56484 14989 56618 15001
rect 56484 14937 56525 14989
rect 56577 14937 56618 14989
rect 56484 14925 56618 14937
rect 56484 14873 56525 14925
rect 56577 14873 56618 14925
rect 56484 14861 56618 14873
rect 56484 14809 56525 14861
rect 56577 14809 56618 14861
rect 56484 14797 56618 14809
rect 56484 14745 56525 14797
rect 56577 14745 56618 14797
rect 56484 14733 56618 14745
rect 56484 14681 56525 14733
rect 56577 14681 56618 14733
rect 56484 14669 56618 14681
rect 56484 14617 56525 14669
rect 56577 14617 56618 14669
rect 56484 14605 56618 14617
rect 56484 14553 56525 14605
rect 56577 14553 56618 14605
rect 56484 14541 56618 14553
rect 56484 14489 56525 14541
rect 56577 14489 56618 14541
rect 56484 14477 56618 14489
rect 56484 14425 56525 14477
rect 56577 14425 56618 14477
rect 56484 14413 56618 14425
rect 56484 14361 56525 14413
rect 56577 14361 56618 14413
rect 56484 14349 56618 14361
rect 56484 14297 56525 14349
rect 56577 14297 56618 14349
rect 56484 14285 56618 14297
rect 56484 14233 56525 14285
rect 56577 14233 56618 14285
rect 56484 14221 56618 14233
rect 56484 14169 56525 14221
rect 56577 14169 56618 14221
rect 56484 14157 56618 14169
rect 56484 14105 56525 14157
rect 56577 14105 56618 14157
rect 56484 14093 56618 14105
rect 56484 14041 56525 14093
rect 56577 14041 56618 14093
rect 56484 14029 56618 14041
rect 56484 13977 56525 14029
rect 56577 13977 56618 14029
rect 56484 13965 56618 13977
rect 56484 13913 56525 13965
rect 56577 13913 56618 13965
rect 56484 13882 56618 13913
rect 54915 11940 55151 13657
rect 54905 11912 55161 11940
rect 54905 11732 54943 11912
rect 55123 11732 55161 11912
rect 54905 11704 55161 11732
<< via1 >>
rect 41712 101954 41892 102134
rect 40269 100688 40321 100740
rect 40269 100624 40321 100676
rect 40269 100560 40321 100612
rect 40269 100496 40321 100548
rect 40269 100432 40321 100484
rect 40269 100368 40321 100420
rect 40269 100304 40321 100356
rect 40269 100240 40321 100292
rect 40269 100176 40321 100228
rect 40269 100112 40321 100164
rect 40269 100048 40321 100100
rect 40269 99984 40321 100036
rect 40269 99920 40321 99972
rect 40269 99856 40321 99908
rect 40269 99792 40321 99844
rect 40269 99728 40321 99780
rect 40269 99664 40321 99716
rect 40269 99600 40321 99652
rect 40269 99536 40321 99588
rect 40269 99472 40321 99524
rect 40269 99408 40321 99460
rect 40269 99344 40321 99396
rect 40269 99280 40321 99332
rect 69728 101925 69908 102105
rect 81778 101926 81958 102106
rect 43270 100694 43322 100746
rect 43270 100630 43322 100682
rect 43270 100566 43322 100618
rect 43270 100502 43322 100554
rect 43270 100438 43322 100490
rect 43270 100374 43322 100426
rect 43270 100310 43322 100362
rect 43270 100246 43322 100298
rect 43270 100182 43322 100234
rect 43270 100118 43322 100170
rect 43270 100054 43322 100106
rect 43270 99990 43322 100042
rect 43270 99926 43322 99978
rect 43270 99862 43322 99914
rect 43270 99798 43322 99850
rect 43270 99734 43322 99786
rect 43270 99670 43322 99722
rect 43270 99606 43322 99658
rect 43270 99542 43322 99594
rect 43270 99478 43322 99530
rect 43270 99414 43322 99466
rect 43270 99350 43322 99402
rect 43270 99286 43322 99338
rect 40269 99216 40321 99268
rect 40269 99152 40321 99204
rect 40269 99088 40321 99140
rect 40269 99024 40321 99076
rect 40269 98960 40321 99012
rect 40269 98896 40321 98948
rect 40269 98832 40321 98884
rect 43270 99222 43322 99274
rect 43270 99158 43322 99210
rect 43270 99094 43322 99146
rect 43270 99030 43322 99082
rect 43270 98966 43322 99018
rect 43270 98902 43322 98954
rect 43270 98838 43322 98890
rect 40269 98768 40321 98820
rect 40269 98704 40321 98756
rect 40269 98640 40321 98692
rect 40269 98576 40321 98628
rect 40269 98512 40321 98564
rect 40269 98448 40321 98500
rect 40269 98384 40321 98436
rect 40269 98320 40321 98372
rect 40269 98256 40321 98308
rect 40269 98192 40321 98244
rect 40269 98128 40321 98180
rect 40269 98064 40321 98116
rect 40269 98000 40321 98052
rect 40269 97936 40321 97988
rect 40269 97872 40321 97924
rect 40269 97808 40321 97860
rect 40269 97744 40321 97796
rect 40269 97680 40321 97732
rect 40269 97616 40321 97668
rect 40269 97552 40321 97604
rect 40269 97488 40321 97540
rect 40269 97424 40321 97476
rect 43270 98774 43322 98826
rect 43270 98710 43322 98762
rect 43270 98646 43322 98698
rect 43270 98582 43322 98634
rect 43270 98518 43322 98570
rect 43270 98454 43322 98506
rect 43270 98390 43322 98442
rect 43270 98326 43322 98378
rect 43270 98262 43322 98314
rect 43270 98198 43322 98250
rect 43270 98134 43322 98186
rect 43270 98070 43322 98122
rect 43270 98006 43322 98058
rect 43270 97942 43322 97994
rect 43270 97878 43322 97930
rect 43270 97814 43322 97866
rect 43270 97750 43322 97802
rect 43270 97686 43322 97738
rect 43270 97622 43322 97674
rect 43270 97558 43322 97610
rect 43270 97494 43322 97546
rect 43270 97430 43322 97482
rect 68243 100686 68359 100742
rect 68243 100652 68283 100686
rect 68283 100652 68317 100686
rect 68317 100652 68359 100686
rect 68243 100614 68359 100652
rect 68243 100580 68283 100614
rect 68283 100580 68317 100614
rect 68317 100580 68359 100614
rect 68243 100542 68359 100580
rect 68243 100508 68283 100542
rect 68283 100508 68317 100542
rect 68317 100508 68359 100542
rect 68243 100470 68359 100508
rect 68243 100436 68283 100470
rect 68283 100436 68317 100470
rect 68317 100436 68359 100470
rect 68243 100398 68359 100436
rect 68243 100364 68283 100398
rect 68283 100364 68317 100398
rect 68317 100364 68359 100398
rect 68243 100326 68359 100364
rect 68243 100292 68283 100326
rect 68283 100292 68317 100326
rect 68317 100292 68359 100326
rect 68243 100254 68359 100292
rect 68243 100220 68283 100254
rect 68283 100220 68317 100254
rect 68317 100220 68359 100254
rect 68243 100182 68359 100220
rect 68243 100148 68283 100182
rect 68283 100148 68317 100182
rect 68317 100148 68359 100182
rect 68243 100110 68359 100148
rect 68243 100076 68283 100110
rect 68283 100076 68317 100110
rect 68317 100076 68359 100110
rect 68243 100038 68359 100076
rect 68243 100004 68283 100038
rect 68283 100004 68317 100038
rect 68317 100004 68359 100038
rect 68243 99966 68359 100004
rect 68243 99932 68283 99966
rect 68283 99932 68317 99966
rect 68317 99932 68359 99966
rect 68243 99894 68359 99932
rect 68243 99860 68283 99894
rect 68283 99860 68317 99894
rect 68317 99860 68359 99894
rect 68243 99822 68359 99860
rect 68243 99788 68283 99822
rect 68283 99788 68317 99822
rect 68317 99788 68359 99822
rect 68243 99750 68359 99788
rect 68243 99716 68283 99750
rect 68283 99716 68317 99750
rect 68317 99716 68359 99750
rect 68243 99678 68359 99716
rect 68243 99644 68283 99678
rect 68283 99644 68317 99678
rect 68317 99644 68359 99678
rect 68243 99606 68359 99644
rect 68243 99572 68283 99606
rect 68283 99572 68317 99606
rect 68317 99572 68359 99606
rect 68243 99534 68359 99572
rect 68243 99500 68283 99534
rect 68283 99500 68317 99534
rect 68317 99500 68359 99534
rect 68243 99462 68359 99500
rect 68243 99428 68283 99462
rect 68283 99428 68317 99462
rect 68317 99428 68359 99462
rect 68243 99390 68359 99428
rect 68243 99356 68283 99390
rect 68283 99356 68317 99390
rect 68317 99356 68359 99390
rect 68243 99318 68359 99356
rect 68243 99284 68283 99318
rect 68283 99284 68317 99318
rect 68317 99284 68359 99318
rect 68243 99246 68359 99284
rect 68243 99212 68283 99246
rect 68283 99212 68317 99246
rect 68317 99212 68359 99246
rect 68243 99174 68359 99212
rect 68243 99140 68283 99174
rect 68283 99140 68317 99174
rect 68317 99140 68359 99174
rect 68243 99102 68359 99140
rect 68243 99068 68283 99102
rect 68283 99068 68317 99102
rect 68317 99068 68359 99102
rect 68243 99030 68359 99068
rect 68243 98996 68283 99030
rect 68283 98996 68317 99030
rect 68317 98996 68359 99030
rect 68243 98958 68359 98996
rect 68243 98924 68283 98958
rect 68283 98924 68317 98958
rect 68317 98924 68359 98958
rect 68243 98886 68359 98924
rect 68243 98852 68283 98886
rect 68283 98852 68317 98886
rect 68317 98852 68359 98886
rect 68243 98814 68359 98852
rect 68243 98780 68283 98814
rect 68283 98780 68317 98814
rect 68317 98780 68359 98814
rect 68243 98742 68359 98780
rect 68243 98708 68283 98742
rect 68283 98708 68317 98742
rect 68317 98708 68359 98742
rect 68243 98670 68359 98708
rect 68243 98636 68283 98670
rect 68283 98636 68317 98670
rect 68317 98636 68359 98670
rect 68243 98598 68359 98636
rect 68243 98564 68283 98598
rect 68283 98564 68317 98598
rect 68317 98564 68359 98598
rect 68243 98526 68359 98564
rect 68243 98492 68283 98526
rect 68283 98492 68317 98526
rect 68317 98492 68359 98526
rect 68243 98454 68359 98492
rect 68243 98420 68283 98454
rect 68283 98420 68317 98454
rect 68317 98420 68359 98454
rect 68243 98382 68359 98420
rect 68243 98348 68283 98382
rect 68283 98348 68317 98382
rect 68317 98348 68359 98382
rect 68243 98310 68359 98348
rect 68243 98276 68283 98310
rect 68283 98276 68317 98310
rect 68317 98276 68359 98310
rect 68243 98238 68359 98276
rect 68243 98204 68283 98238
rect 68283 98204 68317 98238
rect 68317 98204 68359 98238
rect 68243 98166 68359 98204
rect 68243 98132 68283 98166
rect 68283 98132 68317 98166
rect 68317 98132 68359 98166
rect 68243 98094 68359 98132
rect 68243 98060 68283 98094
rect 68283 98060 68317 98094
rect 68317 98060 68359 98094
rect 68243 98022 68359 98060
rect 68243 97988 68283 98022
rect 68283 97988 68317 98022
rect 68317 97988 68359 98022
rect 68243 97950 68359 97988
rect 68243 97916 68283 97950
rect 68283 97916 68317 97950
rect 68317 97916 68359 97950
rect 68243 97878 68359 97916
rect 68243 97844 68283 97878
rect 68283 97844 68317 97878
rect 68317 97844 68359 97878
rect 68243 97806 68359 97844
rect 68243 97772 68283 97806
rect 68283 97772 68317 97806
rect 68317 97772 68359 97806
rect 68243 97734 68359 97772
rect 68243 97700 68283 97734
rect 68283 97700 68317 97734
rect 68317 97700 68359 97734
rect 68243 97662 68359 97700
rect 68243 97628 68283 97662
rect 68283 97628 68317 97662
rect 68317 97628 68359 97662
rect 68243 97590 68359 97628
rect 68243 97556 68283 97590
rect 68283 97556 68317 97590
rect 68317 97556 68359 97590
rect 68243 97518 68359 97556
rect 68243 97484 68283 97518
rect 68283 97484 68317 97518
rect 68317 97484 68359 97518
rect 68243 97426 68359 97484
rect 71244 97439 71360 100755
rect 40436 95766 40488 95818
rect 41614 95762 41666 95814
rect 41831 95769 41883 95821
rect 42965 95766 43017 95818
rect 40546 94262 40598 94314
rect 41660 94248 41712 94300
rect 41873 94249 41925 94301
rect 43037 94249 43089 94301
rect 41678 92464 41730 92516
rect 41678 92400 41730 92452
rect 41678 92336 41730 92388
rect 41141 92211 41193 92263
rect 41141 92147 41193 92199
rect 41678 92272 41730 92324
rect 41678 92208 41730 92260
rect 42225 92214 42277 92266
rect 42225 92150 42277 92202
rect 40523 91577 40575 91629
rect 41678 91571 41730 91623
rect 42796 91582 42848 91634
rect 47213 87366 47265 87418
rect 47277 87366 47329 87418
rect 47341 87366 47393 87418
rect 47405 87366 47457 87418
rect 47469 87366 47521 87418
rect 47533 87366 47585 87418
rect 47597 87366 47649 87418
rect 49024 87368 49076 87420
rect 49088 87368 49140 87420
rect 49152 87368 49204 87420
rect 49216 87368 49268 87420
rect 49280 87368 49332 87420
rect 49344 87368 49396 87420
rect 49408 87368 49460 87420
rect 50819 87364 50871 87416
rect 50883 87364 50935 87416
rect 50947 87364 50999 87416
rect 51011 87364 51063 87416
rect 51075 87364 51127 87416
rect 51139 87364 51191 87416
rect 51203 87364 51255 87416
rect 52618 87362 52670 87414
rect 52682 87362 52734 87414
rect 52746 87362 52798 87414
rect 52810 87362 52862 87414
rect 52874 87362 52926 87414
rect 52938 87362 52990 87414
rect 53002 87362 53054 87414
rect 50185 87018 50365 87198
rect 54409 87366 54461 87418
rect 54473 87366 54525 87418
rect 54537 87366 54589 87418
rect 54601 87366 54653 87418
rect 54665 87366 54717 87418
rect 54729 87366 54781 87418
rect 54793 87366 54845 87418
rect 56211 87362 56263 87414
rect 56275 87362 56327 87414
rect 56339 87362 56391 87414
rect 56403 87362 56455 87414
rect 56467 87362 56519 87414
rect 56531 87362 56583 87414
rect 56595 87362 56647 87414
rect 57866 87044 58366 87224
rect 48543 78559 48595 78611
rect 50234 78560 50286 78612
rect 51939 78559 51991 78611
rect 53735 78559 53787 78611
rect 55564 78559 55616 78611
rect 47421 78367 47473 78419
rect 47485 78367 47537 78419
rect 47549 78367 47601 78419
rect 49216 78366 49268 78418
rect 49280 78366 49332 78418
rect 49344 78366 49396 78418
rect 51016 78368 51068 78420
rect 51080 78368 51132 78420
rect 51144 78368 51196 78420
rect 52814 78367 52866 78419
rect 52878 78367 52930 78419
rect 52942 78367 52994 78419
rect 54612 78368 54664 78420
rect 54676 78368 54728 78420
rect 54740 78368 54792 78420
rect 56415 78367 56467 78419
rect 56479 78367 56531 78419
rect 56543 78367 56595 78419
rect 57276 78368 57328 78420
rect 42317 77564 42369 77616
rect 42381 77564 42433 77616
rect 49550 77564 49602 77616
rect 50111 77564 50163 77616
rect 50175 77564 50227 77616
rect 57469 84768 57585 84830
rect 57469 84734 57504 84768
rect 57504 84734 57538 84768
rect 57538 84734 57585 84768
rect 57469 84696 57585 84734
rect 57469 84662 57504 84696
rect 57504 84662 57538 84696
rect 57538 84662 57585 84696
rect 57469 84624 57585 84662
rect 57469 84590 57504 84624
rect 57504 84590 57538 84624
rect 57538 84590 57585 84624
rect 57469 84552 57585 84590
rect 57469 84518 57504 84552
rect 57504 84518 57538 84552
rect 57538 84518 57585 84552
rect 57469 84480 57585 84518
rect 57469 84446 57504 84480
rect 57504 84446 57538 84480
rect 57538 84446 57585 84480
rect 57469 84408 57585 84446
rect 57469 84374 57504 84408
rect 57504 84374 57538 84408
rect 57538 84374 57585 84408
rect 57469 84336 57585 84374
rect 57469 84302 57504 84336
rect 57504 84302 57538 84336
rect 57538 84302 57585 84336
rect 57469 84264 57585 84302
rect 57469 84230 57504 84264
rect 57504 84230 57538 84264
rect 57538 84230 57585 84264
rect 57469 84192 57585 84230
rect 57469 84158 57504 84192
rect 57504 84158 57538 84192
rect 57538 84158 57585 84192
rect 57469 84120 57585 84158
rect 57469 84086 57504 84120
rect 57504 84086 57538 84120
rect 57538 84086 57585 84120
rect 57469 84048 57585 84086
rect 57469 84014 57504 84048
rect 57504 84014 57538 84048
rect 57538 84014 57585 84048
rect 57469 83976 57585 84014
rect 57469 83942 57504 83976
rect 57504 83942 57538 83976
rect 57538 83942 57585 83976
rect 57469 83904 57585 83942
rect 57469 83870 57504 83904
rect 57504 83870 57538 83904
rect 57538 83870 57585 83904
rect 57469 83832 57585 83870
rect 57469 83798 57504 83832
rect 57504 83798 57538 83832
rect 57538 83798 57585 83832
rect 57469 83760 57585 83798
rect 57469 83726 57504 83760
rect 57504 83726 57538 83760
rect 57538 83726 57585 83760
rect 57469 83688 57585 83726
rect 57469 83654 57504 83688
rect 57504 83654 57538 83688
rect 57538 83654 57585 83688
rect 57469 83616 57585 83654
rect 57469 83582 57504 83616
rect 57504 83582 57538 83616
rect 57538 83582 57585 83616
rect 57469 83544 57585 83582
rect 57469 83510 57504 83544
rect 57504 83510 57538 83544
rect 57538 83510 57585 83544
rect 57469 83472 57585 83510
rect 57469 83438 57504 83472
rect 57504 83438 57538 83472
rect 57538 83438 57585 83472
rect 57469 83400 57585 83438
rect 57469 83366 57504 83400
rect 57504 83366 57538 83400
rect 57538 83366 57585 83400
rect 57469 83328 57585 83366
rect 57469 83294 57504 83328
rect 57504 83294 57538 83328
rect 57538 83294 57585 83328
rect 57469 83256 57585 83294
rect 57469 83222 57504 83256
rect 57504 83222 57538 83256
rect 57538 83222 57585 83256
rect 57469 83184 57585 83222
rect 57469 83150 57504 83184
rect 57504 83150 57538 83184
rect 57538 83150 57585 83184
rect 57469 83112 57585 83150
rect 57469 83078 57504 83112
rect 57504 83078 57538 83112
rect 57538 83078 57585 83112
rect 57469 83040 57585 83078
rect 57469 83006 57504 83040
rect 57504 83006 57538 83040
rect 57538 83006 57585 83040
rect 57469 82968 57585 83006
rect 57469 82934 57504 82968
rect 57504 82934 57538 82968
rect 57538 82934 57585 82968
rect 57469 82896 57585 82934
rect 57469 82862 57504 82896
rect 57504 82862 57538 82896
rect 57538 82862 57585 82896
rect 57469 82824 57585 82862
rect 57469 82790 57504 82824
rect 57504 82790 57538 82824
rect 57538 82790 57585 82824
rect 57469 82752 57585 82790
rect 57469 82718 57504 82752
rect 57504 82718 57538 82752
rect 57538 82718 57585 82752
rect 57469 82680 57585 82718
rect 57469 82646 57504 82680
rect 57504 82646 57538 82680
rect 57538 82646 57585 82680
rect 57469 82608 57585 82646
rect 57469 82574 57504 82608
rect 57504 82574 57538 82608
rect 57538 82574 57585 82608
rect 57469 82536 57585 82574
rect 57469 82502 57504 82536
rect 57504 82502 57538 82536
rect 57538 82502 57585 82536
rect 57469 82464 57585 82502
rect 57469 82430 57504 82464
rect 57504 82430 57538 82464
rect 57538 82430 57585 82464
rect 57469 82392 57585 82430
rect 57469 82358 57504 82392
rect 57504 82358 57538 82392
rect 57538 82358 57585 82392
rect 57469 82320 57585 82358
rect 57469 82286 57504 82320
rect 57504 82286 57538 82320
rect 57538 82286 57585 82320
rect 57469 82248 57585 82286
rect 57469 82214 57504 82248
rect 57504 82214 57538 82248
rect 57538 82214 57585 82248
rect 57469 82176 57585 82214
rect 57469 82142 57504 82176
rect 57504 82142 57538 82176
rect 57538 82142 57585 82176
rect 57469 82104 57585 82142
rect 57469 82070 57504 82104
rect 57504 82070 57538 82104
rect 57538 82070 57585 82104
rect 57469 82032 57585 82070
rect 57469 81998 57504 82032
rect 57504 81998 57538 82032
rect 57538 81998 57585 82032
rect 57469 81960 57585 81998
rect 57469 81926 57504 81960
rect 57504 81926 57538 81960
rect 57538 81926 57585 81960
rect 57469 81888 57585 81926
rect 57469 81854 57504 81888
rect 57504 81854 57538 81888
rect 57538 81854 57585 81888
rect 57469 81816 57585 81854
rect 57469 81782 57504 81816
rect 57504 81782 57538 81816
rect 57538 81782 57585 81816
rect 57469 81744 57585 81782
rect 57469 81710 57504 81744
rect 57504 81710 57538 81744
rect 57538 81710 57585 81744
rect 57469 81672 57585 81710
rect 57469 81638 57504 81672
rect 57504 81638 57538 81672
rect 57538 81638 57585 81672
rect 57469 81600 57585 81638
rect 57469 81566 57504 81600
rect 57504 81566 57538 81600
rect 57538 81566 57585 81600
rect 57469 81528 57585 81566
rect 57469 81494 57504 81528
rect 57504 81494 57538 81528
rect 57538 81494 57585 81528
rect 57469 81456 57585 81494
rect 57469 81422 57504 81456
rect 57504 81422 57538 81456
rect 57538 81422 57585 81456
rect 57469 81384 57585 81422
rect 57469 81350 57504 81384
rect 57504 81350 57538 81384
rect 57538 81350 57585 81384
rect 57469 81312 57585 81350
rect 57469 81278 57504 81312
rect 57504 81278 57538 81312
rect 57538 81278 57585 81312
rect 57469 81240 57585 81278
rect 57469 81206 57504 81240
rect 57504 81206 57538 81240
rect 57538 81206 57585 81240
rect 57469 81168 57585 81206
rect 57469 81134 57504 81168
rect 57504 81134 57538 81168
rect 57538 81134 57585 81168
rect 57469 81096 57585 81134
rect 57469 81062 57504 81096
rect 57504 81062 57538 81096
rect 57538 81062 57585 81096
rect 57469 81024 57585 81062
rect 57469 80990 57504 81024
rect 57504 80990 57538 81024
rect 57538 80990 57585 81024
rect 57469 80952 57585 80990
rect 57469 80918 57504 80952
rect 57504 80918 57538 80952
rect 57538 80918 57585 80952
rect 57469 80880 57585 80918
rect 57469 80846 57504 80880
rect 57504 80846 57538 80880
rect 57538 80846 57585 80880
rect 57469 80808 57585 80846
rect 57469 80774 57504 80808
rect 57504 80774 57538 80808
rect 57538 80774 57585 80808
rect 57469 80736 57585 80774
rect 57469 80702 57504 80736
rect 57504 80702 57538 80736
rect 57538 80702 57585 80736
rect 57469 80664 57585 80702
rect 57469 80630 57504 80664
rect 57504 80630 57538 80664
rect 57538 80630 57585 80664
rect 57469 80592 57585 80630
rect 57469 80558 57504 80592
rect 57504 80558 57538 80592
rect 57538 80558 57585 80592
rect 57469 80520 57585 80558
rect 57469 80486 57504 80520
rect 57504 80486 57538 80520
rect 57538 80486 57585 80520
rect 57469 80448 57585 80486
rect 57469 80414 57504 80448
rect 57504 80414 57538 80448
rect 57538 80414 57585 80448
rect 57469 80376 57585 80414
rect 57469 80342 57504 80376
rect 57504 80342 57538 80376
rect 57538 80342 57585 80376
rect 57469 80304 57585 80342
rect 57469 80270 57504 80304
rect 57504 80270 57538 80304
rect 57538 80270 57585 80304
rect 57469 80232 57585 80270
rect 57469 80198 57504 80232
rect 57504 80198 57538 80232
rect 57538 80198 57585 80232
rect 57469 80160 57585 80198
rect 57469 80126 57504 80160
rect 57504 80126 57538 80160
rect 57538 80126 57585 80160
rect 57469 80088 57585 80126
rect 57469 80054 57504 80088
rect 57504 80054 57538 80088
rect 57538 80054 57585 80088
rect 57469 80016 57585 80054
rect 57469 79982 57504 80016
rect 57504 79982 57538 80016
rect 57538 79982 57585 80016
rect 57469 79944 57585 79982
rect 57469 79910 57504 79944
rect 57504 79910 57538 79944
rect 57538 79910 57585 79944
rect 57469 79872 57585 79910
rect 57469 79838 57504 79872
rect 57504 79838 57538 79872
rect 57538 79838 57585 79872
rect 57469 79800 57585 79838
rect 57469 79766 57504 79800
rect 57504 79766 57538 79800
rect 57538 79766 57585 79800
rect 57469 79728 57585 79766
rect 57469 79694 57504 79728
rect 57504 79694 57538 79728
rect 57538 79694 57585 79728
rect 57469 79656 57585 79694
rect 57469 79622 57504 79656
rect 57504 79622 57538 79656
rect 57538 79622 57585 79656
rect 57469 79584 57585 79622
rect 57469 79550 57504 79584
rect 57504 79550 57538 79584
rect 57538 79550 57585 79584
rect 57469 79512 57585 79550
rect 57469 79478 57504 79512
rect 57504 79478 57538 79512
rect 57538 79478 57585 79512
rect 57469 79440 57585 79478
rect 57469 79406 57504 79440
rect 57504 79406 57538 79440
rect 57538 79406 57585 79440
rect 57469 79368 57585 79406
rect 57469 79334 57504 79368
rect 57504 79334 57538 79368
rect 57538 79334 57585 79368
rect 57469 79296 57585 79334
rect 57469 79262 57504 79296
rect 57504 79262 57538 79296
rect 57538 79262 57585 79296
rect 57469 79224 57585 79262
rect 57469 79190 57504 79224
rect 57504 79190 57538 79224
rect 57538 79190 57585 79224
rect 57469 79152 57585 79190
rect 57469 79118 57504 79152
rect 57504 79118 57538 79152
rect 57538 79118 57585 79152
rect 57469 79080 57585 79118
rect 57469 79046 57504 79080
rect 57504 79046 57538 79080
rect 57538 79046 57585 79080
rect 57469 79008 57585 79046
rect 57469 78974 57504 79008
rect 57504 78974 57538 79008
rect 57538 78974 57585 79008
rect 57469 78936 57585 78974
rect 57469 78902 57504 78936
rect 57504 78902 57538 78936
rect 57538 78902 57585 78936
rect 57469 78864 57585 78902
rect 57469 78830 57504 78864
rect 57504 78830 57538 78864
rect 57538 78830 57585 78864
rect 57469 78792 57585 78830
rect 57469 78758 57504 78792
rect 57504 78758 57538 78792
rect 57538 78758 57585 78792
rect 57469 78720 57585 78758
rect 57469 78686 57504 78720
rect 57504 78686 57538 78720
rect 57538 78686 57585 78720
rect 57469 78648 57585 78686
rect 57469 78614 57504 78648
rect 57504 78614 57538 78648
rect 57538 78614 57585 78648
rect 57469 78576 57585 78614
rect 57469 78542 57504 78576
rect 57504 78542 57538 78576
rect 57538 78542 57585 78576
rect 57469 78504 57585 78542
rect 57469 78470 57504 78504
rect 57504 78470 57538 78504
rect 57538 78470 57585 78504
rect 57469 78432 57585 78470
rect 57469 78398 57504 78432
rect 57504 78398 57538 78432
rect 57538 78398 57585 78432
rect 57469 78360 57585 78398
rect 57469 78326 57504 78360
rect 57504 78326 57538 78360
rect 57538 78326 57585 78360
rect 57469 78288 57585 78326
rect 57469 78254 57504 78288
rect 57504 78254 57538 78288
rect 57538 78254 57585 78288
rect 57469 78216 57585 78254
rect 57469 78182 57504 78216
rect 57504 78182 57538 78216
rect 57538 78182 57585 78216
rect 57469 78144 57585 78182
rect 57469 78110 57504 78144
rect 57504 78110 57538 78144
rect 57538 78110 57585 78144
rect 57469 78072 57585 78110
rect 57469 78038 57504 78072
rect 57504 78038 57538 78072
rect 57538 78038 57585 78072
rect 57469 78000 57585 78038
rect 57469 77966 57504 78000
rect 57504 77966 57538 78000
rect 57538 77966 57585 78000
rect 57469 77928 57585 77966
rect 57469 77894 57504 77928
rect 57504 77894 57538 77928
rect 57538 77894 57585 77928
rect 57469 77856 57585 77894
rect 57469 77822 57504 77856
rect 57504 77822 57538 77856
rect 57538 77822 57585 77856
rect 57469 77784 57585 77822
rect 57469 77750 57504 77784
rect 57504 77750 57538 77784
rect 57538 77750 57585 77784
rect 57469 77712 57585 77750
rect 57469 77678 57504 77712
rect 57504 77678 57538 77712
rect 57538 77678 57585 77712
rect 57469 77640 57585 77678
rect 57469 77606 57504 77640
rect 57504 77606 57538 77640
rect 57538 77606 57585 77640
rect 57469 77568 57585 77606
rect 57469 77534 57504 77568
rect 57504 77534 57538 77568
rect 57538 77534 57585 77568
rect 57469 77496 57585 77534
rect 57469 77462 57504 77496
rect 57504 77462 57538 77496
rect 57538 77462 57585 77496
rect 57469 77424 57585 77462
rect 57469 77390 57504 77424
rect 57504 77390 57538 77424
rect 57538 77390 57585 77424
rect 57469 77352 57585 77390
rect 57469 77318 57504 77352
rect 57504 77318 57538 77352
rect 57538 77318 57585 77352
rect 57469 77280 57585 77318
rect 57469 77246 57504 77280
rect 57504 77246 57538 77280
rect 57538 77246 57585 77280
rect 57469 77208 57585 77246
rect 57469 77174 57504 77208
rect 57504 77174 57538 77208
rect 57538 77174 57585 77208
rect 57469 77162 57585 77174
rect 47702 76956 47754 77008
rect 47766 76956 47818 77008
rect 48256 75191 48308 75243
rect 48256 75127 48308 75179
rect 48256 75063 48308 75115
rect 47702 74901 47754 74953
rect 47766 74901 47818 74953
rect 50111 74899 50163 74951
rect 50175 74899 50227 74951
rect 51416 75010 53196 75086
rect 53735 75010 54555 75065
rect 55442 75010 56326 75055
rect 51416 74976 51487 75010
rect 51487 74976 51521 75010
rect 51521 74976 51559 75010
rect 51559 74976 51593 75010
rect 51593 74976 51631 75010
rect 51631 74976 51665 75010
rect 51665 74976 51703 75010
rect 51703 74976 51737 75010
rect 51737 74976 51775 75010
rect 51775 74976 51809 75010
rect 51809 74976 51847 75010
rect 51847 74976 51881 75010
rect 51881 74976 51919 75010
rect 51919 74976 51953 75010
rect 51953 74976 51991 75010
rect 51991 74976 52025 75010
rect 52025 74976 52063 75010
rect 52063 74976 52097 75010
rect 52097 74976 52135 75010
rect 52135 74976 52169 75010
rect 52169 74976 52207 75010
rect 52207 74976 52241 75010
rect 52241 74976 52279 75010
rect 52279 74976 52313 75010
rect 52313 74976 52351 75010
rect 52351 74976 52385 75010
rect 52385 74976 52423 75010
rect 52423 74976 52457 75010
rect 52457 74976 52495 75010
rect 52495 74976 52529 75010
rect 52529 74976 52567 75010
rect 52567 74976 52601 75010
rect 52601 74976 52639 75010
rect 52639 74976 52673 75010
rect 52673 74976 52711 75010
rect 52711 74976 52745 75010
rect 52745 74976 52783 75010
rect 52783 74976 52817 75010
rect 52817 74976 52855 75010
rect 52855 74976 52889 75010
rect 52889 74976 52927 75010
rect 52927 74976 52961 75010
rect 52961 74976 52999 75010
rect 52999 74976 53033 75010
rect 53033 74976 53071 75010
rect 53071 74976 53105 75010
rect 53105 74976 53143 75010
rect 53143 74976 53177 75010
rect 53177 74976 53196 75010
rect 53735 74976 53753 75010
rect 53753 74976 53791 75010
rect 53791 74976 53825 75010
rect 53825 74976 53863 75010
rect 53863 74976 53897 75010
rect 53897 74976 53935 75010
rect 53935 74976 53969 75010
rect 53969 74976 54007 75010
rect 54007 74976 54041 75010
rect 54041 74976 54079 75010
rect 54079 74976 54113 75010
rect 54113 74976 54151 75010
rect 54151 74976 54185 75010
rect 54185 74976 54223 75010
rect 54223 74976 54257 75010
rect 54257 74976 54295 75010
rect 54295 74976 54329 75010
rect 54329 74976 54367 75010
rect 54367 74976 54401 75010
rect 54401 74976 54439 75010
rect 54439 74976 54473 75010
rect 54473 74976 54511 75010
rect 54511 74976 54545 75010
rect 54545 74976 54555 75010
rect 55442 74976 55447 75010
rect 55447 74976 55481 75010
rect 55481 74976 55519 75010
rect 55519 74976 55553 75010
rect 55553 74976 55591 75010
rect 55591 74976 55625 75010
rect 55625 74976 55663 75010
rect 55663 74976 55697 75010
rect 55697 74976 55735 75010
rect 55735 74976 55769 75010
rect 55769 74976 55807 75010
rect 55807 74976 55841 75010
rect 55841 74976 55879 75010
rect 55879 74976 55913 75010
rect 55913 74976 55951 75010
rect 55951 74976 55985 75010
rect 55985 74976 56023 75010
rect 56023 74976 56057 75010
rect 56057 74976 56095 75010
rect 56095 74976 56129 75010
rect 56129 74976 56167 75010
rect 56167 74976 56201 75010
rect 56201 74976 56239 75010
rect 56239 74976 56273 75010
rect 56273 74976 56311 75010
rect 56311 74976 56326 75010
rect 51416 74906 53196 74976
rect 53735 74949 54555 74976
rect 55442 74939 56326 74976
rect 48241 74740 48293 74792
rect 48241 74676 48293 74728
rect 48241 74612 48293 74664
rect 48241 74548 48293 74600
rect 48241 74484 48293 74536
rect 48241 74420 48293 74472
rect 30042 73684 30094 73736
rect 30106 73684 30158 73736
rect 30170 73684 30222 73736
rect 30234 73684 30286 73736
rect 30298 73684 30350 73736
rect 30689 73420 30741 73429
rect 30753 73420 30805 73429
rect 30817 73420 30869 73429
rect 30881 73420 30933 73429
rect 30689 73386 30717 73420
rect 30717 73386 30741 73420
rect 30753 73386 30789 73420
rect 30789 73386 30805 73420
rect 30817 73386 30823 73420
rect 30823 73386 30861 73420
rect 30861 73386 30869 73420
rect 30881 73386 30895 73420
rect 30895 73386 30933 73420
rect 30689 73377 30741 73386
rect 30753 73377 30805 73386
rect 30817 73377 30869 73386
rect 30881 73377 30933 73386
rect 31040 73435 31047 73440
rect 31047 73435 31081 73440
rect 31081 73435 31092 73440
rect 31040 73388 31092 73435
rect 31128 73142 31180 73194
rect 31192 73142 31244 73194
rect 31256 73142 31308 73194
rect 31320 73142 31372 73194
rect 31384 73142 31436 73194
rect 51164 71804 51344 74736
rect 57025 74735 57205 74783
rect 57025 74701 57119 74735
rect 57119 74701 57153 74735
rect 57153 74701 57205 74735
rect 57025 74663 57205 74701
rect 57025 74629 57119 74663
rect 57119 74629 57153 74663
rect 57153 74629 57205 74663
rect 57025 74591 57205 74629
rect 57025 74557 57119 74591
rect 57119 74557 57153 74591
rect 57153 74557 57205 74591
rect 57025 74519 57205 74557
rect 57025 74485 57119 74519
rect 57119 74485 57153 74519
rect 57153 74485 57205 74519
rect 57025 74447 57205 74485
rect 57025 74413 57119 74447
rect 57119 74413 57153 74447
rect 57153 74413 57205 74447
rect 57025 74375 57205 74413
rect 57025 74341 57119 74375
rect 57119 74341 57153 74375
rect 57153 74341 57205 74375
rect 57025 74303 57205 74341
rect 57025 74269 57119 74303
rect 57119 74269 57153 74303
rect 57153 74269 57205 74303
rect 57025 74231 57205 74269
rect 57025 74197 57119 74231
rect 57119 74197 57153 74231
rect 57153 74197 57205 74231
rect 57025 74159 57205 74197
rect 57025 74125 57119 74159
rect 57119 74125 57153 74159
rect 57153 74125 57205 74159
rect 57025 74087 57205 74125
rect 57025 74053 57119 74087
rect 57119 74053 57153 74087
rect 57153 74053 57205 74087
rect 57025 74015 57205 74053
rect 57025 73981 57119 74015
rect 57119 73981 57153 74015
rect 57153 73981 57205 74015
rect 57025 73943 57205 73981
rect 57025 73909 57119 73943
rect 57119 73909 57153 73943
rect 57153 73909 57205 73943
rect 57025 73871 57205 73909
rect 57025 73837 57119 73871
rect 57119 73837 57153 73871
rect 57153 73837 57205 73871
rect 57025 73799 57205 73837
rect 57025 73765 57119 73799
rect 57119 73765 57153 73799
rect 57153 73765 57205 73799
rect 57025 73727 57205 73765
rect 57025 73693 57119 73727
rect 57119 73693 57153 73727
rect 57153 73693 57205 73727
rect 57025 73655 57205 73693
rect 57025 73621 57119 73655
rect 57119 73621 57153 73655
rect 57153 73621 57205 73655
rect 57025 73583 57205 73621
rect 57025 73549 57119 73583
rect 57119 73549 57153 73583
rect 57153 73549 57205 73583
rect 57025 73511 57205 73549
rect 57025 73477 57119 73511
rect 57119 73477 57153 73511
rect 57153 73477 57205 73511
rect 57025 73439 57205 73477
rect 57025 73405 57119 73439
rect 57119 73405 57153 73439
rect 57153 73405 57205 73439
rect 57025 73367 57205 73405
rect 57025 73333 57119 73367
rect 57119 73333 57153 73367
rect 57153 73333 57205 73367
rect 57025 73295 57205 73333
rect 57025 73261 57119 73295
rect 57119 73261 57153 73295
rect 57153 73261 57205 73295
rect 57025 73223 57205 73261
rect 57025 73189 57119 73223
rect 57119 73189 57153 73223
rect 57153 73189 57205 73223
rect 57025 73151 57205 73189
rect 57025 73117 57119 73151
rect 57119 73117 57153 73151
rect 57153 73117 57205 73151
rect 57025 73079 57205 73117
rect 57025 73045 57119 73079
rect 57119 73045 57153 73079
rect 57153 73045 57205 73079
rect 57025 73007 57205 73045
rect 57025 72973 57119 73007
rect 57119 72973 57153 73007
rect 57153 72973 57205 73007
rect 57025 72935 57205 72973
rect 57025 72901 57119 72935
rect 57119 72901 57153 72935
rect 57153 72901 57205 72935
rect 57025 72863 57205 72901
rect 57025 72829 57119 72863
rect 57119 72829 57153 72863
rect 57153 72829 57205 72863
rect 57025 72791 57205 72829
rect 57025 72757 57119 72791
rect 57119 72757 57153 72791
rect 57153 72757 57205 72791
rect 57025 72719 57205 72757
rect 57025 72685 57119 72719
rect 57119 72685 57153 72719
rect 57153 72685 57205 72719
rect 57025 72647 57205 72685
rect 57025 72613 57119 72647
rect 57119 72613 57153 72647
rect 57153 72613 57205 72647
rect 57025 72575 57205 72613
rect 57025 72541 57119 72575
rect 57119 72541 57153 72575
rect 57153 72541 57205 72575
rect 57025 72503 57205 72541
rect 57025 72469 57119 72503
rect 57119 72469 57153 72503
rect 57153 72469 57205 72503
rect 57025 72431 57205 72469
rect 57025 72397 57119 72431
rect 57119 72397 57153 72431
rect 57153 72397 57205 72431
rect 57025 72359 57205 72397
rect 57025 72325 57119 72359
rect 57119 72325 57153 72359
rect 57153 72325 57205 72359
rect 57025 72287 57205 72325
rect 57025 72253 57119 72287
rect 57119 72253 57153 72287
rect 57153 72253 57205 72287
rect 57025 72215 57205 72253
rect 57025 72181 57119 72215
rect 57119 72181 57153 72215
rect 57153 72181 57205 72215
rect 57025 72143 57205 72181
rect 57025 72109 57119 72143
rect 57119 72109 57153 72143
rect 57153 72109 57205 72143
rect 57025 72071 57205 72109
rect 57025 72037 57119 72071
rect 57119 72037 57153 72071
rect 57153 72037 57205 72071
rect 57025 71999 57205 72037
rect 57025 71965 57119 71999
rect 57119 71965 57153 71999
rect 57153 71965 57205 71999
rect 57025 71927 57205 71965
rect 57025 71893 57119 71927
rect 57119 71893 57153 71927
rect 57153 71893 57205 71927
rect 57025 71855 57205 71893
rect 57025 71821 57119 71855
rect 57119 71821 57153 71855
rect 57153 71821 57205 71855
rect 57025 71787 57205 71821
rect 67272 71662 67644 84834
rect 30029 67266 30081 67318
rect 30029 67202 30081 67254
rect 30029 67138 30081 67190
rect 30029 67074 30081 67126
rect 30029 67010 30081 67062
rect 43631 67025 43683 67077
rect 30029 66946 30081 66998
rect 30029 66882 30081 66934
rect 30029 66818 30081 66870
rect 30029 66125 30081 66177
rect 30029 66061 30081 66113
rect 30029 65997 30081 66049
rect 30029 65933 30081 65985
rect 30029 65869 30081 65921
rect 30029 65805 30081 65857
rect 30029 65741 30081 65793
rect 30029 65677 30081 65729
rect 30029 65613 30081 65665
rect 30029 65549 30081 65601
rect 30029 65485 30081 65537
rect 30029 65421 30081 65473
rect 30029 65357 30081 65409
rect 30029 65293 30081 65345
rect 30029 65229 30081 65281
rect 30029 65165 30081 65217
rect 30029 65101 30081 65153
rect 30029 65037 30081 65089
rect 30034 64599 30086 64651
rect 30034 64535 30086 64587
rect 30034 64471 30086 64523
rect 30034 64407 30086 64459
rect 30034 64343 30086 64395
rect 30034 64279 30086 64331
rect 30034 64215 30086 64267
rect 30034 64151 30086 64203
rect 30034 64087 30086 64139
rect 30034 64023 30086 64075
rect 30034 63959 30086 64011
rect 30034 63895 30086 63947
rect 30034 63831 30086 63883
rect 30034 63767 30086 63819
rect 30034 63703 30086 63755
rect 30034 63639 30086 63691
rect 30034 63575 30086 63627
rect 30034 63511 30086 63563
rect 38223 63490 38275 63542
rect 38223 63426 38275 63478
rect 38223 63362 38275 63414
rect 38223 63298 38275 63350
rect 38223 63234 38275 63286
rect 25288 63136 25340 63172
rect 25288 63120 25299 63136
rect 25299 63120 25333 63136
rect 25333 63120 25340 63136
rect 38223 63170 38275 63222
rect 25288 63102 25299 63108
rect 25299 63102 25333 63108
rect 25333 63102 25340 63108
rect 25288 63064 25340 63102
rect 25288 63056 25299 63064
rect 25299 63056 25333 63064
rect 25333 63056 25340 63064
rect 25288 63030 25299 63044
rect 25299 63030 25333 63044
rect 25333 63030 25340 63044
rect 25288 62992 25340 63030
rect 25288 62958 25299 62980
rect 25299 62958 25333 62980
rect 25333 62958 25340 62980
rect 25288 62928 25340 62958
rect 25288 62886 25299 62916
rect 25299 62886 25333 62916
rect 25333 62886 25340 62916
rect 25288 62864 25340 62886
rect 25289 62572 25341 62617
rect 25289 62565 25299 62572
rect 25299 62565 25333 62572
rect 25333 62565 25341 62572
rect 25289 62538 25299 62553
rect 25299 62538 25333 62553
rect 25333 62538 25341 62553
rect 25289 62501 25341 62538
rect 25289 62466 25299 62489
rect 25299 62466 25333 62489
rect 25333 62466 25341 62489
rect 25289 62437 25341 62466
rect 25289 62394 25299 62425
rect 25299 62394 25333 62425
rect 25333 62394 25341 62425
rect 25289 62373 25341 62394
rect 25289 62356 25341 62361
rect 25289 62322 25299 62356
rect 25299 62322 25333 62356
rect 25333 62322 25341 62356
rect 25289 62309 25341 62322
rect 25289 62284 25341 62297
rect 25289 62250 25299 62284
rect 25299 62250 25333 62284
rect 25333 62250 25341 62284
rect 25289 62245 25341 62250
rect 30028 63088 30080 63140
rect 30028 63024 30080 63076
rect 30028 62960 30080 63012
rect 30028 62896 30080 62948
rect 30028 62832 30080 62884
rect 30028 62768 30080 62820
rect 30028 62704 30080 62756
rect 30028 62640 30080 62692
rect 30028 62576 30080 62628
rect 30028 62512 30080 62564
rect 30028 62448 30080 62500
rect 27494 62377 27546 62429
rect 27558 62377 27610 62429
rect 27622 62377 27674 62429
rect 27686 62377 27738 62429
rect 27750 62377 27802 62429
rect 27814 62377 27866 62429
rect 27878 62377 27930 62429
rect 30028 62384 30080 62436
rect 30028 62320 30080 62372
rect 25289 62181 25341 62233
rect 26070 62220 26122 62272
rect 26134 62220 26186 62272
rect 30028 62256 30080 62308
rect 38223 63106 38275 63158
rect 38223 63042 38275 63094
rect 38223 62978 38275 63030
rect 38223 62914 38275 62966
rect 38223 62850 38275 62902
rect 38223 62786 38275 62838
rect 38223 62722 38275 62774
rect 38223 62658 38275 62710
rect 38223 62594 38275 62646
rect 38223 62530 38275 62582
rect 38223 62466 38275 62518
rect 38223 62402 38275 62454
rect 38223 62338 38275 62390
rect 38223 62274 38275 62326
rect 38223 62210 38275 62262
rect 38223 62146 38275 62198
rect 38223 62082 38275 62134
rect 38223 62018 38275 62070
rect 38223 61954 38275 62006
rect 38223 61890 38275 61942
rect 38223 61826 38275 61878
rect 38223 61762 38275 61814
rect 38223 61698 38275 61750
rect 38223 61634 38275 61686
rect 21604 61382 21784 61562
rect 38223 61570 38275 61622
rect 38223 61506 38275 61558
rect 26901 61439 26953 61491
rect 26965 61439 27017 61491
rect 38223 61442 38275 61494
rect 38223 61378 38275 61430
rect 27446 61287 27498 61339
rect 27510 61287 27562 61339
rect 27574 61287 27626 61339
rect 27638 61287 27690 61339
rect 27702 61287 27754 61339
rect 27766 61287 27818 61339
rect 27830 61287 27882 61339
rect 27894 61287 27946 61339
rect 30031 61321 30083 61373
rect 30031 61257 30083 61309
rect 30031 61193 30083 61245
rect 30031 61129 30083 61181
rect 30031 61065 30083 61117
rect 30031 61001 30083 61053
rect 30031 60937 30083 60989
rect 30031 60873 30083 60925
rect 30031 60809 30083 60861
rect 30031 60745 30083 60797
rect 30031 60681 30083 60733
rect 30031 60617 30083 60669
rect 30031 60553 30083 60605
rect 30031 60489 30083 60541
rect 38223 61314 38275 61366
rect 38223 61250 38275 61302
rect 38223 61186 38275 61238
rect 38223 61122 38275 61174
rect 38223 61058 38275 61110
rect 38223 60994 38275 61046
rect 38223 60930 38275 60982
rect 38223 60866 38275 60918
rect 38223 60802 38275 60854
rect 38223 60738 38275 60790
rect 38223 60674 38275 60726
rect 38223 60610 38275 60662
rect 38223 60546 38275 60598
rect 38223 60482 38275 60534
rect 38223 60418 38275 60470
rect 38223 60354 38275 60406
rect 38223 60290 38275 60342
rect 38223 60226 38275 60278
rect 30031 60112 30083 60164
rect 38223 60162 38275 60214
rect 30031 60048 30083 60100
rect 30031 59984 30083 60036
rect 30031 59920 30083 59972
rect 30031 59856 30083 59908
rect 30031 59792 30083 59844
rect 30031 59728 30083 59780
rect 30031 59664 30083 59716
rect 30031 59600 30083 59652
rect 30031 59536 30083 59588
rect 30031 59472 30083 59524
rect 30031 59408 30083 59460
rect 30031 59344 30083 59396
rect 30031 59280 30083 59332
rect 30031 59216 30083 59268
rect 30031 59152 30083 59204
rect 30031 59088 30083 59140
rect 30031 59024 30083 59076
rect 30028 58634 30080 58686
rect 30028 58570 30080 58622
rect 30028 58506 30080 58558
rect 30028 58442 30080 58494
rect 30028 58378 30080 58430
rect 30028 58314 30080 58366
rect 30028 58250 30080 58302
rect 30028 58186 30080 58238
rect 30028 58122 30080 58174
rect 30028 58058 30080 58110
rect 30028 57994 30080 58046
rect 30028 57930 30080 57982
rect 30028 57866 30080 57918
rect 30028 57802 30080 57854
rect 30028 57738 30080 57790
rect 30028 57674 30080 57726
rect 30028 57610 30080 57662
rect 30028 57546 30080 57598
rect 30023 56852 30075 56904
rect 30023 56788 30075 56840
rect 30023 56724 30075 56776
rect 30023 56660 30075 56712
rect 30023 56596 30075 56648
rect 30023 56532 30075 56584
rect 30023 56468 30075 56520
rect 30023 56404 30075 56456
rect 44407 66362 44459 66414
rect 51181 63842 51361 70294
rect 47702 63769 47754 63821
rect 47766 63769 47818 63821
rect 50111 63769 50163 63821
rect 50175 63769 50227 63821
rect 47731 58640 47783 58692
rect 51432 63795 56924 63868
rect 51432 63761 51474 63795
rect 51474 63761 51508 63795
rect 51508 63761 51546 63795
rect 51546 63761 51580 63795
rect 51580 63761 51618 63795
rect 51618 63761 51652 63795
rect 51652 63761 51690 63795
rect 51690 63761 51724 63795
rect 51724 63761 51762 63795
rect 51762 63761 51796 63795
rect 51796 63761 51834 63795
rect 51834 63761 51868 63795
rect 51868 63761 51906 63795
rect 51906 63761 51940 63795
rect 51940 63761 51978 63795
rect 51978 63761 52012 63795
rect 52012 63761 52050 63795
rect 52050 63761 52084 63795
rect 52084 63761 52122 63795
rect 52122 63761 52156 63795
rect 52156 63761 52194 63795
rect 52194 63761 52228 63795
rect 52228 63761 52266 63795
rect 52266 63761 52300 63795
rect 52300 63761 52338 63795
rect 52338 63761 52372 63795
rect 52372 63761 52410 63795
rect 52410 63761 52444 63795
rect 52444 63761 52482 63795
rect 52482 63761 52516 63795
rect 52516 63761 52554 63795
rect 52554 63761 52588 63795
rect 52588 63761 52626 63795
rect 52626 63761 52660 63795
rect 52660 63761 52698 63795
rect 52698 63761 52732 63795
rect 52732 63761 52770 63795
rect 52770 63761 52804 63795
rect 52804 63761 52842 63795
rect 52842 63761 52876 63795
rect 52876 63761 52914 63795
rect 52914 63761 52948 63795
rect 52948 63761 52986 63795
rect 52986 63761 53020 63795
rect 53020 63761 53058 63795
rect 53058 63761 53092 63795
rect 53092 63761 53130 63795
rect 53130 63761 53164 63795
rect 53164 63761 53202 63795
rect 53202 63761 53236 63795
rect 53236 63761 53274 63795
rect 53274 63761 53308 63795
rect 53308 63761 53346 63795
rect 53346 63761 53380 63795
rect 53380 63761 53418 63795
rect 53418 63761 53452 63795
rect 53452 63761 53490 63795
rect 53490 63761 53524 63795
rect 53524 63761 53562 63795
rect 53562 63761 53596 63795
rect 53596 63761 53634 63795
rect 53634 63761 53668 63795
rect 53668 63761 53706 63795
rect 53706 63761 53740 63795
rect 53740 63761 53778 63795
rect 53778 63761 53812 63795
rect 53812 63761 53850 63795
rect 53850 63761 53884 63795
rect 53884 63761 53922 63795
rect 53922 63761 53956 63795
rect 53956 63761 53994 63795
rect 53994 63761 54028 63795
rect 54028 63761 54066 63795
rect 54066 63761 54100 63795
rect 54100 63761 54138 63795
rect 54138 63761 54172 63795
rect 54172 63761 54210 63795
rect 54210 63761 54244 63795
rect 54244 63761 54282 63795
rect 54282 63761 54316 63795
rect 54316 63761 54354 63795
rect 54354 63761 54388 63795
rect 54388 63761 54426 63795
rect 54426 63761 54460 63795
rect 54460 63761 54498 63795
rect 54498 63761 54532 63795
rect 54532 63761 54570 63795
rect 54570 63761 54604 63795
rect 54604 63761 54642 63795
rect 54642 63761 54676 63795
rect 54676 63761 54714 63795
rect 54714 63761 54748 63795
rect 54748 63761 54786 63795
rect 54786 63761 54820 63795
rect 54820 63761 54858 63795
rect 54858 63761 54892 63795
rect 54892 63761 54930 63795
rect 54930 63761 54964 63795
rect 54964 63761 55002 63795
rect 55002 63761 55036 63795
rect 55036 63761 55074 63795
rect 55074 63761 55108 63795
rect 55108 63761 55146 63795
rect 55146 63761 55180 63795
rect 55180 63761 55218 63795
rect 55218 63761 55252 63795
rect 55252 63761 55290 63795
rect 55290 63761 55324 63795
rect 55324 63761 55362 63795
rect 55362 63761 55396 63795
rect 55396 63761 55434 63795
rect 55434 63761 55468 63795
rect 55468 63761 55506 63795
rect 55506 63761 55540 63795
rect 55540 63761 55578 63795
rect 55578 63761 55612 63795
rect 55612 63761 55650 63795
rect 55650 63761 55684 63795
rect 55684 63761 55722 63795
rect 55722 63761 55756 63795
rect 55756 63761 55794 63795
rect 55794 63761 55828 63795
rect 55828 63761 55866 63795
rect 55866 63761 55900 63795
rect 55900 63761 55938 63795
rect 55938 63761 55972 63795
rect 55972 63761 56010 63795
rect 56010 63761 56044 63795
rect 56044 63761 56082 63795
rect 56082 63761 56116 63795
rect 56116 63761 56154 63795
rect 56154 63761 56188 63795
rect 56188 63761 56226 63795
rect 56226 63761 56260 63795
rect 56260 63761 56298 63795
rect 56298 63761 56332 63795
rect 56332 63761 56370 63795
rect 56370 63761 56404 63795
rect 56404 63761 56442 63795
rect 56442 63761 56476 63795
rect 56476 63761 56514 63795
rect 56514 63761 56548 63795
rect 56548 63761 56586 63795
rect 56586 63761 56620 63795
rect 56620 63761 56658 63795
rect 56658 63761 56692 63795
rect 56692 63761 56730 63795
rect 56730 63761 56764 63795
rect 56764 63761 56802 63795
rect 56802 63761 56836 63795
rect 56836 63761 56874 63795
rect 56874 63761 56908 63795
rect 56908 63761 56924 63795
rect 51432 63688 56924 63761
rect 57455 69807 57635 69865
rect 57455 69773 57504 69807
rect 57504 69773 57538 69807
rect 57538 69773 57635 69807
rect 57455 69735 57635 69773
rect 57455 69701 57504 69735
rect 57504 69701 57538 69735
rect 57538 69701 57635 69735
rect 57455 69663 57635 69701
rect 57455 69629 57504 69663
rect 57504 69629 57538 69663
rect 57538 69629 57635 69663
rect 57455 69591 57635 69629
rect 57455 69557 57504 69591
rect 57504 69557 57538 69591
rect 57538 69557 57635 69591
rect 57455 69519 57635 69557
rect 57455 69485 57504 69519
rect 57504 69485 57538 69519
rect 57538 69485 57635 69519
rect 57455 69447 57635 69485
rect 57455 69413 57504 69447
rect 57504 69413 57538 69447
rect 57538 69413 57635 69447
rect 57455 69375 57635 69413
rect 57455 69341 57504 69375
rect 57504 69341 57538 69375
rect 57538 69341 57635 69375
rect 57455 69303 57635 69341
rect 57455 69269 57504 69303
rect 57504 69269 57538 69303
rect 57538 69269 57635 69303
rect 57455 69231 57635 69269
rect 57455 69197 57504 69231
rect 57504 69197 57538 69231
rect 57538 69197 57635 69231
rect 57455 69159 57635 69197
rect 57455 69125 57504 69159
rect 57504 69125 57538 69159
rect 57538 69125 57635 69159
rect 57455 69087 57635 69125
rect 57455 69053 57504 69087
rect 57504 69053 57538 69087
rect 57538 69053 57635 69087
rect 57455 69015 57635 69053
rect 57455 68981 57504 69015
rect 57504 68981 57538 69015
rect 57538 68981 57635 69015
rect 57455 68943 57635 68981
rect 57455 68909 57504 68943
rect 57504 68909 57538 68943
rect 57538 68909 57635 68943
rect 57455 68871 57635 68909
rect 57455 68837 57504 68871
rect 57504 68837 57538 68871
rect 57538 68837 57635 68871
rect 57455 68799 57635 68837
rect 57455 68765 57504 68799
rect 57504 68765 57538 68799
rect 57538 68765 57635 68799
rect 57455 68727 57635 68765
rect 57455 68693 57504 68727
rect 57504 68693 57538 68727
rect 57538 68693 57635 68727
rect 57455 68655 57635 68693
rect 57455 68621 57504 68655
rect 57504 68621 57538 68655
rect 57538 68621 57635 68655
rect 57455 68583 57635 68621
rect 57455 68549 57504 68583
rect 57504 68549 57538 68583
rect 57538 68549 57635 68583
rect 57455 68511 57635 68549
rect 57455 68477 57504 68511
rect 57504 68477 57538 68511
rect 57538 68477 57635 68511
rect 57455 68439 57635 68477
rect 57455 68405 57504 68439
rect 57504 68405 57538 68439
rect 57538 68405 57635 68439
rect 57455 68341 57635 68405
rect 57468 65348 57584 65403
rect 57468 65314 57504 65348
rect 57504 65314 57538 65348
rect 57538 65314 57584 65348
rect 57468 65276 57584 65314
rect 57468 65242 57504 65276
rect 57504 65242 57538 65276
rect 57538 65242 57584 65276
rect 57468 65204 57584 65242
rect 57468 65170 57504 65204
rect 57504 65170 57538 65204
rect 57538 65170 57584 65204
rect 57468 65132 57584 65170
rect 57468 65098 57504 65132
rect 57504 65098 57538 65132
rect 57538 65098 57584 65132
rect 57468 65060 57584 65098
rect 57468 65026 57504 65060
rect 57504 65026 57538 65060
rect 57538 65026 57584 65060
rect 57468 64988 57584 65026
rect 57468 64954 57504 64988
rect 57504 64954 57538 64988
rect 57538 64954 57584 64988
rect 57468 64916 57584 64954
rect 57468 64882 57504 64916
rect 57504 64882 57538 64916
rect 57538 64882 57584 64916
rect 57468 64844 57584 64882
rect 57468 64810 57504 64844
rect 57504 64810 57538 64844
rect 57538 64810 57584 64844
rect 57468 64772 57584 64810
rect 57468 64738 57504 64772
rect 57504 64738 57538 64772
rect 57538 64738 57584 64772
rect 57468 64700 57584 64738
rect 57468 64666 57504 64700
rect 57504 64666 57538 64700
rect 57538 64666 57584 64700
rect 57468 64628 57584 64666
rect 57468 64594 57504 64628
rect 57504 64594 57538 64628
rect 57538 64594 57584 64628
rect 57468 64556 57584 64594
rect 57468 64522 57504 64556
rect 57504 64522 57538 64556
rect 57538 64522 57584 64556
rect 57468 64484 57584 64522
rect 57468 64450 57504 64484
rect 57504 64450 57538 64484
rect 57538 64450 57584 64484
rect 57468 64412 57584 64450
rect 57468 64378 57504 64412
rect 57504 64378 57538 64412
rect 57538 64378 57584 64412
rect 57468 64340 57584 64378
rect 57468 64306 57504 64340
rect 57504 64306 57538 64340
rect 57538 64306 57584 64340
rect 57468 64268 57584 64306
rect 57468 64234 57504 64268
rect 57504 64234 57538 64268
rect 57538 64234 57584 64268
rect 57468 64196 57584 64234
rect 57468 64162 57504 64196
rect 57504 64162 57538 64196
rect 57538 64162 57584 64196
rect 57468 64124 57584 64162
rect 57468 64090 57504 64124
rect 57504 64090 57538 64124
rect 57538 64090 57584 64124
rect 57468 63879 57584 64090
rect 59622 62821 59674 62873
rect 59622 62757 59674 62809
rect 59622 62693 59674 62745
rect 57193 62530 57245 62582
rect 58330 62530 58382 62582
rect 59726 62532 59778 62584
rect 62461 62532 62513 62584
rect 59632 62364 59684 62416
rect 59632 62300 59684 62352
rect 59632 62236 59684 62288
rect 59632 62172 59684 62224
rect 59632 62108 59684 62160
rect 62461 62119 62513 62171
rect 59632 62044 59684 62096
rect 57193 61615 57245 61667
rect 60527 61615 60579 61667
rect 59744 61171 59796 61223
rect 59268 61115 59320 61167
rect 59268 61051 59320 61103
rect 59268 60987 59320 61039
rect 59268 60923 59320 60975
rect 57193 60780 57245 60832
rect 57983 60780 58035 60832
rect 59269 60615 59321 60667
rect 59269 60551 59321 60603
rect 59269 60487 59321 60539
rect 59269 60423 59321 60475
rect 59269 60359 59321 60411
rect 59269 60295 59321 60347
rect 60048 60055 60100 60107
rect 60112 60055 60164 60107
rect 60176 60055 60228 60107
rect 60240 60055 60292 60107
rect 60304 60055 60356 60107
rect 60368 60055 60420 60107
rect 67305 63889 67613 70149
rect 74531 88708 74583 88760
rect 74531 88644 74583 88696
rect 74531 88580 74583 88632
rect 74531 88516 74583 88568
rect 74531 88452 74583 88504
rect 74531 88388 74583 88440
rect 74531 88324 74583 88376
rect 74531 88260 74583 88312
rect 74531 88196 74583 88248
rect 81059 88708 81111 88760
rect 81059 88644 81111 88696
rect 81059 88580 81111 88632
rect 81059 88516 81111 88568
rect 81059 88452 81111 88504
rect 81059 88388 81111 88440
rect 81059 88324 81111 88376
rect 81059 88260 81111 88312
rect 81059 88196 81111 88248
rect 88675 88708 88727 88760
rect 88675 88644 88727 88696
rect 88675 88580 88727 88632
rect 88675 88516 88727 88568
rect 88675 88452 88727 88504
rect 88675 88388 88727 88440
rect 88675 88324 88727 88376
rect 88675 88260 88727 88312
rect 88675 88196 88727 88248
rect 75076 86705 75128 86757
rect 75076 86641 75128 86693
rect 75076 86577 75128 86629
rect 75076 86513 75128 86565
rect 75076 86449 75128 86501
rect 75076 86385 75128 86437
rect 75076 86321 75128 86373
rect 75076 86257 75128 86309
rect 75076 86193 75128 86245
rect 76164 86705 76216 86757
rect 76164 86641 76216 86693
rect 76164 86577 76216 86629
rect 76164 86513 76216 86565
rect 76164 86449 76216 86501
rect 76164 86385 76216 86437
rect 76164 86321 76216 86373
rect 76164 86257 76216 86309
rect 76164 86193 76216 86245
rect 78340 86705 78392 86757
rect 78340 86641 78392 86693
rect 78340 86577 78392 86629
rect 78340 86513 78392 86565
rect 78340 86449 78392 86501
rect 78340 86385 78392 86437
rect 78340 86321 78392 86373
rect 78340 86257 78392 86309
rect 78340 86193 78392 86245
rect 79428 86705 79480 86757
rect 79428 86641 79480 86693
rect 79428 86577 79480 86629
rect 79428 86513 79480 86565
rect 79428 86449 79480 86501
rect 79428 86385 79480 86437
rect 79428 86321 79480 86373
rect 79428 86257 79480 86309
rect 79428 86193 79480 86245
rect 80516 86705 80568 86757
rect 80516 86641 80568 86693
rect 80516 86577 80568 86629
rect 80516 86513 80568 86565
rect 80516 86449 80568 86501
rect 80516 86385 80568 86437
rect 80516 86321 80568 86373
rect 80516 86257 80568 86309
rect 80516 86193 80568 86245
rect 81604 86705 81656 86757
rect 81604 86641 81656 86693
rect 81604 86577 81656 86629
rect 81604 86513 81656 86565
rect 81604 86449 81656 86501
rect 81604 86385 81656 86437
rect 81604 86321 81656 86373
rect 81604 86257 81656 86309
rect 81604 86193 81656 86245
rect 82692 86705 82744 86757
rect 82692 86641 82744 86693
rect 82692 86577 82744 86629
rect 82692 86513 82744 86565
rect 82692 86449 82744 86501
rect 82692 86385 82744 86437
rect 82692 86321 82744 86373
rect 82692 86257 82744 86309
rect 82692 86193 82744 86245
rect 83780 86705 83832 86757
rect 83780 86641 83832 86693
rect 83780 86577 83832 86629
rect 83780 86513 83832 86565
rect 83780 86449 83832 86501
rect 83780 86385 83832 86437
rect 83780 86321 83832 86373
rect 83780 86257 83832 86309
rect 83780 86193 83832 86245
rect 85956 86705 86008 86757
rect 85956 86641 86008 86693
rect 85956 86577 86008 86629
rect 85956 86513 86008 86565
rect 85956 86449 86008 86501
rect 85956 86385 86008 86437
rect 85956 86321 86008 86373
rect 85956 86257 86008 86309
rect 85956 86193 86008 86245
rect 87044 86705 87096 86757
rect 87044 86641 87096 86693
rect 87044 86577 87096 86629
rect 87044 86513 87096 86565
rect 87044 86449 87096 86501
rect 87044 86385 87096 86437
rect 87044 86321 87096 86373
rect 87044 86257 87096 86309
rect 87044 86193 87096 86245
rect 88132 86705 88184 86757
rect 88132 86641 88184 86693
rect 88132 86577 88184 86629
rect 88132 86513 88184 86565
rect 88132 86449 88184 86501
rect 88132 86385 88184 86437
rect 88132 86321 88184 86373
rect 88132 86257 88184 86309
rect 88132 86193 88184 86245
rect 74531 84708 74583 84760
rect 74531 84644 74583 84696
rect 74531 84580 74583 84632
rect 74531 84516 74583 84568
rect 74531 84452 74583 84504
rect 74531 84388 74583 84440
rect 74531 84324 74583 84376
rect 74531 84260 74583 84312
rect 74531 84196 74583 84248
rect 75619 84708 75671 84760
rect 75619 84644 75671 84696
rect 75619 84580 75671 84632
rect 75619 84516 75671 84568
rect 75619 84452 75671 84504
rect 75619 84388 75671 84440
rect 75619 84324 75671 84376
rect 75619 84260 75671 84312
rect 75619 84196 75671 84248
rect 76707 84708 76759 84760
rect 76707 84644 76759 84696
rect 76707 84580 76759 84632
rect 76707 84516 76759 84568
rect 76707 84452 76759 84504
rect 76707 84388 76759 84440
rect 76707 84324 76759 84376
rect 76707 84260 76759 84312
rect 76707 84196 76759 84248
rect 77795 84708 77847 84760
rect 77795 84644 77847 84696
rect 77795 84580 77847 84632
rect 77795 84516 77847 84568
rect 77795 84452 77847 84504
rect 77795 84388 77847 84440
rect 77795 84324 77847 84376
rect 77795 84260 77847 84312
rect 77795 84196 77847 84248
rect 78883 84708 78935 84760
rect 78883 84644 78935 84696
rect 78883 84580 78935 84632
rect 78883 84516 78935 84568
rect 78883 84452 78935 84504
rect 78883 84388 78935 84440
rect 78883 84324 78935 84376
rect 78883 84260 78935 84312
rect 78883 84196 78935 84248
rect 79971 84708 80023 84760
rect 79971 84644 80023 84696
rect 79971 84580 80023 84632
rect 79971 84516 80023 84568
rect 79971 84452 80023 84504
rect 79971 84388 80023 84440
rect 79971 84324 80023 84376
rect 79971 84260 80023 84312
rect 79971 84196 80023 84248
rect 81059 84708 81111 84760
rect 81059 84644 81111 84696
rect 81059 84580 81111 84632
rect 81059 84516 81111 84568
rect 81059 84452 81111 84504
rect 81059 84388 81111 84440
rect 81059 84324 81111 84376
rect 81059 84260 81111 84312
rect 81059 84196 81111 84248
rect 82147 84708 82199 84760
rect 82147 84644 82199 84696
rect 82147 84580 82199 84632
rect 82147 84516 82199 84568
rect 82147 84452 82199 84504
rect 82147 84388 82199 84440
rect 82147 84324 82199 84376
rect 82147 84260 82199 84312
rect 82147 84196 82199 84248
rect 83235 84708 83287 84760
rect 83235 84644 83287 84696
rect 83235 84580 83287 84632
rect 83235 84516 83287 84568
rect 83235 84452 83287 84504
rect 83235 84388 83287 84440
rect 83235 84324 83287 84376
rect 83235 84260 83287 84312
rect 83235 84196 83287 84248
rect 84323 84708 84375 84760
rect 84323 84644 84375 84696
rect 84323 84580 84375 84632
rect 84323 84516 84375 84568
rect 84323 84452 84375 84504
rect 84323 84388 84375 84440
rect 84323 84324 84375 84376
rect 84323 84260 84375 84312
rect 84323 84196 84375 84248
rect 85411 84708 85463 84760
rect 85411 84644 85463 84696
rect 85411 84580 85463 84632
rect 85411 84516 85463 84568
rect 85411 84452 85463 84504
rect 85411 84388 85463 84440
rect 85411 84324 85463 84376
rect 85411 84260 85463 84312
rect 85411 84196 85463 84248
rect 86499 84708 86551 84760
rect 86499 84644 86551 84696
rect 86499 84580 86551 84632
rect 86499 84516 86551 84568
rect 86499 84452 86551 84504
rect 86499 84388 86551 84440
rect 86499 84324 86551 84376
rect 86499 84260 86551 84312
rect 86499 84196 86551 84248
rect 87587 84708 87639 84760
rect 87587 84644 87639 84696
rect 87587 84580 87639 84632
rect 87587 84516 87639 84568
rect 87587 84452 87639 84504
rect 87587 84388 87639 84440
rect 87587 84324 87639 84376
rect 87587 84260 87639 84312
rect 87587 84196 87639 84248
rect 88675 84708 88727 84760
rect 88675 84644 88727 84696
rect 88675 84580 88727 84632
rect 88675 84516 88727 84568
rect 88675 84452 88727 84504
rect 88675 84388 88727 84440
rect 88675 84324 88727 84376
rect 88675 84260 88727 84312
rect 88675 84196 88727 84248
rect 75076 82705 75128 82757
rect 75076 82641 75128 82693
rect 75076 82577 75128 82629
rect 75076 82513 75128 82565
rect 75076 82449 75128 82501
rect 75076 82385 75128 82437
rect 75076 82321 75128 82373
rect 75076 82257 75128 82309
rect 75076 82193 75128 82245
rect 76164 82705 76216 82757
rect 76164 82641 76216 82693
rect 76164 82577 76216 82629
rect 76164 82513 76216 82565
rect 76164 82449 76216 82501
rect 76164 82385 76216 82437
rect 76164 82321 76216 82373
rect 76164 82257 76216 82309
rect 76164 82193 76216 82245
rect 77252 82705 77304 82757
rect 77252 82641 77304 82693
rect 77252 82577 77304 82629
rect 77252 82513 77304 82565
rect 77252 82449 77304 82501
rect 77252 82385 77304 82437
rect 77252 82321 77304 82373
rect 77252 82257 77304 82309
rect 77252 82193 77304 82245
rect 78340 82705 78392 82757
rect 78340 82641 78392 82693
rect 78340 82577 78392 82629
rect 78340 82513 78392 82565
rect 78340 82449 78392 82501
rect 78340 82385 78392 82437
rect 78340 82321 78392 82373
rect 78340 82257 78392 82309
rect 78340 82193 78392 82245
rect 79428 82705 79480 82757
rect 79428 82641 79480 82693
rect 79428 82577 79480 82629
rect 79428 82513 79480 82565
rect 79428 82449 79480 82501
rect 79428 82385 79480 82437
rect 79428 82321 79480 82373
rect 79428 82257 79480 82309
rect 79428 82193 79480 82245
rect 80516 82705 80568 82757
rect 80516 82641 80568 82693
rect 80516 82577 80568 82629
rect 80516 82513 80568 82565
rect 80516 82449 80568 82501
rect 80516 82385 80568 82437
rect 80516 82321 80568 82373
rect 80516 82257 80568 82309
rect 80516 82193 80568 82245
rect 81604 82705 81656 82757
rect 81604 82641 81656 82693
rect 81604 82577 81656 82629
rect 81604 82513 81656 82565
rect 81604 82449 81656 82501
rect 81604 82385 81656 82437
rect 81604 82321 81656 82373
rect 81604 82257 81656 82309
rect 81604 82193 81656 82245
rect 82692 82705 82744 82757
rect 82692 82641 82744 82693
rect 82692 82577 82744 82629
rect 82692 82513 82744 82565
rect 82692 82449 82744 82501
rect 82692 82385 82744 82437
rect 82692 82321 82744 82373
rect 82692 82257 82744 82309
rect 82692 82193 82744 82245
rect 83780 82705 83832 82757
rect 83780 82641 83832 82693
rect 83780 82577 83832 82629
rect 83780 82513 83832 82565
rect 83780 82449 83832 82501
rect 83780 82385 83832 82437
rect 83780 82321 83832 82373
rect 83780 82257 83832 82309
rect 83780 82193 83832 82245
rect 84868 82705 84920 82757
rect 84868 82641 84920 82693
rect 84868 82577 84920 82629
rect 84868 82513 84920 82565
rect 84868 82449 84920 82501
rect 84868 82385 84920 82437
rect 84868 82321 84920 82373
rect 84868 82257 84920 82309
rect 84868 82193 84920 82245
rect 85956 82705 86008 82757
rect 85956 82641 86008 82693
rect 85956 82577 86008 82629
rect 85956 82513 86008 82565
rect 85956 82449 86008 82501
rect 85956 82385 86008 82437
rect 85956 82321 86008 82373
rect 85956 82257 86008 82309
rect 85956 82193 86008 82245
rect 87044 82705 87096 82757
rect 87044 82641 87096 82693
rect 87044 82577 87096 82629
rect 87044 82513 87096 82565
rect 87044 82449 87096 82501
rect 87044 82385 87096 82437
rect 87044 82321 87096 82373
rect 87044 82257 87096 82309
rect 87044 82193 87096 82245
rect 88132 82705 88184 82757
rect 88132 82641 88184 82693
rect 88132 82577 88184 82629
rect 88132 82513 88184 82565
rect 88132 82449 88184 82501
rect 88132 82385 88184 82437
rect 88132 82321 88184 82373
rect 88132 82257 88184 82309
rect 88132 82193 88184 82245
rect 74531 80708 74583 80760
rect 74531 80644 74583 80696
rect 74531 80580 74583 80632
rect 74531 80516 74583 80568
rect 74531 80452 74583 80504
rect 74531 80388 74583 80440
rect 74531 80324 74583 80376
rect 74531 80260 74583 80312
rect 74531 80196 74583 80248
rect 75619 80708 75671 80760
rect 75619 80644 75671 80696
rect 75619 80580 75671 80632
rect 75619 80516 75671 80568
rect 75619 80452 75671 80504
rect 75619 80388 75671 80440
rect 75619 80324 75671 80376
rect 75619 80260 75671 80312
rect 75619 80196 75671 80248
rect 76707 80708 76759 80760
rect 76707 80644 76759 80696
rect 76707 80580 76759 80632
rect 76707 80516 76759 80568
rect 76707 80452 76759 80504
rect 76707 80388 76759 80440
rect 76707 80324 76759 80376
rect 76707 80260 76759 80312
rect 76707 80196 76759 80248
rect 77795 80708 77847 80760
rect 77795 80644 77847 80696
rect 77795 80580 77847 80632
rect 77795 80516 77847 80568
rect 77795 80452 77847 80504
rect 77795 80388 77847 80440
rect 77795 80324 77847 80376
rect 77795 80260 77847 80312
rect 77795 80196 77847 80248
rect 78883 80708 78935 80760
rect 78883 80644 78935 80696
rect 78883 80580 78935 80632
rect 78883 80516 78935 80568
rect 78883 80452 78935 80504
rect 78883 80388 78935 80440
rect 78883 80324 78935 80376
rect 78883 80260 78935 80312
rect 78883 80196 78935 80248
rect 79971 80708 80023 80760
rect 79971 80644 80023 80696
rect 79971 80580 80023 80632
rect 79971 80516 80023 80568
rect 79971 80452 80023 80504
rect 79971 80388 80023 80440
rect 79971 80324 80023 80376
rect 79971 80260 80023 80312
rect 79971 80196 80023 80248
rect 81059 80708 81111 80760
rect 81059 80644 81111 80696
rect 81059 80580 81111 80632
rect 81059 80516 81111 80568
rect 81059 80452 81111 80504
rect 81059 80388 81111 80440
rect 81059 80324 81111 80376
rect 81059 80260 81111 80312
rect 81059 80196 81111 80248
rect 82147 80708 82199 80760
rect 82147 80644 82199 80696
rect 82147 80580 82199 80632
rect 82147 80516 82199 80568
rect 82147 80452 82199 80504
rect 82147 80388 82199 80440
rect 82147 80324 82199 80376
rect 82147 80260 82199 80312
rect 82147 80196 82199 80248
rect 83235 80708 83287 80760
rect 83235 80644 83287 80696
rect 83235 80580 83287 80632
rect 83235 80516 83287 80568
rect 83235 80452 83287 80504
rect 83235 80388 83287 80440
rect 83235 80324 83287 80376
rect 83235 80260 83287 80312
rect 83235 80196 83287 80248
rect 84323 80708 84375 80760
rect 84323 80644 84375 80696
rect 84323 80580 84375 80632
rect 84323 80516 84375 80568
rect 84323 80452 84375 80504
rect 84323 80388 84375 80440
rect 84323 80324 84375 80376
rect 84323 80260 84375 80312
rect 84323 80196 84375 80248
rect 85411 80708 85463 80760
rect 85411 80644 85463 80696
rect 85411 80580 85463 80632
rect 85411 80516 85463 80568
rect 85411 80452 85463 80504
rect 85411 80388 85463 80440
rect 85411 80324 85463 80376
rect 85411 80260 85463 80312
rect 85411 80196 85463 80248
rect 86499 80708 86551 80760
rect 86499 80644 86551 80696
rect 86499 80580 86551 80632
rect 86499 80516 86551 80568
rect 86499 80452 86551 80504
rect 86499 80388 86551 80440
rect 86499 80324 86551 80376
rect 86499 80260 86551 80312
rect 86499 80196 86551 80248
rect 87587 80708 87639 80760
rect 87587 80644 87639 80696
rect 87587 80580 87639 80632
rect 87587 80516 87639 80568
rect 87587 80452 87639 80504
rect 87587 80388 87639 80440
rect 87587 80324 87639 80376
rect 87587 80260 87639 80312
rect 87587 80196 87639 80248
rect 88675 80708 88727 80760
rect 88675 80644 88727 80696
rect 88675 80580 88727 80632
rect 88675 80516 88727 80568
rect 88675 80452 88727 80504
rect 88675 80388 88727 80440
rect 88675 80324 88727 80376
rect 88675 80260 88727 80312
rect 88675 80196 88727 80248
rect 75076 78705 75128 78757
rect 75076 78641 75128 78693
rect 75076 78577 75128 78629
rect 75076 78513 75128 78565
rect 75076 78449 75128 78501
rect 75076 78385 75128 78437
rect 75076 78321 75128 78373
rect 75076 78257 75128 78309
rect 75076 78193 75128 78245
rect 76164 78705 76216 78757
rect 76164 78641 76216 78693
rect 76164 78577 76216 78629
rect 76164 78513 76216 78565
rect 76164 78449 76216 78501
rect 76164 78385 76216 78437
rect 76164 78321 76216 78373
rect 76164 78257 76216 78309
rect 76164 78193 76216 78245
rect 77252 78705 77304 78757
rect 77252 78641 77304 78693
rect 77252 78577 77304 78629
rect 77252 78513 77304 78565
rect 77252 78449 77304 78501
rect 77252 78385 77304 78437
rect 77252 78321 77304 78373
rect 77252 78257 77304 78309
rect 77252 78193 77304 78245
rect 78340 78705 78392 78757
rect 78340 78641 78392 78693
rect 78340 78577 78392 78629
rect 78340 78513 78392 78565
rect 78340 78449 78392 78501
rect 78340 78385 78392 78437
rect 78340 78321 78392 78373
rect 78340 78257 78392 78309
rect 78340 78193 78392 78245
rect 79428 78705 79480 78757
rect 79428 78641 79480 78693
rect 79428 78577 79480 78629
rect 79428 78513 79480 78565
rect 79428 78449 79480 78501
rect 79428 78385 79480 78437
rect 79428 78321 79480 78373
rect 79428 78257 79480 78309
rect 79428 78193 79480 78245
rect 80516 78705 80568 78757
rect 80516 78641 80568 78693
rect 80516 78577 80568 78629
rect 80516 78513 80568 78565
rect 80516 78449 80568 78501
rect 80516 78385 80568 78437
rect 80516 78321 80568 78373
rect 80516 78257 80568 78309
rect 80516 78193 80568 78245
rect 81604 78705 81656 78757
rect 81604 78641 81656 78693
rect 81604 78577 81656 78629
rect 81604 78513 81656 78565
rect 81604 78449 81656 78501
rect 81604 78385 81656 78437
rect 81604 78321 81656 78373
rect 81604 78257 81656 78309
rect 81604 78193 81656 78245
rect 82692 78705 82744 78757
rect 82692 78641 82744 78693
rect 82692 78577 82744 78629
rect 82692 78513 82744 78565
rect 82692 78449 82744 78501
rect 82692 78385 82744 78437
rect 82692 78321 82744 78373
rect 82692 78257 82744 78309
rect 82692 78193 82744 78245
rect 83780 78705 83832 78757
rect 83780 78641 83832 78693
rect 83780 78577 83832 78629
rect 83780 78513 83832 78565
rect 83780 78449 83832 78501
rect 83780 78385 83832 78437
rect 83780 78321 83832 78373
rect 83780 78257 83832 78309
rect 83780 78193 83832 78245
rect 84868 78705 84920 78757
rect 84868 78641 84920 78693
rect 84868 78577 84920 78629
rect 84868 78513 84920 78565
rect 84868 78449 84920 78501
rect 84868 78385 84920 78437
rect 84868 78321 84920 78373
rect 84868 78257 84920 78309
rect 84868 78193 84920 78245
rect 85956 78705 86008 78757
rect 85956 78641 86008 78693
rect 85956 78577 86008 78629
rect 85956 78513 86008 78565
rect 85956 78449 86008 78501
rect 85956 78385 86008 78437
rect 85956 78321 86008 78373
rect 85956 78257 86008 78309
rect 85956 78193 86008 78245
rect 87044 78705 87096 78757
rect 87044 78641 87096 78693
rect 87044 78577 87096 78629
rect 87044 78513 87096 78565
rect 87044 78449 87096 78501
rect 87044 78385 87096 78437
rect 87044 78321 87096 78373
rect 87044 78257 87096 78309
rect 87044 78193 87096 78245
rect 88132 78705 88184 78757
rect 88132 78641 88184 78693
rect 88132 78577 88184 78629
rect 88132 78513 88184 78565
rect 88132 78449 88184 78501
rect 88132 78385 88184 78437
rect 88132 78321 88184 78373
rect 88132 78257 88184 78309
rect 88132 78193 88184 78245
rect 74531 76708 74583 76760
rect 74531 76644 74583 76696
rect 74531 76580 74583 76632
rect 74531 76516 74583 76568
rect 74531 76452 74583 76504
rect 74531 76388 74583 76440
rect 74531 76324 74583 76376
rect 74531 76260 74583 76312
rect 74531 76196 74583 76248
rect 75619 76708 75671 76760
rect 75619 76644 75671 76696
rect 75619 76580 75671 76632
rect 75619 76516 75671 76568
rect 75619 76452 75671 76504
rect 75619 76388 75671 76440
rect 75619 76324 75671 76376
rect 75619 76260 75671 76312
rect 75619 76196 75671 76248
rect 76707 76708 76759 76760
rect 76707 76644 76759 76696
rect 76707 76580 76759 76632
rect 76707 76516 76759 76568
rect 76707 76452 76759 76504
rect 76707 76388 76759 76440
rect 76707 76324 76759 76376
rect 76707 76260 76759 76312
rect 76707 76196 76759 76248
rect 77795 76708 77847 76760
rect 77795 76644 77847 76696
rect 77795 76580 77847 76632
rect 77795 76516 77847 76568
rect 77795 76452 77847 76504
rect 77795 76388 77847 76440
rect 77795 76324 77847 76376
rect 77795 76260 77847 76312
rect 77795 76196 77847 76248
rect 78883 76708 78935 76760
rect 78883 76644 78935 76696
rect 78883 76580 78935 76632
rect 78883 76516 78935 76568
rect 78883 76452 78935 76504
rect 78883 76388 78935 76440
rect 78883 76324 78935 76376
rect 78883 76260 78935 76312
rect 78883 76196 78935 76248
rect 79971 76708 80023 76760
rect 79971 76644 80023 76696
rect 79971 76580 80023 76632
rect 79971 76516 80023 76568
rect 79971 76452 80023 76504
rect 79971 76388 80023 76440
rect 79971 76324 80023 76376
rect 79971 76260 80023 76312
rect 79971 76196 80023 76248
rect 81059 76708 81111 76760
rect 81059 76644 81111 76696
rect 81059 76580 81111 76632
rect 81059 76516 81111 76568
rect 81059 76452 81111 76504
rect 81059 76388 81111 76440
rect 81059 76324 81111 76376
rect 81059 76260 81111 76312
rect 81059 76196 81111 76248
rect 82147 76708 82199 76760
rect 82147 76644 82199 76696
rect 82147 76580 82199 76632
rect 82147 76516 82199 76568
rect 82147 76452 82199 76504
rect 82147 76388 82199 76440
rect 82147 76324 82199 76376
rect 82147 76260 82199 76312
rect 82147 76196 82199 76248
rect 83235 76708 83287 76760
rect 83235 76644 83287 76696
rect 83235 76580 83287 76632
rect 83235 76516 83287 76568
rect 83235 76452 83287 76504
rect 83235 76388 83287 76440
rect 83235 76324 83287 76376
rect 83235 76260 83287 76312
rect 83235 76196 83287 76248
rect 84323 76708 84375 76760
rect 84323 76644 84375 76696
rect 84323 76580 84375 76632
rect 84323 76516 84375 76568
rect 84323 76452 84375 76504
rect 84323 76388 84375 76440
rect 84323 76324 84375 76376
rect 84323 76260 84375 76312
rect 84323 76196 84375 76248
rect 85411 76708 85463 76760
rect 85411 76644 85463 76696
rect 85411 76580 85463 76632
rect 85411 76516 85463 76568
rect 85411 76452 85463 76504
rect 85411 76388 85463 76440
rect 85411 76324 85463 76376
rect 85411 76260 85463 76312
rect 85411 76196 85463 76248
rect 86499 76708 86551 76760
rect 86499 76644 86551 76696
rect 86499 76580 86551 76632
rect 86499 76516 86551 76568
rect 86499 76452 86551 76504
rect 86499 76388 86551 76440
rect 86499 76324 86551 76376
rect 86499 76260 86551 76312
rect 86499 76196 86551 76248
rect 87587 76708 87639 76760
rect 87587 76644 87639 76696
rect 87587 76580 87639 76632
rect 87587 76516 87639 76568
rect 87587 76452 87639 76504
rect 87587 76388 87639 76440
rect 87587 76324 87639 76376
rect 87587 76260 87639 76312
rect 87587 76196 87639 76248
rect 88675 76708 88727 76760
rect 88675 76644 88727 76696
rect 88675 76580 88727 76632
rect 88675 76516 88727 76568
rect 88675 76452 88727 76504
rect 88675 76388 88727 76440
rect 88675 76324 88727 76376
rect 88675 76260 88727 76312
rect 88675 76196 88727 76248
rect 75076 74705 75128 74757
rect 75076 74641 75128 74693
rect 75076 74577 75128 74629
rect 75076 74513 75128 74565
rect 75076 74449 75128 74501
rect 75076 74385 75128 74437
rect 75076 74321 75128 74373
rect 75076 74257 75128 74309
rect 75076 74193 75128 74245
rect 77252 74705 77304 74757
rect 77252 74641 77304 74693
rect 77252 74577 77304 74629
rect 77252 74513 77304 74565
rect 77252 74449 77304 74501
rect 77252 74385 77304 74437
rect 77252 74321 77304 74373
rect 77252 74257 77304 74309
rect 77252 74193 77304 74245
rect 78340 74705 78392 74757
rect 78340 74641 78392 74693
rect 78340 74577 78392 74629
rect 78340 74513 78392 74565
rect 78340 74449 78392 74501
rect 78340 74385 78392 74437
rect 78340 74321 78392 74373
rect 78340 74257 78392 74309
rect 78340 74193 78392 74245
rect 80516 74705 80568 74757
rect 80516 74641 80568 74693
rect 80516 74577 80568 74629
rect 80516 74513 80568 74565
rect 80516 74449 80568 74501
rect 80516 74385 80568 74437
rect 80516 74321 80568 74373
rect 80516 74257 80568 74309
rect 80516 74193 80568 74245
rect 81604 74705 81656 74757
rect 81604 74641 81656 74693
rect 81604 74577 81656 74629
rect 81604 74513 81656 74565
rect 81604 74449 81656 74501
rect 81604 74385 81656 74437
rect 81604 74321 81656 74373
rect 81604 74257 81656 74309
rect 81604 74193 81656 74245
rect 82692 74705 82744 74757
rect 82692 74641 82744 74693
rect 82692 74577 82744 74629
rect 82692 74513 82744 74565
rect 82692 74449 82744 74501
rect 82692 74385 82744 74437
rect 82692 74321 82744 74373
rect 82692 74257 82744 74309
rect 82692 74193 82744 74245
rect 84868 74705 84920 74757
rect 84868 74641 84920 74693
rect 84868 74577 84920 74629
rect 84868 74513 84920 74565
rect 84868 74449 84920 74501
rect 84868 74385 84920 74437
rect 84868 74321 84920 74373
rect 84868 74257 84920 74309
rect 84868 74193 84920 74245
rect 85956 74705 86008 74757
rect 85956 74641 86008 74693
rect 85956 74577 86008 74629
rect 85956 74513 86008 74565
rect 85956 74449 86008 74501
rect 85956 74385 86008 74437
rect 85956 74321 86008 74373
rect 85956 74257 86008 74309
rect 85956 74193 86008 74245
rect 88132 74705 88184 74757
rect 88132 74641 88184 74693
rect 88132 74577 88184 74629
rect 88132 74513 88184 74565
rect 88132 74449 88184 74501
rect 88132 74385 88184 74437
rect 88132 74321 88184 74373
rect 88132 74257 88184 74309
rect 88132 74193 88184 74245
rect 74531 72708 74583 72760
rect 74531 72644 74583 72696
rect 74531 72580 74583 72632
rect 74531 72516 74583 72568
rect 74531 72452 74583 72504
rect 74531 72388 74583 72440
rect 74531 72324 74583 72376
rect 74531 72260 74583 72312
rect 74531 72196 74583 72248
rect 75619 72708 75671 72760
rect 75619 72644 75671 72696
rect 75619 72580 75671 72632
rect 75619 72516 75671 72568
rect 75619 72452 75671 72504
rect 75619 72388 75671 72440
rect 75619 72324 75671 72376
rect 75619 72260 75671 72312
rect 75619 72196 75671 72248
rect 76707 72708 76759 72760
rect 76707 72644 76759 72696
rect 76707 72580 76759 72632
rect 76707 72516 76759 72568
rect 76707 72452 76759 72504
rect 76707 72388 76759 72440
rect 76707 72324 76759 72376
rect 76707 72260 76759 72312
rect 76707 72196 76759 72248
rect 77795 72708 77847 72760
rect 77795 72644 77847 72696
rect 77795 72580 77847 72632
rect 77795 72516 77847 72568
rect 77795 72452 77847 72504
rect 77795 72388 77847 72440
rect 77795 72324 77847 72376
rect 77795 72260 77847 72312
rect 77795 72196 77847 72248
rect 78883 72708 78935 72760
rect 78883 72644 78935 72696
rect 78883 72580 78935 72632
rect 78883 72516 78935 72568
rect 78883 72452 78935 72504
rect 78883 72388 78935 72440
rect 78883 72324 78935 72376
rect 78883 72260 78935 72312
rect 78883 72196 78935 72248
rect 79971 72708 80023 72760
rect 79971 72644 80023 72696
rect 79971 72580 80023 72632
rect 79971 72516 80023 72568
rect 79971 72452 80023 72504
rect 79971 72388 80023 72440
rect 79971 72324 80023 72376
rect 79971 72260 80023 72312
rect 79971 72196 80023 72248
rect 81059 72708 81111 72760
rect 81059 72644 81111 72696
rect 81059 72580 81111 72632
rect 81059 72516 81111 72568
rect 81059 72452 81111 72504
rect 81059 72388 81111 72440
rect 81059 72324 81111 72376
rect 81059 72260 81111 72312
rect 81059 72196 81111 72248
rect 86499 72708 86551 72760
rect 86499 72644 86551 72696
rect 86499 72580 86551 72632
rect 86499 72516 86551 72568
rect 86499 72452 86551 72504
rect 86499 72388 86551 72440
rect 86499 72324 86551 72376
rect 86499 72260 86551 72312
rect 86499 72196 86551 72248
rect 87587 72708 87639 72760
rect 87587 72644 87639 72696
rect 87587 72580 87639 72632
rect 87587 72516 87639 72568
rect 87587 72452 87639 72504
rect 87587 72388 87639 72440
rect 87587 72324 87639 72376
rect 87587 72260 87639 72312
rect 87587 72196 87639 72248
rect 88675 72708 88727 72760
rect 88675 72644 88727 72696
rect 88675 72580 88727 72632
rect 88675 72516 88727 72568
rect 88675 72452 88727 72504
rect 88675 72388 88727 72440
rect 88675 72324 88727 72376
rect 88675 72260 88727 72312
rect 88675 72196 88727 72248
rect 75076 70705 75128 70757
rect 75076 70641 75128 70693
rect 75076 70577 75128 70629
rect 75076 70513 75128 70565
rect 75076 70449 75128 70501
rect 75076 70385 75128 70437
rect 75076 70321 75128 70373
rect 75076 70257 75128 70309
rect 75076 70193 75128 70245
rect 76164 70705 76216 70757
rect 76164 70641 76216 70693
rect 76164 70577 76216 70629
rect 76164 70513 76216 70565
rect 76164 70449 76216 70501
rect 76164 70385 76216 70437
rect 76164 70321 76216 70373
rect 76164 70257 76216 70309
rect 76164 70193 76216 70245
rect 77252 70705 77304 70757
rect 77252 70641 77304 70693
rect 77252 70577 77304 70629
rect 77252 70513 77304 70565
rect 77252 70449 77304 70501
rect 77252 70385 77304 70437
rect 77252 70321 77304 70373
rect 77252 70257 77304 70309
rect 77252 70193 77304 70245
rect 78340 70705 78392 70757
rect 78340 70641 78392 70693
rect 78340 70577 78392 70629
rect 78340 70513 78392 70565
rect 78340 70449 78392 70501
rect 78340 70385 78392 70437
rect 78340 70321 78392 70373
rect 78340 70257 78392 70309
rect 78340 70193 78392 70245
rect 79428 70705 79480 70757
rect 79428 70641 79480 70693
rect 79428 70577 79480 70629
rect 79428 70513 79480 70565
rect 79428 70449 79480 70501
rect 79428 70385 79480 70437
rect 79428 70321 79480 70373
rect 79428 70257 79480 70309
rect 79428 70193 79480 70245
rect 81604 70705 81656 70757
rect 81604 70641 81656 70693
rect 81604 70577 81656 70629
rect 81604 70513 81656 70565
rect 81604 70449 81656 70501
rect 81604 70385 81656 70437
rect 81604 70321 81656 70373
rect 81604 70257 81656 70309
rect 81604 70193 81656 70245
rect 82692 70705 82744 70757
rect 82692 70641 82744 70693
rect 82692 70577 82744 70629
rect 82692 70513 82744 70565
rect 82692 70449 82744 70501
rect 82692 70385 82744 70437
rect 82692 70321 82744 70373
rect 82692 70257 82744 70309
rect 82692 70193 82744 70245
rect 83780 70705 83832 70757
rect 83780 70641 83832 70693
rect 83780 70577 83832 70629
rect 83780 70513 83832 70565
rect 83780 70449 83832 70501
rect 83780 70385 83832 70437
rect 83780 70321 83832 70373
rect 83780 70257 83832 70309
rect 83780 70193 83832 70245
rect 84868 70705 84920 70757
rect 84868 70641 84920 70693
rect 84868 70577 84920 70629
rect 84868 70513 84920 70565
rect 84868 70449 84920 70501
rect 84868 70385 84920 70437
rect 84868 70321 84920 70373
rect 84868 70257 84920 70309
rect 84868 70193 84920 70245
rect 85956 70705 86008 70757
rect 85956 70641 86008 70693
rect 85956 70577 86008 70629
rect 85956 70513 86008 70565
rect 85956 70449 86008 70501
rect 85956 70385 86008 70437
rect 85956 70321 86008 70373
rect 85956 70257 86008 70309
rect 85956 70193 86008 70245
rect 87044 70705 87096 70757
rect 87044 70641 87096 70693
rect 87044 70577 87096 70629
rect 87044 70513 87096 70565
rect 87044 70449 87096 70501
rect 87044 70385 87096 70437
rect 87044 70321 87096 70373
rect 87044 70257 87096 70309
rect 87044 70193 87096 70245
rect 88132 70705 88184 70757
rect 88132 70641 88184 70693
rect 88132 70577 88184 70629
rect 88132 70513 88184 70565
rect 88132 70449 88184 70501
rect 88132 70385 88184 70437
rect 88132 70321 88184 70373
rect 88132 70257 88184 70309
rect 88132 70193 88184 70245
rect 75345 69712 75397 69764
rect 75891 69712 75943 69764
rect 76437 69703 76489 69755
rect 76982 69702 77034 69754
rect 78613 69690 78665 69742
rect 79156 69687 79208 69739
rect 79698 69686 79750 69738
rect 80245 69691 80297 69743
rect 82963 69702 83015 69754
rect 83506 69706 83558 69758
rect 84048 69700 84100 69752
rect 84605 69691 84657 69743
rect 86229 69702 86281 69754
rect 86773 69695 86825 69747
rect 87323 69699 87375 69751
rect 87856 69699 87908 69751
rect 101874 69036 101926 69088
rect 101938 69036 101990 69088
rect 102002 69036 102054 69088
rect 102066 69036 102118 69088
rect 102130 69036 102182 69088
rect 102194 69036 102246 69088
rect 102258 69036 102310 69088
rect 102322 69036 102374 69088
rect 96657 68855 96709 68907
rect 97689 68838 97741 68852
rect 97689 68804 97697 68838
rect 97697 68804 97731 68838
rect 97731 68804 97741 68838
rect 97689 68800 97741 68804
rect 98089 68832 98141 68841
rect 98089 68798 98099 68832
rect 98099 68798 98133 68832
rect 98133 68798 98141 68832
rect 98089 68789 98141 68798
rect 98246 68838 98298 68845
rect 98246 68804 98255 68838
rect 98255 68804 98289 68838
rect 98289 68804 98298 68838
rect 98246 68793 98298 68804
rect 97988 68773 98040 68784
rect 97988 68739 97999 68773
rect 97999 68739 98033 68773
rect 98033 68739 98040 68773
rect 97988 68732 98040 68739
rect 96657 68665 96709 68717
rect 103416 68753 103596 68933
rect 98635 68490 98687 68542
rect 98699 68490 98751 68542
rect 98763 68490 98815 68542
rect 98827 68490 98879 68542
rect 98891 68490 98943 68542
rect 101873 67885 101925 67937
rect 101937 67885 101989 67937
rect 102001 67885 102053 67937
rect 102065 67885 102117 67937
rect 102129 67885 102181 67937
rect 102193 67885 102245 67937
rect 102257 67885 102309 67937
rect 102321 67885 102373 67937
rect 96657 67705 96709 67757
rect 97689 67688 97741 67702
rect 97689 67654 97697 67688
rect 97697 67654 97731 67688
rect 97731 67654 97741 67688
rect 97689 67650 97741 67654
rect 98089 67682 98141 67691
rect 98089 67648 98099 67682
rect 98099 67648 98133 67682
rect 98133 67648 98141 67682
rect 98089 67639 98141 67648
rect 98246 67688 98298 67695
rect 98246 67654 98255 67688
rect 98255 67654 98289 67688
rect 98289 67654 98298 67688
rect 98246 67643 98298 67654
rect 97988 67623 98040 67634
rect 97988 67589 97999 67623
rect 97999 67589 98033 67623
rect 98033 67589 98040 67623
rect 97988 67582 98040 67589
rect 96657 67515 96709 67567
rect 103404 67602 103584 67782
rect 98633 67340 98685 67392
rect 98697 67340 98749 67392
rect 98761 67340 98813 67392
rect 98825 67340 98877 67392
rect 98889 67340 98941 67392
rect 101863 65343 101915 65395
rect 101927 65343 101979 65395
rect 101991 65343 102043 65395
rect 102055 65343 102107 65395
rect 102119 65343 102171 65395
rect 102183 65343 102235 65395
rect 102247 65343 102299 65395
rect 102311 65343 102363 65395
rect 96657 65165 96709 65217
rect 97689 65148 97741 65162
rect 97689 65114 97697 65148
rect 97697 65114 97731 65148
rect 97731 65114 97741 65148
rect 97689 65110 97741 65114
rect 98089 65142 98141 65151
rect 98089 65108 98099 65142
rect 98099 65108 98133 65142
rect 98133 65108 98141 65142
rect 98089 65099 98141 65108
rect 98246 65148 98298 65155
rect 98246 65114 98255 65148
rect 98255 65114 98289 65148
rect 98289 65114 98298 65148
rect 98246 65103 98298 65114
rect 97988 65083 98040 65094
rect 97988 65049 97999 65083
rect 97999 65049 98033 65083
rect 98033 65049 98040 65083
rect 97988 65042 98040 65049
rect 96657 64975 96709 65027
rect 103262 65070 103442 65250
rect 98551 64799 98603 64851
rect 98615 64799 98667 64851
rect 98679 64799 98731 64851
rect 98743 64799 98795 64851
rect 98807 64799 98859 64851
rect 101863 64073 101915 64125
rect 101927 64073 101979 64125
rect 101991 64073 102043 64125
rect 102055 64073 102107 64125
rect 102119 64073 102171 64125
rect 102183 64073 102235 64125
rect 102247 64073 102299 64125
rect 102311 64073 102363 64125
rect 96657 63895 96709 63947
rect 97689 63878 97741 63892
rect 97689 63844 97697 63878
rect 97697 63844 97731 63878
rect 97731 63844 97741 63878
rect 97689 63840 97741 63844
rect 98089 63872 98141 63881
rect 98089 63838 98099 63872
rect 98099 63838 98133 63872
rect 98133 63838 98141 63872
rect 98089 63829 98141 63838
rect 98246 63878 98298 63885
rect 98246 63844 98255 63878
rect 98255 63844 98289 63878
rect 98289 63844 98298 63878
rect 98246 63833 98298 63844
rect 97988 63813 98040 63824
rect 97988 63779 97999 63813
rect 97999 63779 98033 63813
rect 98033 63779 98040 63813
rect 97988 63772 98040 63779
rect 96657 63705 96709 63757
rect 103233 63780 103413 63960
rect 98549 63530 98601 63582
rect 98613 63530 98665 63582
rect 98677 63530 98729 63582
rect 98741 63530 98793 63582
rect 98805 63530 98857 63582
rect 64204 63024 64384 63204
rect 69664 63024 69844 63204
rect 64336 62119 64388 62171
rect 62529 61171 62581 61223
rect 63801 61171 63853 61223
rect 60700 60058 60752 60110
rect 60764 60058 60816 60110
rect 60828 60058 60880 60110
rect 62175 60057 62227 60109
rect 62239 60057 62291 60109
rect 62303 60057 62355 60109
rect 62367 60057 62419 60109
rect 66528 61615 66580 61667
rect 62691 60058 62743 60110
rect 62755 60058 62807 60110
rect 62819 60058 62871 60110
rect 64050 60050 64102 60102
rect 64114 60050 64166 60102
rect 64178 60050 64230 60102
rect 64504 60057 64556 60109
rect 64568 60057 64620 60109
rect 64632 60057 64684 60109
rect 64696 60057 64748 60109
rect 66042 60056 66094 60108
rect 66106 60056 66158 60108
rect 66170 60056 66222 60108
rect 66234 60056 66286 60108
rect 66298 60056 66350 60108
rect 66362 60056 66414 60108
rect 66692 60053 66744 60105
rect 66756 60053 66808 60105
rect 66820 60053 66872 60105
rect 62530 58984 62582 59036
rect 64342 58982 64394 59034
rect 60839 57820 60891 57872
rect 50152 57143 50204 57195
rect 50111 55775 50163 55827
rect 50175 55775 50227 55827
rect 62530 58389 62582 58441
rect 64342 58389 64394 58441
rect 62530 57525 62582 57577
rect 64528 57533 64580 57585
rect 66839 57820 66891 57872
rect 61454 54396 61506 54448
rect 65428 54401 65480 54453
rect 47703 54269 47755 54321
rect 47767 54269 47819 54321
rect 44407 53716 44459 53768
rect 26901 53187 27017 53303
rect 38577 53187 38693 53303
rect 43631 53293 43683 53345
rect 59051 52772 59103 52824
rect 59115 52772 59167 52824
rect 65060 52810 65112 52862
rect 51014 52572 51066 52624
rect 51078 52572 51130 52624
rect 60499 52559 60551 52611
rect 41405 52059 41457 52111
rect 41405 51995 41457 52047
rect 43111 52036 43163 52088
rect 26070 51829 26186 51945
rect 37717 51829 37833 51945
rect 41405 51931 41457 51983
rect 41405 51867 41457 51919
rect 41405 51803 41457 51855
rect 41405 51739 41457 51791
rect 41405 51675 41457 51727
rect 44715 52029 44767 52081
rect 44715 51965 44767 52017
rect 44715 51901 44767 51953
rect 44715 51837 44767 51889
rect 44715 51773 44767 51825
rect 44715 51709 44767 51761
rect 38774 51539 38826 51591
rect 39465 51544 39581 51660
rect 42188 51541 42240 51593
rect 44722 51372 44774 51424
rect 44722 51308 44774 51360
rect 42690 51229 42742 51281
rect 44722 51244 44774 51296
rect 38774 51062 38826 51114
rect 38219 50724 38271 50776
rect 18913 50558 18965 50610
rect 18977 50558 19029 50610
rect 19041 50558 19093 50610
rect 19105 50558 19157 50610
rect 19169 50558 19221 50610
rect 19233 50558 19285 50610
rect 19297 50558 19349 50610
rect 19361 50558 19413 50610
rect 19425 50558 19477 50610
rect 19489 50558 19541 50610
rect 19553 50558 19605 50610
rect 19617 50558 19669 50610
rect 19681 50558 19733 50610
rect 19745 50558 19797 50610
rect 19809 50558 19861 50610
rect 19873 50558 19925 50610
rect 19937 50558 19989 50610
rect 20001 50558 20053 50610
rect 20065 50558 20117 50610
rect 20129 50558 20181 50610
rect 20193 50558 20245 50610
rect 20257 50558 20309 50610
rect 20321 50558 20373 50610
rect 20385 50558 20437 50610
rect 20449 50558 20501 50610
rect 20513 50558 20565 50610
rect 20577 50558 20629 50610
rect 20641 50558 20693 50610
rect 20705 50558 20757 50610
rect 20769 50558 20821 50610
rect 20833 50558 20885 50610
rect 20897 50558 20949 50610
rect 20961 50558 21013 50610
rect 21025 50558 21077 50610
rect 21089 50558 21141 50610
rect 21153 50558 21205 50610
rect 21217 50558 21269 50610
rect 21281 50558 21333 50610
rect 21345 50558 21397 50610
rect 21409 50558 21461 50610
rect 21473 50558 21525 50610
rect 21537 50558 21589 50610
rect 21601 50558 21653 50610
rect 21665 50558 21717 50610
rect 21729 50558 21781 50610
rect 21793 50558 21845 50610
rect 21857 50558 21909 50610
rect 21921 50558 21973 50610
rect 21985 50558 22037 50610
rect 22049 50558 22101 50610
rect 22113 50558 22165 50610
rect 22177 50558 22229 50610
rect 38218 49941 38270 49993
rect 31659 49420 31711 49472
rect 31659 49356 31711 49408
rect 31659 49292 31711 49344
rect 31659 49228 31711 49280
rect 16529 48985 16709 49165
rect 24109 49012 24225 49128
rect 31659 48889 31711 48941
rect 31659 48825 31711 48877
rect 31659 48761 31711 48813
rect 18919 47550 18971 47602
rect 18983 47550 19035 47602
rect 19047 47550 19099 47602
rect 19111 47550 19163 47602
rect 19175 47550 19227 47602
rect 19239 47550 19291 47602
rect 19303 47550 19355 47602
rect 19367 47550 19419 47602
rect 19431 47550 19483 47602
rect 19495 47550 19547 47602
rect 19559 47550 19611 47602
rect 19623 47550 19675 47602
rect 19687 47550 19739 47602
rect 19751 47550 19803 47602
rect 19815 47550 19867 47602
rect 19879 47550 19931 47602
rect 19943 47550 19995 47602
rect 20007 47550 20059 47602
rect 20071 47550 20123 47602
rect 20135 47550 20187 47602
rect 20199 47550 20251 47602
rect 20263 47550 20315 47602
rect 20327 47550 20379 47602
rect 20391 47550 20443 47602
rect 20455 47550 20507 47602
rect 20519 47550 20571 47602
rect 20583 47550 20635 47602
rect 20647 47550 20699 47602
rect 20711 47550 20763 47602
rect 20775 47550 20827 47602
rect 20839 47550 20891 47602
rect 20903 47550 20955 47602
rect 20967 47550 21019 47602
rect 21031 47550 21083 47602
rect 21095 47550 21147 47602
rect 21159 47550 21211 47602
rect 21223 47550 21275 47602
rect 21287 47550 21339 47602
rect 21351 47550 21403 47602
rect 21415 47550 21467 47602
rect 21479 47550 21531 47602
rect 21543 47550 21595 47602
rect 21607 47550 21659 47602
rect 21671 47550 21723 47602
rect 21735 47550 21787 47602
rect 21799 47550 21851 47602
rect 21863 47550 21915 47602
rect 21927 47550 21979 47602
rect 21991 47550 22043 47602
rect 22055 47550 22107 47602
rect 22119 47550 22171 47602
rect 22183 47550 22235 47602
rect 42188 51053 42240 51105
rect 39844 50724 39896 50776
rect 47084 50552 47136 50604
rect 47148 50552 47200 50604
rect 43111 50436 43163 50488
rect 39465 50315 39581 50431
rect 44719 50427 44771 50479
rect 44719 50363 44771 50415
rect 41387 50222 41439 50274
rect 41387 50158 41439 50210
rect 41387 50094 41439 50146
rect 44719 50299 44771 50351
rect 44719 50235 44771 50287
rect 44719 50171 44771 50223
rect 44719 50107 44771 50159
rect 42188 49937 42240 49989
rect 44715 49773 44767 49825
rect 59052 49784 59104 49836
rect 59116 49784 59168 49836
rect 44715 49709 44767 49761
rect 42690 49629 42742 49681
rect 44715 49645 44767 49697
rect 41388 49388 41440 49440
rect 41388 49324 41440 49376
rect 41388 49260 41440 49312
rect 41388 49196 41440 49248
rect 41388 49132 41440 49184
rect 41388 49068 41440 49120
rect 53599 49378 53651 49430
rect 53663 49378 53715 49430
rect 39465 48902 39581 49018
rect 43111 48836 43163 48888
rect 44707 48677 44759 48729
rect 44707 48613 44759 48665
rect 44707 48549 44759 48601
rect 44707 48485 44759 48537
rect 38774 48421 38826 48473
rect 42186 48411 42238 48463
rect 44711 48181 44763 48233
rect 38219 48082 38271 48134
rect 39837 48082 39889 48134
rect 44711 48117 44763 48169
rect 42690 48029 42742 48081
rect 44711 48053 44763 48105
rect 66499 52556 66551 52608
rect 65060 49784 65112 49836
rect 62817 48546 62869 48598
rect 62817 48482 62869 48534
rect 62817 48418 62869 48470
rect 62817 48354 62869 48406
rect 62817 48290 62869 48342
rect 62817 48226 62869 48278
rect 60499 48065 60551 48117
rect 39465 47673 39581 47789
rect 41376 47581 41428 47633
rect 41376 47517 41428 47569
rect 41376 47453 41428 47505
rect 62743 48061 62795 48113
rect 64117 48065 64169 48117
rect 66499 48065 66551 48117
rect 99959 48115 100011 48167
rect 100023 48115 100075 48167
rect 100087 48115 100139 48167
rect 100151 48115 100203 48167
rect 100215 48115 100267 48167
rect 100279 48115 100331 48167
rect 100343 48115 100395 48167
rect 100407 48115 100459 48167
rect 100471 48115 100523 48167
rect 100535 48115 100587 48167
rect 100599 48115 100651 48167
rect 100663 48115 100715 48167
rect 100727 48115 100779 48167
rect 100791 48115 100843 48167
rect 100855 48115 100907 48167
rect 100919 48115 100971 48167
rect 100983 48115 101035 48167
rect 101047 48115 101099 48167
rect 101111 48115 101163 48167
rect 101175 48115 101227 48167
rect 101239 48115 101291 48167
rect 101303 48115 101355 48167
rect 101367 48115 101419 48167
rect 101431 48115 101483 48167
rect 101495 48115 101547 48167
rect 101559 48115 101611 48167
rect 101623 48115 101675 48167
rect 101687 48115 101739 48167
rect 101751 48115 101803 48167
rect 101815 48115 101867 48167
rect 101879 48115 101931 48167
rect 101943 48115 101995 48167
rect 102007 48115 102059 48167
rect 102071 48115 102123 48167
rect 102135 48115 102187 48167
rect 102199 48115 102251 48167
rect 102263 48115 102315 48167
rect 102327 48115 102379 48167
rect 102391 48115 102443 48167
rect 102455 48115 102507 48167
rect 102519 48115 102571 48167
rect 102583 48115 102635 48167
rect 102647 48115 102699 48167
rect 102711 48115 102763 48167
rect 102775 48115 102827 48167
rect 102839 48115 102891 48167
rect 102903 48115 102955 48167
rect 102967 48115 103019 48167
rect 103031 48115 103083 48167
rect 103095 48115 103147 48167
rect 103159 48115 103211 48167
rect 103223 48115 103275 48167
rect 92252 47830 92304 47882
rect 96451 47663 96503 47715
rect 94923 47579 94975 47631
rect 94923 47515 94975 47567
rect 96451 47599 96503 47651
rect 96451 47535 96503 47587
rect 43111 47236 43163 47288
rect 44714 47223 44766 47275
rect 44714 47159 44766 47211
rect 44714 47095 44766 47147
rect 65901 47297 65953 47349
rect 65965 47297 66017 47349
rect 44714 47031 44766 47083
rect 59650 47027 59702 47079
rect 67302 47027 67354 47079
rect 44714 46967 44766 47019
rect 44714 46903 44766 46955
rect 42186 46741 42238 46793
rect 45499 46740 45551 46792
rect 45563 46740 45615 46792
rect 44711 46571 44763 46623
rect 44711 46507 44763 46559
rect 42690 46429 42742 46481
rect 44711 46443 44763 46495
rect 51014 45635 51066 45687
rect 51078 45635 51130 45687
rect 53599 44773 53651 44825
rect 53663 44773 53715 44825
rect 18953 43022 19005 43074
rect 19017 43022 19069 43074
rect 19081 43022 19133 43074
rect 19145 43022 19197 43074
rect 19209 43022 19261 43074
rect 19273 43022 19325 43074
rect 19337 43022 19389 43074
rect 19401 43022 19453 43074
rect 19465 43022 19517 43074
rect 19529 43022 19581 43074
rect 19593 43022 19645 43074
rect 19657 43022 19709 43074
rect 19721 43022 19773 43074
rect 19785 43022 19837 43074
rect 19849 43022 19901 43074
rect 19913 43022 19965 43074
rect 19977 43022 20029 43074
rect 20041 43022 20093 43074
rect 20105 43022 20157 43074
rect 20169 43022 20221 43074
rect 20233 43022 20285 43074
rect 20297 43022 20349 43074
rect 20361 43022 20413 43074
rect 20425 43022 20477 43074
rect 20489 43022 20541 43074
rect 20553 43022 20605 43074
rect 20617 43022 20669 43074
rect 20681 43022 20733 43074
rect 20745 43022 20797 43074
rect 20809 43022 20861 43074
rect 20873 43022 20925 43074
rect 20937 43022 20989 43074
rect 21001 43022 21053 43074
rect 21065 43022 21117 43074
rect 21129 43022 21181 43074
rect 21193 43022 21245 43074
rect 21257 43022 21309 43074
rect 21321 43022 21373 43074
rect 21385 43022 21437 43074
rect 21449 43022 21501 43074
rect 21513 43022 21565 43074
rect 21577 43022 21629 43074
rect 21641 43022 21693 43074
rect 21705 43022 21757 43074
rect 21769 43022 21821 43074
rect 21833 43022 21885 43074
rect 21897 43022 21949 43074
rect 21961 43022 22013 43074
rect 22025 43022 22077 43074
rect 22089 43022 22141 43074
rect 22153 43022 22205 43074
rect 31648 41866 31700 41918
rect 31648 41802 31700 41854
rect 31648 41738 31700 41790
rect 31648 41674 31700 41726
rect 16526 41444 16706 41624
rect 56656 44073 56708 44125
rect 56656 44009 56708 44061
rect 58784 43374 58836 43426
rect 58784 43310 58836 43362
rect 25970 41482 26086 41598
rect 57333 41736 57385 41788
rect 56279 41489 56331 41541
rect 31654 41346 31706 41398
rect 31654 41282 31706 41334
rect 31654 41218 31706 41270
rect 61491 46007 61543 46059
rect 65322 46007 65374 46059
rect 61491 44915 61543 44967
rect 65322 44915 65374 44967
rect 62494 44073 62546 44125
rect 62494 44009 62546 44061
rect 66494 44073 66546 44125
rect 66494 44009 66546 44061
rect 60495 43310 60547 43362
rect 60161 43070 60213 43122
rect 61965 43064 62273 43180
rect 64494 43374 64546 43426
rect 64494 43310 64546 43362
rect 64185 43070 64237 43122
rect 56655 41185 56707 41237
rect 56655 41121 56707 41173
rect 58784 41185 58836 41237
rect 58784 41121 58836 41173
rect 61395 41253 61447 41305
rect 66081 43070 66133 43122
rect 94930 47162 94982 47214
rect 94930 47098 94982 47150
rect 94930 47034 94982 47086
rect 94930 46970 94982 47022
rect 96446 47168 96498 47220
rect 96446 47104 96498 47156
rect 96446 47040 96498 47092
rect 96446 46976 96498 47028
rect 92194 46632 92374 46812
rect 92862 46695 92914 46747
rect 92926 46695 92978 46747
rect 92990 46695 93042 46747
rect 93054 46695 93106 46747
rect 96451 46337 96503 46389
rect 94929 46243 94981 46295
rect 94929 46179 94981 46231
rect 96451 46273 96503 46325
rect 96451 46209 96503 46261
rect 104678 46548 104858 46728
rect 94924 45782 94976 45834
rect 94924 45718 94976 45770
rect 94924 45654 94976 45706
rect 96452 45802 96504 45854
rect 96452 45738 96504 45790
rect 96452 45674 96504 45726
rect 96452 45610 96504 45662
rect 92252 45549 92304 45601
rect 99957 45119 100009 45171
rect 100021 45119 100073 45171
rect 100085 45119 100137 45171
rect 100149 45119 100201 45171
rect 100213 45119 100265 45171
rect 100277 45119 100329 45171
rect 100341 45119 100393 45171
rect 100405 45119 100457 45171
rect 100469 45119 100521 45171
rect 100533 45119 100585 45171
rect 100597 45119 100649 45171
rect 100661 45119 100713 45171
rect 100725 45119 100777 45171
rect 100789 45119 100841 45171
rect 100853 45119 100905 45171
rect 100917 45119 100969 45171
rect 100981 45119 101033 45171
rect 101045 45119 101097 45171
rect 101109 45119 101161 45171
rect 101173 45119 101225 45171
rect 101237 45119 101289 45171
rect 101301 45119 101353 45171
rect 101365 45119 101417 45171
rect 101429 45119 101481 45171
rect 101493 45119 101545 45171
rect 101557 45119 101609 45171
rect 101621 45119 101673 45171
rect 101685 45119 101737 45171
rect 101749 45119 101801 45171
rect 101813 45119 101865 45171
rect 101877 45119 101929 45171
rect 101941 45119 101993 45171
rect 102005 45119 102057 45171
rect 102069 45119 102121 45171
rect 102133 45119 102185 45171
rect 102197 45119 102249 45171
rect 102261 45119 102313 45171
rect 102325 45119 102377 45171
rect 102389 45119 102441 45171
rect 102453 45119 102505 45171
rect 102517 45119 102569 45171
rect 102581 45119 102633 45171
rect 102645 45119 102697 45171
rect 102709 45119 102761 45171
rect 102773 45119 102825 45171
rect 102837 45119 102889 45171
rect 102901 45119 102953 45171
rect 102965 45119 103017 45171
rect 103029 45119 103081 45171
rect 103093 45119 103145 45171
rect 103157 45119 103209 45171
rect 103221 45119 103273 45171
rect 71788 44991 71840 45043
rect 80770 44180 80822 44232
rect 69473 44011 69589 44127
rect 68395 43312 68511 43428
rect 80789 43346 80841 43398
rect 67332 43022 67384 43074
rect 65380 42682 65432 42734
rect 70674 42652 70726 42704
rect 80758 42392 80810 42444
rect 80789 41516 80841 41568
rect 64493 41323 64545 41375
rect 63327 41253 63379 41305
rect 64493 41259 64545 41311
rect 66496 41323 66548 41375
rect 66496 41259 66548 41311
rect 70985 41323 71037 41375
rect 70985 41259 71037 41311
rect 71790 41047 71842 41099
rect 60493 40830 60545 40882
rect 60493 40766 60545 40818
rect 62493 40830 62545 40882
rect 62493 40766 62545 40818
rect 70377 40830 70429 40882
rect 70377 40766 70429 40818
rect 53174 40252 53226 40304
rect 57355 40274 68223 40454
rect 18923 40027 18975 40079
rect 18987 40027 19039 40079
rect 19051 40027 19103 40079
rect 19115 40027 19167 40079
rect 19179 40027 19231 40079
rect 19243 40027 19295 40079
rect 19307 40027 19359 40079
rect 19371 40027 19423 40079
rect 19435 40027 19487 40079
rect 19499 40027 19551 40079
rect 19563 40027 19615 40079
rect 19627 40027 19679 40079
rect 19691 40027 19743 40079
rect 19755 40027 19807 40079
rect 19819 40027 19871 40079
rect 19883 40027 19935 40079
rect 19947 40027 19999 40079
rect 20011 40027 20063 40079
rect 20075 40027 20127 40079
rect 20139 40027 20191 40079
rect 20203 40027 20255 40079
rect 20267 40027 20319 40079
rect 20331 40027 20383 40079
rect 20395 40027 20447 40079
rect 20459 40027 20511 40079
rect 20523 40027 20575 40079
rect 20587 40027 20639 40079
rect 20651 40027 20703 40079
rect 20715 40027 20767 40079
rect 20779 40027 20831 40079
rect 20843 40027 20895 40079
rect 20907 40027 20959 40079
rect 20971 40027 21023 40079
rect 21035 40027 21087 40079
rect 21099 40027 21151 40079
rect 21163 40027 21215 40079
rect 21227 40027 21279 40079
rect 21291 40027 21343 40079
rect 21355 40027 21407 40079
rect 21419 40027 21471 40079
rect 21483 40027 21535 40079
rect 21547 40027 21599 40079
rect 21611 40027 21663 40079
rect 21675 40027 21727 40079
rect 21739 40027 21791 40079
rect 21803 40027 21855 40079
rect 21867 40027 21919 40079
rect 21931 40027 21983 40079
rect 21995 40027 22047 40079
rect 22059 40027 22111 40079
rect 22123 40027 22175 40079
rect 22187 40027 22239 40079
rect 51314 39672 51366 39724
rect 53180 39105 53232 39157
rect 56416 39106 56468 39158
rect 53965 38950 54017 39002
rect 53965 38886 54017 38938
rect 53965 38822 54017 38874
rect 53965 38758 54017 38810
rect 31587 38393 31639 38445
rect 31587 38329 31639 38381
rect 31587 38265 31639 38317
rect 52201 38401 52253 38453
rect 52201 38337 52253 38389
rect 52201 38273 52253 38325
rect 31587 38201 31639 38253
rect 24109 38002 24225 38118
rect 44036 38105 44088 38157
rect 50556 38105 50608 38157
rect 53180 38109 53232 38161
rect 38877 38037 38929 38089
rect 31586 37867 31638 37919
rect 31586 37803 31638 37855
rect 31586 37739 31638 37791
rect 52193 37944 52245 37996
rect 52193 37880 52245 37932
rect 52193 37816 52245 37868
rect 52193 37752 52245 37804
rect 55301 37085 55353 37137
rect 55301 37021 55353 37073
rect 55301 36957 55353 37009
rect 50556 36856 50608 36908
rect 51249 36856 51301 36908
rect 55301 36893 55353 36945
rect 55301 36829 55353 36881
rect 55301 36765 55353 36817
rect 53180 36605 53232 36657
rect 56815 36607 56867 36659
rect 55602 36373 55654 36425
rect 51249 36183 51301 36235
rect 55342 35490 55394 35542
rect 55342 35426 55394 35478
rect 55342 35362 55394 35414
rect 55342 35298 55394 35350
rect 55342 35234 55394 35286
rect 55342 35170 55394 35222
rect 53679 35004 53731 35056
rect 56815 35005 56867 35057
rect 51249 34913 51301 34965
rect 50954 34791 51006 34843
rect 51018 34791 51070 34843
rect 51082 34791 51134 34843
rect 51418 34790 51470 34842
rect 51482 34790 51534 34842
rect 51546 34790 51598 34842
rect 51610 34790 51662 34842
rect 55602 34747 55654 34799
rect 57143 40139 57259 40182
rect 57143 40105 57182 40139
rect 57182 40105 57216 40139
rect 57216 40105 57259 40139
rect 57143 40067 57259 40105
rect 57143 40033 57182 40067
rect 57182 40033 57216 40067
rect 57216 40033 57259 40067
rect 57143 39995 57259 40033
rect 57143 39961 57182 39995
rect 57182 39961 57216 39995
rect 57216 39961 57259 39995
rect 57143 39923 57259 39961
rect 57143 39889 57182 39923
rect 57182 39889 57216 39923
rect 57216 39889 57259 39923
rect 57143 39851 57259 39889
rect 57143 39817 57182 39851
rect 57182 39817 57216 39851
rect 57216 39817 57259 39851
rect 57143 39779 57259 39817
rect 57143 39745 57182 39779
rect 57182 39745 57216 39779
rect 57216 39745 57259 39779
rect 57143 39707 57259 39745
rect 57143 39673 57182 39707
rect 57182 39673 57216 39707
rect 57216 39673 57259 39707
rect 57143 39635 57259 39673
rect 57143 39601 57182 39635
rect 57182 39601 57216 39635
rect 57216 39601 57259 39635
rect 57143 39563 57259 39601
rect 57143 39529 57182 39563
rect 57182 39529 57216 39563
rect 57216 39529 57259 39563
rect 57143 39491 57259 39529
rect 57143 39457 57182 39491
rect 57182 39457 57216 39491
rect 57216 39457 57259 39491
rect 57143 39419 57259 39457
rect 57143 39385 57182 39419
rect 57182 39385 57216 39419
rect 57216 39385 57259 39419
rect 57143 39347 57259 39385
rect 57143 39313 57182 39347
rect 57182 39313 57216 39347
rect 57216 39313 57259 39347
rect 57143 39275 57259 39313
rect 57143 39241 57182 39275
rect 57182 39241 57216 39275
rect 57216 39241 57259 39275
rect 57143 39203 57259 39241
rect 57143 39169 57182 39203
rect 57182 39169 57216 39203
rect 57216 39169 57259 39203
rect 57143 39131 57259 39169
rect 57143 39097 57182 39131
rect 57182 39097 57216 39131
rect 57216 39097 57259 39131
rect 57143 39059 57259 39097
rect 57143 39025 57182 39059
rect 57182 39025 57216 39059
rect 57216 39025 57259 39059
rect 57143 38987 57259 39025
rect 57143 38953 57182 38987
rect 57182 38953 57216 38987
rect 57216 38953 57259 38987
rect 57143 38915 57259 38953
rect 57143 38881 57182 38915
rect 57182 38881 57216 38915
rect 57216 38881 57259 38915
rect 57143 38843 57259 38881
rect 57143 38809 57182 38843
rect 57182 38809 57216 38843
rect 57216 38809 57259 38843
rect 57143 38771 57259 38809
rect 57143 38737 57182 38771
rect 57182 38737 57216 38771
rect 57216 38737 57259 38771
rect 57143 38699 57259 38737
rect 57143 38665 57182 38699
rect 57182 38665 57216 38699
rect 57216 38665 57259 38699
rect 57143 38627 57259 38665
rect 57143 38593 57182 38627
rect 57182 38593 57216 38627
rect 57216 38593 57259 38627
rect 57143 38555 57259 38593
rect 57143 38521 57182 38555
rect 57182 38521 57216 38555
rect 57216 38521 57259 38555
rect 57143 38483 57259 38521
rect 57143 38449 57182 38483
rect 57182 38449 57216 38483
rect 57216 38449 57259 38483
rect 57143 38411 57259 38449
rect 57143 38377 57182 38411
rect 57182 38377 57216 38411
rect 57216 38377 57259 38411
rect 57143 38339 57259 38377
rect 57143 38305 57182 38339
rect 57182 38305 57216 38339
rect 57216 38305 57259 38339
rect 57143 38267 57259 38305
rect 57143 38233 57182 38267
rect 57182 38233 57216 38267
rect 57216 38233 57259 38267
rect 57143 38195 57259 38233
rect 57143 38161 57182 38195
rect 57182 38161 57216 38195
rect 57216 38161 57259 38195
rect 57143 38123 57259 38161
rect 57143 38089 57182 38123
rect 57182 38089 57216 38123
rect 57216 38089 57259 38123
rect 57143 38051 57259 38089
rect 57143 38017 57182 38051
rect 57182 38017 57216 38051
rect 57216 38017 57259 38051
rect 57143 37979 57259 38017
rect 57143 37945 57182 37979
rect 57182 37945 57216 37979
rect 57216 37945 57259 37979
rect 57143 37907 57259 37945
rect 57143 37873 57182 37907
rect 57182 37873 57216 37907
rect 57216 37873 57259 37907
rect 57143 37835 57259 37873
rect 57143 37801 57182 37835
rect 57182 37801 57216 37835
rect 57216 37801 57259 37835
rect 57143 37763 57259 37801
rect 57143 37729 57182 37763
rect 57182 37729 57216 37763
rect 57216 37729 57259 37763
rect 57143 37691 57259 37729
rect 57143 37657 57182 37691
rect 57182 37657 57216 37691
rect 57216 37657 57259 37691
rect 57143 37619 57259 37657
rect 57143 37585 57182 37619
rect 57182 37585 57216 37619
rect 57216 37585 57259 37619
rect 57143 37547 57259 37585
rect 57143 37513 57182 37547
rect 57182 37513 57216 37547
rect 57216 37513 57259 37547
rect 57143 37475 57259 37513
rect 57143 37441 57182 37475
rect 57182 37441 57216 37475
rect 57216 37441 57259 37475
rect 57143 37403 57259 37441
rect 57143 37369 57182 37403
rect 57182 37369 57216 37403
rect 57216 37369 57259 37403
rect 57143 37331 57259 37369
rect 57143 37297 57182 37331
rect 57182 37297 57216 37331
rect 57216 37297 57259 37331
rect 57143 37259 57259 37297
rect 57143 37225 57182 37259
rect 57182 37225 57216 37259
rect 57216 37225 57259 37259
rect 57143 37187 57259 37225
rect 57143 37153 57182 37187
rect 57182 37153 57216 37187
rect 57216 37153 57259 37187
rect 57143 37115 57259 37153
rect 57143 37081 57182 37115
rect 57182 37081 57216 37115
rect 57216 37081 57259 37115
rect 57143 37043 57259 37081
rect 57143 37009 57182 37043
rect 57182 37009 57216 37043
rect 57216 37009 57259 37043
rect 57143 36971 57259 37009
rect 57143 36937 57182 36971
rect 57182 36937 57216 36971
rect 57216 36937 57259 36971
rect 57143 36899 57259 36937
rect 57143 36865 57182 36899
rect 57182 36865 57216 36899
rect 57216 36865 57259 36899
rect 57143 36827 57259 36865
rect 57143 36793 57182 36827
rect 57182 36793 57216 36827
rect 57216 36793 57259 36827
rect 57143 36755 57259 36793
rect 57143 36721 57182 36755
rect 57182 36721 57216 36755
rect 57216 36721 57259 36755
rect 57143 36683 57259 36721
rect 57143 36649 57182 36683
rect 57182 36649 57216 36683
rect 57216 36649 57259 36683
rect 57143 36611 57259 36649
rect 57143 36577 57182 36611
rect 57182 36577 57216 36611
rect 57216 36577 57259 36611
rect 57143 36539 57259 36577
rect 57143 36505 57182 36539
rect 57182 36505 57216 36539
rect 57216 36505 57259 36539
rect 57143 36467 57259 36505
rect 57143 36433 57182 36467
rect 57182 36433 57216 36467
rect 57216 36433 57259 36467
rect 57143 36395 57259 36433
rect 57143 36361 57182 36395
rect 57182 36361 57216 36395
rect 57216 36361 57259 36395
rect 57143 36323 57259 36361
rect 57143 36289 57182 36323
rect 57182 36289 57216 36323
rect 57216 36289 57259 36323
rect 57143 36251 57259 36289
rect 57143 36217 57182 36251
rect 57182 36217 57216 36251
rect 57216 36217 57259 36251
rect 57143 36179 57259 36217
rect 57143 36145 57182 36179
rect 57182 36145 57216 36179
rect 57216 36145 57259 36179
rect 57143 36107 57259 36145
rect 57143 36073 57182 36107
rect 57182 36073 57216 36107
rect 57216 36073 57259 36107
rect 57143 36035 57259 36073
rect 57143 36001 57182 36035
rect 57182 36001 57216 36035
rect 57216 36001 57259 36035
rect 57143 35963 57259 36001
rect 57143 35929 57182 35963
rect 57182 35929 57216 35963
rect 57216 35929 57259 35963
rect 57143 35891 57259 35929
rect 57143 35857 57182 35891
rect 57182 35857 57216 35891
rect 57216 35857 57259 35891
rect 57143 35819 57259 35857
rect 57143 35785 57182 35819
rect 57182 35785 57216 35819
rect 57216 35785 57259 35819
rect 57143 35747 57259 35785
rect 57143 35713 57182 35747
rect 57182 35713 57216 35747
rect 57216 35713 57259 35747
rect 57143 35675 57259 35713
rect 57143 35641 57182 35675
rect 57182 35641 57216 35675
rect 57216 35641 57259 35675
rect 57143 35603 57259 35641
rect 57143 35569 57182 35603
rect 57182 35569 57216 35603
rect 57216 35569 57259 35603
rect 57143 35531 57259 35569
rect 57143 35497 57182 35531
rect 57182 35497 57216 35531
rect 57216 35497 57259 35531
rect 57143 35459 57259 35497
rect 57143 35425 57182 35459
rect 57182 35425 57216 35459
rect 57216 35425 57259 35459
rect 57143 35387 57259 35425
rect 57143 35353 57182 35387
rect 57182 35353 57216 35387
rect 57216 35353 57259 35387
rect 57143 35315 57259 35353
rect 57143 35281 57182 35315
rect 57182 35281 57216 35315
rect 57216 35281 57259 35315
rect 57143 35243 57259 35281
rect 57143 35209 57182 35243
rect 57182 35209 57216 35243
rect 57216 35209 57259 35243
rect 57143 35171 57259 35209
rect 57143 35137 57182 35171
rect 57182 35137 57216 35171
rect 57216 35137 57259 35171
rect 57143 35099 57259 35137
rect 57143 35065 57182 35099
rect 57182 35065 57216 35099
rect 57216 35065 57259 35099
rect 57143 35027 57259 35065
rect 57143 34993 57182 35027
rect 57182 34993 57216 35027
rect 57216 34993 57259 35027
rect 57143 34955 57259 34993
rect 57143 34921 57182 34955
rect 57182 34921 57216 34955
rect 57216 34921 57259 34955
rect 57143 34883 57259 34921
rect 57143 34849 57182 34883
rect 57182 34849 57216 34883
rect 57216 34849 57259 34883
rect 57143 34811 57259 34849
rect 57143 34777 57182 34811
rect 57182 34777 57216 34811
rect 57216 34777 57259 34811
rect 57143 34739 57259 34777
rect 57143 34705 57182 34739
rect 57182 34705 57216 34739
rect 57216 34705 57259 34739
rect 57143 34690 57259 34705
rect 68355 40144 68471 40185
rect 68355 40110 68397 40144
rect 68397 40110 68431 40144
rect 68431 40110 68471 40144
rect 68355 40072 68471 40110
rect 68355 40038 68397 40072
rect 68397 40038 68431 40072
rect 68431 40038 68471 40072
rect 68355 40000 68471 40038
rect 68355 39966 68397 40000
rect 68397 39966 68431 40000
rect 68431 39966 68471 40000
rect 68355 39928 68471 39966
rect 68355 39894 68397 39928
rect 68397 39894 68431 39928
rect 68431 39894 68471 39928
rect 68355 39856 68471 39894
rect 68355 39822 68397 39856
rect 68397 39822 68431 39856
rect 68431 39822 68471 39856
rect 68355 39784 68471 39822
rect 68355 39750 68397 39784
rect 68397 39750 68431 39784
rect 68431 39750 68471 39784
rect 68355 39712 68471 39750
rect 68355 39678 68397 39712
rect 68397 39678 68431 39712
rect 68431 39678 68471 39712
rect 68355 39640 68471 39678
rect 68355 39606 68397 39640
rect 68397 39606 68431 39640
rect 68431 39606 68471 39640
rect 68355 39568 68471 39606
rect 68355 39534 68397 39568
rect 68397 39534 68431 39568
rect 68431 39534 68471 39568
rect 68355 39496 68471 39534
rect 68355 39462 68397 39496
rect 68397 39462 68431 39496
rect 68431 39462 68471 39496
rect 68355 39424 68471 39462
rect 68355 39390 68397 39424
rect 68397 39390 68431 39424
rect 68431 39390 68471 39424
rect 68355 39352 68471 39390
rect 68355 39318 68397 39352
rect 68397 39318 68431 39352
rect 68431 39318 68471 39352
rect 68355 39280 68471 39318
rect 68355 39246 68397 39280
rect 68397 39246 68431 39280
rect 68431 39246 68471 39280
rect 68355 39208 68471 39246
rect 68355 39174 68397 39208
rect 68397 39174 68431 39208
rect 68431 39174 68471 39208
rect 68355 39136 68471 39174
rect 68355 39102 68397 39136
rect 68397 39102 68431 39136
rect 68431 39102 68471 39136
rect 68355 39064 68471 39102
rect 68355 39030 68397 39064
rect 68397 39030 68431 39064
rect 68431 39030 68471 39064
rect 68355 38992 68471 39030
rect 68355 38958 68397 38992
rect 68397 38958 68431 38992
rect 68431 38958 68471 38992
rect 68355 38920 68471 38958
rect 68355 38886 68397 38920
rect 68397 38886 68431 38920
rect 68431 38886 68471 38920
rect 68355 38848 68471 38886
rect 68355 38814 68397 38848
rect 68397 38814 68431 38848
rect 68431 38814 68471 38848
rect 68355 38776 68471 38814
rect 68355 38742 68397 38776
rect 68397 38742 68431 38776
rect 68431 38742 68471 38776
rect 68355 38704 68471 38742
rect 68355 38670 68397 38704
rect 68397 38670 68431 38704
rect 68431 38670 68471 38704
rect 68355 38632 68471 38670
rect 68355 38598 68397 38632
rect 68397 38598 68431 38632
rect 68431 38598 68471 38632
rect 68355 38560 68471 38598
rect 68355 38526 68397 38560
rect 68397 38526 68431 38560
rect 68431 38526 68471 38560
rect 68355 38488 68471 38526
rect 68355 38469 68397 38488
rect 68397 38469 68431 38488
rect 68431 38469 68471 38488
rect 80786 39752 80838 39804
rect 78028 39460 78080 39512
rect 71790 39192 71842 39244
rect 68356 37942 68472 37968
rect 68356 37908 68397 37942
rect 68397 37908 68431 37942
rect 68431 37908 68472 37942
rect 68356 37870 68472 37908
rect 68356 37836 68397 37870
rect 68397 37836 68431 37870
rect 68431 37836 68472 37870
rect 68356 37798 68472 37836
rect 68356 37764 68397 37798
rect 68397 37764 68431 37798
rect 68431 37764 68472 37798
rect 68356 37726 68472 37764
rect 68356 37692 68397 37726
rect 68397 37692 68431 37726
rect 68431 37692 68472 37726
rect 68356 37654 68472 37692
rect 68356 37620 68397 37654
rect 68397 37620 68431 37654
rect 68431 37620 68472 37654
rect 68356 37582 68472 37620
rect 68356 37548 68397 37582
rect 68397 37548 68431 37582
rect 68431 37548 68472 37582
rect 68356 37510 68472 37548
rect 68356 37476 68397 37510
rect 68397 37476 68431 37510
rect 68431 37476 68472 37510
rect 68356 37438 68472 37476
rect 68356 37404 68397 37438
rect 68397 37404 68431 37438
rect 68431 37404 68472 37438
rect 68356 37366 68472 37404
rect 68356 37332 68397 37366
rect 68397 37332 68431 37366
rect 68431 37332 68472 37366
rect 68356 37294 68472 37332
rect 68356 37260 68397 37294
rect 68397 37260 68431 37294
rect 68431 37260 68472 37294
rect 68356 37222 68472 37260
rect 68356 37188 68397 37222
rect 68397 37188 68431 37222
rect 68431 37188 68472 37222
rect 68356 37150 68472 37188
rect 68356 37116 68397 37150
rect 68397 37116 68431 37150
rect 68431 37116 68472 37150
rect 68356 37078 68472 37116
rect 68356 37044 68397 37078
rect 68397 37044 68431 37078
rect 68431 37044 68472 37078
rect 68356 37020 68472 37044
rect 71785 37929 71837 37981
rect 80786 37961 80838 38013
rect 71790 37492 71842 37544
rect 80785 36970 80837 37022
rect 71802 36144 71854 36196
rect 80791 36154 80843 36206
rect 68356 36113 68472 36122
rect 68356 36079 68397 36113
rect 68397 36079 68431 36113
rect 68431 36079 68472 36113
rect 68356 36041 68472 36079
rect 68356 36007 68397 36041
rect 68397 36007 68431 36041
rect 68431 36007 68472 36041
rect 68356 35969 68472 36007
rect 68356 35935 68397 35969
rect 68397 35935 68431 35969
rect 68431 35935 68472 35969
rect 68356 35897 68472 35935
rect 68356 35863 68397 35897
rect 68397 35863 68431 35897
rect 68431 35863 68472 35897
rect 68356 35825 68472 35863
rect 68356 35791 68397 35825
rect 68397 35791 68431 35825
rect 68431 35791 68472 35825
rect 68356 35753 68472 35791
rect 68356 35719 68397 35753
rect 68397 35719 68431 35753
rect 68431 35719 68472 35753
rect 68356 35681 68472 35719
rect 68356 35647 68397 35681
rect 68397 35647 68431 35681
rect 68431 35647 68472 35681
rect 68356 35609 68472 35647
rect 68356 35575 68397 35609
rect 68397 35575 68431 35609
rect 68431 35575 68472 35609
rect 68356 35537 68472 35575
rect 68356 35503 68397 35537
rect 68397 35503 68431 35537
rect 68431 35503 68472 35537
rect 68356 35465 68472 35503
rect 68356 35431 68397 35465
rect 68397 35431 68431 35465
rect 68431 35431 68472 35465
rect 68356 35393 68472 35431
rect 68356 35366 68397 35393
rect 68397 35366 68431 35393
rect 68431 35366 68472 35393
rect 71792 35640 71844 35692
rect 80789 35483 80841 35535
rect 51249 34371 51301 34423
rect 56416 34372 56468 34424
rect 71791 34347 71843 34399
rect 80791 34344 80843 34396
rect 55341 33887 55393 33939
rect 55341 33823 55393 33875
rect 55341 33759 55393 33811
rect 55341 33695 55393 33747
rect 55341 33631 55393 33683
rect 50956 33548 51008 33600
rect 51020 33548 51072 33600
rect 51084 33548 51136 33600
rect 51386 33548 51438 33600
rect 51450 33548 51502 33600
rect 51514 33548 51566 33600
rect 51578 33548 51630 33600
rect 51642 33548 51694 33600
rect 55341 33567 55393 33619
rect 51249 33422 51301 33474
rect 53180 33407 53232 33459
rect 55945 33405 55997 33457
rect 62317 33387 62369 33439
rect 81644 33388 81696 33440
rect 55602 33089 55654 33141
rect 55344 32286 55396 32338
rect 55344 32222 55396 32274
rect 51247 32138 51299 32190
rect 55344 32158 55396 32210
rect 55344 32094 55396 32146
rect 55344 32030 55396 32082
rect 55344 31966 55396 32018
rect 53679 31805 53731 31857
rect 55945 31805 55997 31857
rect 80302 31814 80354 31866
rect 50535 31555 50587 31607
rect 51247 31559 51299 31611
rect 55602 31550 55654 31602
rect 49893 31055 50329 31235
rect 55602 31208 55654 31260
rect 55602 31144 55654 31196
rect 55602 31080 55654 31132
rect 55602 31016 55654 31068
rect 31584 30630 31636 30682
rect 31584 30566 31636 30618
rect 31584 30502 31636 30554
rect 31584 30438 31636 30490
rect 52191 30635 52243 30687
rect 52191 30571 52243 30623
rect 52191 30507 52243 30559
rect 52191 30443 52243 30495
rect 55602 30415 55654 30467
rect 25970 30237 26086 30353
rect 38849 30267 38901 30319
rect 44025 30277 44077 30329
rect 50535 30277 50587 30329
rect 53679 30280 53731 30332
rect 31583 30143 31635 30195
rect 31583 30079 31635 30131
rect 31583 30015 31635 30067
rect 31583 29951 31635 30003
rect 52194 30116 52246 30168
rect 52194 30052 52246 30104
rect 52194 29988 52246 30040
rect 53679 29693 53731 29745
rect 56416 29693 56468 29745
rect 53916 29528 53968 29580
rect 53916 29464 53968 29516
rect 53916 29400 53968 29452
rect 53916 29336 53968 29388
rect 55945 29099 55997 29151
rect 53673 29011 53725 29063
rect 92124 32247 92176 32299
rect 97208 32087 97260 32139
rect 95678 31993 95730 32045
rect 95678 31929 95730 31981
rect 97208 32023 97260 32075
rect 97208 31959 97260 32011
rect 93420 31843 93472 31895
rect 93484 31843 93536 31895
rect 93548 31843 93600 31895
rect 90846 31615 90898 31667
rect 95676 31529 95728 31581
rect 95676 31465 95728 31517
rect 95676 31401 95728 31453
rect 97195 31542 97247 31594
rect 97195 31478 97247 31530
rect 97195 31414 97247 31466
rect 93482 31302 93534 31354
rect 93546 31302 93598 31354
rect 92128 31187 92180 31239
rect 99698 31183 99750 31235
rect 99762 31183 99814 31235
rect 99826 31183 99878 31235
rect 99890 31183 99942 31235
rect 99954 31183 100006 31235
rect 100018 31183 100070 31235
rect 100082 31183 100134 31235
rect 100146 31183 100198 31235
rect 100210 31183 100262 31235
rect 100274 31183 100326 31235
rect 100338 31183 100390 31235
rect 100402 31183 100454 31235
rect 100466 31183 100518 31235
rect 100530 31183 100582 31235
rect 100594 31183 100646 31235
rect 100658 31183 100710 31235
rect 100722 31183 100774 31235
rect 100786 31183 100838 31235
rect 100850 31183 100902 31235
rect 100914 31183 100966 31235
rect 100978 31183 101030 31235
rect 101042 31183 101094 31235
rect 101106 31183 101158 31235
rect 101170 31183 101222 31235
rect 101234 31183 101286 31235
rect 101298 31183 101350 31235
rect 101362 31183 101414 31235
rect 101426 31183 101478 31235
rect 101490 31183 101542 31235
rect 101554 31183 101606 31235
rect 101618 31183 101670 31235
rect 101682 31183 101734 31235
rect 101746 31183 101798 31235
rect 101810 31183 101862 31235
rect 101874 31183 101926 31235
rect 101938 31183 101990 31235
rect 102002 31183 102054 31235
rect 102066 31183 102118 31235
rect 102130 31183 102182 31235
rect 102194 31183 102246 31235
rect 102258 31183 102310 31235
rect 102322 31183 102374 31235
rect 102386 31183 102438 31235
rect 102450 31183 102502 31235
rect 102514 31183 102566 31235
rect 102578 31183 102630 31235
rect 102642 31183 102694 31235
rect 102706 31183 102758 31235
rect 102770 31183 102822 31235
rect 102834 31183 102886 31235
rect 102898 31183 102950 31235
rect 102962 31183 103014 31235
rect 92127 30918 92179 30970
rect 93462 30754 93514 30806
rect 97200 30751 97252 30803
rect 95678 30672 95730 30724
rect 95678 30608 95730 30660
rect 97200 30687 97252 30739
rect 97200 30623 97252 30675
rect 81644 30276 81696 30328
rect 90834 30276 90886 30328
rect 94087 30213 94139 30265
rect 95671 30198 95723 30250
rect 95671 30134 95723 30186
rect 95671 30070 95723 30122
rect 97200 30195 97252 30247
rect 97200 30131 97252 30183
rect 97200 30067 97252 30119
rect 92127 29849 92179 29901
rect 93095 29671 93147 29723
rect 93159 29671 93211 29723
rect 104595 29614 104775 29794
rect 92124 29526 92176 29578
rect 97217 29371 97269 29423
rect 95679 29282 95731 29334
rect 95679 29218 95731 29270
rect 97217 29307 97269 29359
rect 97217 29243 97269 29295
rect 93628 29123 93680 29175
rect 93692 29123 93744 29175
rect 93756 29123 93808 29175
rect 80302 28885 80354 28937
rect 90836 28885 90888 28937
rect 95670 28845 95722 28897
rect 95670 28781 95722 28833
rect 95670 28717 95722 28769
rect 97200 28823 97252 28875
rect 97200 28759 97252 28811
rect 97200 28695 97252 28747
rect 93472 28580 93524 28632
rect 93536 28580 93588 28632
rect 92135 28456 92187 28508
rect 56815 27759 56867 27811
rect 80526 26376 80578 26428
rect 79683 25066 79735 25118
rect 57446 24113 78170 24229
rect 92124 28151 92176 28203
rect 99715 28184 99767 28236
rect 99779 28184 99831 28236
rect 99843 28184 99895 28236
rect 99907 28184 99959 28236
rect 99971 28184 100023 28236
rect 100035 28184 100087 28236
rect 100099 28184 100151 28236
rect 100163 28184 100215 28236
rect 100227 28184 100279 28236
rect 100291 28184 100343 28236
rect 100355 28184 100407 28236
rect 100419 28184 100471 28236
rect 100483 28184 100535 28236
rect 100547 28184 100599 28236
rect 100611 28184 100663 28236
rect 100675 28184 100727 28236
rect 100739 28184 100791 28236
rect 100803 28184 100855 28236
rect 100867 28184 100919 28236
rect 100931 28184 100983 28236
rect 100995 28184 101047 28236
rect 101059 28184 101111 28236
rect 101123 28184 101175 28236
rect 101187 28184 101239 28236
rect 101251 28184 101303 28236
rect 101315 28184 101367 28236
rect 101379 28184 101431 28236
rect 101443 28184 101495 28236
rect 101507 28184 101559 28236
rect 101571 28184 101623 28236
rect 101635 28184 101687 28236
rect 101699 28184 101751 28236
rect 101763 28184 101815 28236
rect 101827 28184 101879 28236
rect 101891 28184 101943 28236
rect 101955 28184 102007 28236
rect 102019 28184 102071 28236
rect 102083 28184 102135 28236
rect 102147 28184 102199 28236
rect 102211 28184 102263 28236
rect 102275 28184 102327 28236
rect 102339 28184 102391 28236
rect 102403 28184 102455 28236
rect 102467 28184 102519 28236
rect 102531 28184 102583 28236
rect 102595 28184 102647 28236
rect 102659 28184 102711 28236
rect 102723 28184 102775 28236
rect 102787 28184 102839 28236
rect 102851 28184 102903 28236
rect 102915 28184 102967 28236
rect 102979 28184 103031 28236
rect 94088 28037 94140 28089
rect 97207 27992 97259 28044
rect 95679 27885 95731 27937
rect 95679 27821 95731 27873
rect 97207 27928 97259 27980
rect 97207 27864 97259 27916
rect 93458 27491 93510 27543
rect 93522 27491 93574 27543
rect 95673 27445 95725 27497
rect 95673 27381 95725 27433
rect 95673 27317 95725 27369
rect 97197 27439 97249 27491
rect 97197 27375 97249 27427
rect 97197 27311 97249 27363
rect 92131 27086 92183 27138
rect 92124 25307 92176 25359
rect 97208 25147 97260 25199
rect 95678 25053 95730 25105
rect 95678 24989 95730 25041
rect 97208 25083 97260 25135
rect 97208 25019 97260 25071
rect 93420 24903 93472 24955
rect 93484 24903 93536 24955
rect 93548 24903 93600 24955
rect 83106 24674 83158 24726
rect 90835 24674 90887 24726
rect 95676 24589 95728 24641
rect 95676 24525 95728 24577
rect 95676 24461 95728 24513
rect 97195 24602 97247 24654
rect 97195 24538 97247 24590
rect 97195 24474 97247 24526
rect 93482 24362 93534 24414
rect 93546 24362 93598 24414
rect 92128 24247 92180 24299
rect 99700 24250 99752 24302
rect 99764 24250 99816 24302
rect 99828 24250 99880 24302
rect 99892 24250 99944 24302
rect 99956 24250 100008 24302
rect 100020 24250 100072 24302
rect 100084 24250 100136 24302
rect 100148 24250 100200 24302
rect 100212 24250 100264 24302
rect 100276 24250 100328 24302
rect 100340 24250 100392 24302
rect 100404 24250 100456 24302
rect 100468 24250 100520 24302
rect 100532 24250 100584 24302
rect 100596 24250 100648 24302
rect 100660 24250 100712 24302
rect 100724 24250 100776 24302
rect 100788 24250 100840 24302
rect 100852 24250 100904 24302
rect 100916 24250 100968 24302
rect 100980 24250 101032 24302
rect 101044 24250 101096 24302
rect 101108 24250 101160 24302
rect 101172 24250 101224 24302
rect 101236 24250 101288 24302
rect 101300 24250 101352 24302
rect 101364 24250 101416 24302
rect 101428 24250 101480 24302
rect 101492 24250 101544 24302
rect 101556 24250 101608 24302
rect 101620 24250 101672 24302
rect 101684 24250 101736 24302
rect 101748 24250 101800 24302
rect 101812 24250 101864 24302
rect 101876 24250 101928 24302
rect 101940 24250 101992 24302
rect 102004 24250 102056 24302
rect 102068 24250 102120 24302
rect 102132 24250 102184 24302
rect 102196 24250 102248 24302
rect 102260 24250 102312 24302
rect 102324 24250 102376 24302
rect 102388 24250 102440 24302
rect 102452 24250 102504 24302
rect 102516 24250 102568 24302
rect 102580 24250 102632 24302
rect 102644 24250 102696 24302
rect 102708 24250 102760 24302
rect 102772 24250 102824 24302
rect 102836 24250 102888 24302
rect 102900 24250 102952 24302
rect 102964 24250 103016 24302
rect 92127 23978 92179 24030
rect 93462 23814 93514 23866
rect 97200 23811 97252 23863
rect 95678 23732 95730 23784
rect 95678 23668 95730 23720
rect 97200 23747 97252 23799
rect 97200 23683 97252 23735
rect 80526 23329 80578 23381
rect 90835 23335 90887 23387
rect 94087 23273 94139 23325
rect 95671 23258 95723 23310
rect 95671 23194 95723 23246
rect 95671 23130 95723 23182
rect 97200 23255 97252 23307
rect 97200 23191 97252 23243
rect 97200 23127 97252 23179
rect 92127 22909 92179 22961
rect 93095 22731 93147 22783
rect 93159 22731 93211 22783
rect 104611 22674 104791 22854
rect 92124 22586 92176 22638
rect 97217 22431 97269 22483
rect 95679 22342 95731 22394
rect 95679 22278 95731 22330
rect 97217 22367 97269 22419
rect 97217 22303 97269 22355
rect 93628 22183 93680 22235
rect 93692 22183 93744 22235
rect 93756 22183 93808 22235
rect 79684 21952 79736 22004
rect 90844 21949 90896 22001
rect 95670 21905 95722 21957
rect 95670 21841 95722 21893
rect 95670 21777 95722 21829
rect 97200 21883 97252 21935
rect 97200 21819 97252 21871
rect 97200 21755 97252 21807
rect 93472 21640 93524 21692
rect 93536 21640 93588 21692
rect 92135 21516 92187 21568
rect 92124 21211 92176 21263
rect 99696 21244 99748 21296
rect 99760 21244 99812 21296
rect 99824 21244 99876 21296
rect 99888 21244 99940 21296
rect 99952 21244 100004 21296
rect 100016 21244 100068 21296
rect 100080 21244 100132 21296
rect 100144 21244 100196 21296
rect 100208 21244 100260 21296
rect 100272 21244 100324 21296
rect 100336 21244 100388 21296
rect 100400 21244 100452 21296
rect 100464 21244 100516 21296
rect 100528 21244 100580 21296
rect 100592 21244 100644 21296
rect 100656 21244 100708 21296
rect 100720 21244 100772 21296
rect 100784 21244 100836 21296
rect 100848 21244 100900 21296
rect 100912 21244 100964 21296
rect 100976 21244 101028 21296
rect 101040 21244 101092 21296
rect 101104 21244 101156 21296
rect 101168 21244 101220 21296
rect 101232 21244 101284 21296
rect 101296 21244 101348 21296
rect 101360 21244 101412 21296
rect 101424 21244 101476 21296
rect 101488 21244 101540 21296
rect 101552 21244 101604 21296
rect 101616 21244 101668 21296
rect 101680 21244 101732 21296
rect 101744 21244 101796 21296
rect 101808 21244 101860 21296
rect 101872 21244 101924 21296
rect 101936 21244 101988 21296
rect 102000 21244 102052 21296
rect 102064 21244 102116 21296
rect 102128 21244 102180 21296
rect 102192 21244 102244 21296
rect 102256 21244 102308 21296
rect 102320 21244 102372 21296
rect 102384 21244 102436 21296
rect 102448 21244 102500 21296
rect 102512 21244 102564 21296
rect 102576 21244 102628 21296
rect 102640 21244 102692 21296
rect 102704 21244 102756 21296
rect 102768 21244 102820 21296
rect 102832 21244 102884 21296
rect 102896 21244 102948 21296
rect 102960 21244 103012 21296
rect 94088 21097 94140 21149
rect 97207 21052 97259 21104
rect 95679 20945 95731 20997
rect 95679 20881 95731 20933
rect 97207 20988 97259 21040
rect 97207 20924 97259 20976
rect 93458 20551 93510 20603
rect 93522 20551 93574 20603
rect 95673 20505 95725 20557
rect 95673 20441 95725 20493
rect 95673 20377 95725 20429
rect 97197 20499 97249 20551
rect 97197 20435 97249 20487
rect 97197 20371 97249 20423
rect 92131 20146 92183 20198
rect 53519 17120 53571 17172
rect 53519 17056 53571 17108
rect 53519 16992 53571 17044
rect 53519 16928 53571 16980
rect 53519 16864 53571 16916
rect 53519 16800 53571 16852
rect 53519 16736 53571 16788
rect 53519 16672 53571 16724
rect 53519 16608 53571 16660
rect 53519 16544 53571 16596
rect 53519 16480 53571 16532
rect 53519 16416 53571 16468
rect 53519 16352 53571 16404
rect 53519 16288 53571 16340
rect 53519 16224 53571 16276
rect 53519 16160 53571 16212
rect 53519 16096 53571 16148
rect 53519 16032 53571 16084
rect 53519 15968 53571 16020
rect 53519 15904 53571 15956
rect 53519 15840 53571 15892
rect 53519 15776 53571 15828
rect 53519 15712 53571 15764
rect 53519 15648 53571 15700
rect 53519 15584 53571 15636
rect 53519 15520 53571 15572
rect 53519 15456 53571 15508
rect 53519 15392 53571 15444
rect 53519 15328 53571 15380
rect 53519 15264 53571 15316
rect 53519 15200 53571 15252
rect 53519 15136 53571 15188
rect 53519 15072 53571 15124
rect 53519 15008 53571 15060
rect 53519 14944 53571 14996
rect 53519 14880 53571 14932
rect 53519 14816 53571 14868
rect 53519 14752 53571 14804
rect 53519 14688 53571 14740
rect 53519 14624 53571 14676
rect 53519 14560 53571 14612
rect 53519 14496 53571 14548
rect 53519 14432 53571 14484
rect 53519 14368 53571 14420
rect 53519 14304 53571 14356
rect 53519 14240 53571 14292
rect 53519 14176 53571 14228
rect 53519 14112 53571 14164
rect 53519 14048 53571 14100
rect 53519 13984 53571 14036
rect 53519 13920 53571 13972
rect 56525 17113 56577 17165
rect 56525 17049 56577 17101
rect 56525 16985 56577 17037
rect 56525 16921 56577 16973
rect 56525 16857 56577 16909
rect 56525 16793 56577 16845
rect 56525 16729 56577 16781
rect 56525 16665 56577 16717
rect 56525 16601 56577 16653
rect 56525 16537 56577 16589
rect 56525 16473 56577 16525
rect 56525 16409 56577 16461
rect 56525 16345 56577 16397
rect 56525 16281 56577 16333
rect 56525 16217 56577 16269
rect 56525 16153 56577 16205
rect 56525 16089 56577 16141
rect 56525 16025 56577 16077
rect 56525 15961 56577 16013
rect 56525 15897 56577 15949
rect 56525 15833 56577 15885
rect 56525 15769 56577 15821
rect 56525 15705 56577 15757
rect 56525 15641 56577 15693
rect 56525 15577 56577 15629
rect 56525 15513 56577 15565
rect 56525 15449 56577 15501
rect 56525 15385 56577 15437
rect 56525 15321 56577 15373
rect 56525 15257 56577 15309
rect 56525 15193 56577 15245
rect 56525 15129 56577 15181
rect 56525 15065 56577 15117
rect 56525 15001 56577 15053
rect 56525 14937 56577 14989
rect 56525 14873 56577 14925
rect 56525 14809 56577 14861
rect 56525 14745 56577 14797
rect 56525 14681 56577 14733
rect 56525 14617 56577 14669
rect 56525 14553 56577 14605
rect 56525 14489 56577 14541
rect 56525 14425 56577 14477
rect 56525 14361 56577 14413
rect 56525 14297 56577 14349
rect 56525 14233 56577 14285
rect 56525 14169 56577 14221
rect 56525 14105 56577 14157
rect 56525 14041 56577 14093
rect 56525 13977 56577 14029
rect 56525 13913 56577 13965
rect 54943 11732 55123 11912
<< metal2 >>
rect 41684 102152 41920 102172
rect 41684 101936 41694 102152
rect 41910 101936 41920 102152
rect 41684 101916 41920 101936
rect 69700 102123 69936 102143
rect 69700 101907 69710 102123
rect 69926 101907 69936 102123
rect 69700 101887 69936 101907
rect 81750 102124 81986 102144
rect 81750 101908 81760 102124
rect 81976 101908 81986 102124
rect 81750 101888 81986 101908
rect 71238 100765 71366 100777
rect 40245 100740 40346 100755
rect 40245 100710 40269 100740
rect 40321 100710 40346 100740
rect 40245 100654 40267 100710
rect 40323 100654 40346 100710
rect 40245 100630 40269 100654
rect 40321 100630 40346 100654
rect 40245 100574 40267 100630
rect 40323 100574 40346 100630
rect 40245 100560 40269 100574
rect 40321 100560 40346 100574
rect 40245 100550 40346 100560
rect 40245 100494 40267 100550
rect 40323 100494 40346 100550
rect 40245 100484 40346 100494
rect 40245 100470 40269 100484
rect 40321 100470 40346 100484
rect 40245 100414 40267 100470
rect 40323 100414 40346 100470
rect 40245 100390 40269 100414
rect 40321 100390 40346 100414
rect 40245 100334 40267 100390
rect 40323 100334 40346 100390
rect 40245 100310 40269 100334
rect 40321 100310 40346 100334
rect 40245 100254 40267 100310
rect 40323 100254 40346 100310
rect 40245 100240 40269 100254
rect 40321 100240 40346 100254
rect 40245 100230 40346 100240
rect 40245 100174 40267 100230
rect 40323 100174 40346 100230
rect 40245 100164 40346 100174
rect 40245 100150 40269 100164
rect 40321 100150 40346 100164
rect 40245 100094 40267 100150
rect 40323 100094 40346 100150
rect 40245 100070 40269 100094
rect 40321 100070 40346 100094
rect 40245 100014 40267 100070
rect 40323 100014 40346 100070
rect 40245 99990 40269 100014
rect 40321 99990 40346 100014
rect 40245 99934 40267 99990
rect 40323 99934 40346 99990
rect 40245 99920 40269 99934
rect 40321 99920 40346 99934
rect 40245 99910 40346 99920
rect 40245 99854 40267 99910
rect 40323 99854 40346 99910
rect 40245 99844 40346 99854
rect 40245 99830 40269 99844
rect 40321 99830 40346 99844
rect 40245 99774 40267 99830
rect 40323 99774 40346 99830
rect 40245 99750 40269 99774
rect 40321 99750 40346 99774
rect 40245 99694 40267 99750
rect 40323 99694 40346 99750
rect 40245 99670 40269 99694
rect 40321 99670 40346 99694
rect 40245 99614 40267 99670
rect 40323 99614 40346 99670
rect 40245 99600 40269 99614
rect 40321 99600 40346 99614
rect 40245 99590 40346 99600
rect 40245 99534 40267 99590
rect 40323 99534 40346 99590
rect 40245 99524 40346 99534
rect 40245 99510 40269 99524
rect 40321 99510 40346 99524
rect 40245 99454 40267 99510
rect 40323 99454 40346 99510
rect 40245 99430 40269 99454
rect 40321 99430 40346 99454
rect 40245 99374 40267 99430
rect 40323 99374 40346 99430
rect 40245 99350 40269 99374
rect 40321 99350 40346 99374
rect 40245 99294 40267 99350
rect 40323 99294 40346 99350
rect 40245 99280 40269 99294
rect 40321 99280 40346 99294
rect 40245 99270 40346 99280
rect 40245 99214 40267 99270
rect 40323 99214 40346 99270
rect 40245 99204 40346 99214
rect 40245 99190 40269 99204
rect 40321 99190 40346 99204
rect 40245 99134 40267 99190
rect 40323 99134 40346 99190
rect 40245 99110 40269 99134
rect 40321 99110 40346 99134
rect 40245 99054 40267 99110
rect 40323 99054 40346 99110
rect 40245 99030 40269 99054
rect 40321 99030 40346 99054
rect 40245 98974 40267 99030
rect 40323 98974 40346 99030
rect 40245 98960 40269 98974
rect 40321 98960 40346 98974
rect 40245 98950 40346 98960
rect 40245 98894 40267 98950
rect 40323 98894 40346 98950
rect 40245 98884 40346 98894
rect 40245 98870 40269 98884
rect 40321 98870 40346 98884
rect 40245 98814 40267 98870
rect 40323 98814 40346 98870
rect 40245 98790 40269 98814
rect 40321 98790 40346 98814
rect 40245 98734 40267 98790
rect 40323 98734 40346 98790
rect 40245 98710 40269 98734
rect 40321 98710 40346 98734
rect 40245 98654 40267 98710
rect 40323 98654 40346 98710
rect 40245 98640 40269 98654
rect 40321 98640 40346 98654
rect 40245 98630 40346 98640
rect 40245 98574 40267 98630
rect 40323 98574 40346 98630
rect 40245 98564 40346 98574
rect 40245 98550 40269 98564
rect 40321 98550 40346 98564
rect 40245 98494 40267 98550
rect 40323 98494 40346 98550
rect 40245 98470 40269 98494
rect 40321 98470 40346 98494
rect 40245 98414 40267 98470
rect 40323 98414 40346 98470
rect 40245 98390 40269 98414
rect 40321 98390 40346 98414
rect 40245 98334 40267 98390
rect 40323 98334 40346 98390
rect 40245 98320 40269 98334
rect 40321 98320 40346 98334
rect 40245 98310 40346 98320
rect 40245 98254 40267 98310
rect 40323 98254 40346 98310
rect 40245 98244 40346 98254
rect 40245 98230 40269 98244
rect 40321 98230 40346 98244
rect 40245 98174 40267 98230
rect 40323 98174 40346 98230
rect 40245 98150 40269 98174
rect 40321 98150 40346 98174
rect 40245 98094 40267 98150
rect 40323 98094 40346 98150
rect 40245 98070 40269 98094
rect 40321 98070 40346 98094
rect 40245 98014 40267 98070
rect 40323 98014 40346 98070
rect 40245 98000 40269 98014
rect 40321 98000 40346 98014
rect 40245 97990 40346 98000
rect 40245 97934 40267 97990
rect 40323 97934 40346 97990
rect 40245 97924 40346 97934
rect 40245 97910 40269 97924
rect 40321 97910 40346 97924
rect 40245 97854 40267 97910
rect 40323 97854 40346 97910
rect 40245 97830 40269 97854
rect 40321 97830 40346 97854
rect 40245 97774 40267 97830
rect 40323 97774 40346 97830
rect 40245 97750 40269 97774
rect 40321 97750 40346 97774
rect 40245 97694 40267 97750
rect 40323 97694 40346 97750
rect 40245 97680 40269 97694
rect 40321 97680 40346 97694
rect 40245 97670 40346 97680
rect 40245 97614 40267 97670
rect 40323 97614 40346 97670
rect 40245 97604 40346 97614
rect 40245 97590 40269 97604
rect 40321 97590 40346 97604
rect 40245 97534 40267 97590
rect 40323 97534 40346 97590
rect 40245 97510 40269 97534
rect 40321 97510 40346 97534
rect 40245 97454 40267 97510
rect 40323 97454 40346 97510
rect 40245 97424 40269 97454
rect 40321 97424 40346 97454
rect 40245 97410 40346 97424
rect 43246 100746 43347 100761
rect 43246 100716 43270 100746
rect 43322 100716 43347 100746
rect 43246 100660 43268 100716
rect 43324 100660 43347 100716
rect 43246 100636 43270 100660
rect 43322 100636 43347 100660
rect 43246 100580 43268 100636
rect 43324 100580 43347 100636
rect 43246 100566 43270 100580
rect 43322 100566 43347 100580
rect 43246 100556 43347 100566
rect 43246 100500 43268 100556
rect 43324 100500 43347 100556
rect 43246 100490 43347 100500
rect 43246 100476 43270 100490
rect 43322 100476 43347 100490
rect 43246 100420 43268 100476
rect 43324 100420 43347 100476
rect 43246 100396 43270 100420
rect 43322 100396 43347 100420
rect 43246 100340 43268 100396
rect 43324 100340 43347 100396
rect 43246 100316 43270 100340
rect 43322 100316 43347 100340
rect 43246 100260 43268 100316
rect 43324 100260 43347 100316
rect 43246 100246 43270 100260
rect 43322 100246 43347 100260
rect 43246 100236 43347 100246
rect 43246 100180 43268 100236
rect 43324 100180 43347 100236
rect 43246 100170 43347 100180
rect 43246 100156 43270 100170
rect 43322 100156 43347 100170
rect 43246 100100 43268 100156
rect 43324 100100 43347 100156
rect 43246 100076 43270 100100
rect 43322 100076 43347 100100
rect 43246 100020 43268 100076
rect 43324 100020 43347 100076
rect 43246 99996 43270 100020
rect 43322 99996 43347 100020
rect 43246 99940 43268 99996
rect 43324 99940 43347 99996
rect 43246 99926 43270 99940
rect 43322 99926 43347 99940
rect 43246 99916 43347 99926
rect 43246 99860 43268 99916
rect 43324 99860 43347 99916
rect 43246 99850 43347 99860
rect 43246 99836 43270 99850
rect 43322 99836 43347 99850
rect 43246 99780 43268 99836
rect 43324 99780 43347 99836
rect 43246 99756 43270 99780
rect 43322 99756 43347 99780
rect 43246 99700 43268 99756
rect 43324 99700 43347 99756
rect 43246 99676 43270 99700
rect 43322 99676 43347 99700
rect 43246 99620 43268 99676
rect 43324 99620 43347 99676
rect 43246 99606 43270 99620
rect 43322 99606 43347 99620
rect 43246 99596 43347 99606
rect 43246 99540 43268 99596
rect 43324 99540 43347 99596
rect 43246 99530 43347 99540
rect 43246 99516 43270 99530
rect 43322 99516 43347 99530
rect 43246 99460 43268 99516
rect 43324 99460 43347 99516
rect 43246 99436 43270 99460
rect 43322 99436 43347 99460
rect 43246 99380 43268 99436
rect 43324 99380 43347 99436
rect 43246 99356 43270 99380
rect 43322 99356 43347 99380
rect 43246 99300 43268 99356
rect 43324 99300 43347 99356
rect 43246 99286 43270 99300
rect 43322 99286 43347 99300
rect 43246 99276 43347 99286
rect 43246 99220 43268 99276
rect 43324 99220 43347 99276
rect 43246 99210 43347 99220
rect 43246 99196 43270 99210
rect 43322 99196 43347 99210
rect 43246 99140 43268 99196
rect 43324 99140 43347 99196
rect 43246 99116 43270 99140
rect 43322 99116 43347 99140
rect 43246 99060 43268 99116
rect 43324 99060 43347 99116
rect 43246 99036 43270 99060
rect 43322 99036 43347 99060
rect 43246 98980 43268 99036
rect 43324 98980 43347 99036
rect 43246 98966 43270 98980
rect 43322 98966 43347 98980
rect 43246 98956 43347 98966
rect 43246 98900 43268 98956
rect 43324 98900 43347 98956
rect 43246 98890 43347 98900
rect 43246 98876 43270 98890
rect 43322 98876 43347 98890
rect 43246 98820 43268 98876
rect 43324 98820 43347 98876
rect 43246 98796 43270 98820
rect 43322 98796 43347 98820
rect 43246 98740 43268 98796
rect 43324 98740 43347 98796
rect 43246 98716 43270 98740
rect 43322 98716 43347 98740
rect 43246 98660 43268 98716
rect 43324 98660 43347 98716
rect 43246 98646 43270 98660
rect 43322 98646 43347 98660
rect 43246 98636 43347 98646
rect 43246 98580 43268 98636
rect 43324 98580 43347 98636
rect 43246 98570 43347 98580
rect 43246 98556 43270 98570
rect 43322 98556 43347 98570
rect 43246 98500 43268 98556
rect 43324 98500 43347 98556
rect 43246 98476 43270 98500
rect 43322 98476 43347 98500
rect 43246 98420 43268 98476
rect 43324 98420 43347 98476
rect 43246 98396 43270 98420
rect 43322 98396 43347 98420
rect 43246 98340 43268 98396
rect 43324 98340 43347 98396
rect 43246 98326 43270 98340
rect 43322 98326 43347 98340
rect 43246 98316 43347 98326
rect 43246 98260 43268 98316
rect 43324 98260 43347 98316
rect 43246 98250 43347 98260
rect 43246 98236 43270 98250
rect 43322 98236 43347 98250
rect 43246 98180 43268 98236
rect 43324 98180 43347 98236
rect 43246 98156 43270 98180
rect 43322 98156 43347 98180
rect 43246 98100 43268 98156
rect 43324 98100 43347 98156
rect 43246 98076 43270 98100
rect 43322 98076 43347 98100
rect 43246 98020 43268 98076
rect 43324 98020 43347 98076
rect 43246 98006 43270 98020
rect 43322 98006 43347 98020
rect 43246 97996 43347 98006
rect 43246 97940 43268 97996
rect 43324 97940 43347 97996
rect 43246 97930 43347 97940
rect 43246 97916 43270 97930
rect 43322 97916 43347 97930
rect 43246 97860 43268 97916
rect 43324 97860 43347 97916
rect 43246 97836 43270 97860
rect 43322 97836 43347 97860
rect 43246 97780 43268 97836
rect 43324 97780 43347 97836
rect 43246 97756 43270 97780
rect 43322 97756 43347 97780
rect 43246 97700 43268 97756
rect 43324 97700 43347 97756
rect 43246 97686 43270 97700
rect 43322 97686 43347 97700
rect 43246 97676 43347 97686
rect 43246 97620 43268 97676
rect 43324 97620 43347 97676
rect 43246 97610 43347 97620
rect 43246 97596 43270 97610
rect 43322 97596 43347 97610
rect 43246 97540 43268 97596
rect 43324 97540 43347 97596
rect 43246 97516 43270 97540
rect 43322 97516 43347 97540
rect 43246 97460 43268 97516
rect 43324 97460 43347 97516
rect 43246 97430 43270 97460
rect 43322 97430 43347 97460
rect 43246 97416 43347 97430
rect 68237 100752 68365 100764
rect 68237 100742 68273 100752
rect 68329 100742 68365 100752
rect 68237 97426 68243 100742
rect 68359 97426 68365 100742
rect 68237 97416 68273 97426
rect 68329 97416 68365 97426
rect 71238 100755 71274 100765
rect 71330 100755 71366 100765
rect 71238 97439 71244 100755
rect 71360 97439 71366 100755
rect 71238 97429 71274 97439
rect 71330 97429 71366 97439
rect 71238 97417 71366 97429
rect 68237 97404 68365 97416
rect 40430 95820 40494 95834
rect 40430 95764 40434 95820
rect 40490 95764 40494 95820
rect 40430 95750 40494 95764
rect 41608 95816 41672 95830
rect 41608 95760 41612 95816
rect 41668 95760 41672 95816
rect 41608 95746 41672 95760
rect 41825 95823 41889 95837
rect 41825 95767 41829 95823
rect 41885 95767 41889 95823
rect 41825 95753 41889 95767
rect 42959 95820 43023 95834
rect 42959 95764 42963 95820
rect 43019 95764 43023 95820
rect 42959 95750 43023 95764
rect 40540 94316 40604 94330
rect 40540 94260 40544 94316
rect 40600 94260 40604 94316
rect 40540 94246 40604 94260
rect 41654 94302 41718 94316
rect 41654 94246 41658 94302
rect 41714 94246 41718 94302
rect 41654 94232 41718 94246
rect 41867 94303 41931 94317
rect 41867 94247 41871 94303
rect 41927 94247 41931 94303
rect 41867 94233 41931 94247
rect 43031 94303 43095 94317
rect 43031 94247 43035 94303
rect 43091 94247 43095 94303
rect 43031 94233 43095 94247
rect 40386 92721 40450 92735
rect 40386 92665 40390 92721
rect 40446 92665 40450 92721
rect 40386 92651 40450 92665
rect 40395 92357 40447 92651
rect 41672 92516 41736 92547
rect 41672 92510 41678 92516
rect 41730 92510 41736 92516
rect 41672 92454 41676 92510
rect 41732 92454 41736 92510
rect 41672 92452 41736 92454
rect 41672 92430 41678 92452
rect 41730 92430 41736 92452
rect 41672 92374 41676 92430
rect 41732 92374 41736 92430
rect 41672 92350 41678 92374
rect 41730 92350 41736 92374
rect 41672 92294 41676 92350
rect 41732 92294 41736 92350
rect 41131 92273 41204 92293
rect 41131 92217 41139 92273
rect 41195 92217 41204 92273
rect 41131 92211 41141 92217
rect 41193 92211 41204 92217
rect 41131 92199 41204 92211
rect 41131 92193 41141 92199
rect 41193 92193 41204 92199
rect 41131 92137 41139 92193
rect 41195 92137 41204 92193
rect 41672 92272 41678 92294
rect 41730 92272 41736 92294
rect 41672 92270 41736 92272
rect 41672 92214 41676 92270
rect 41732 92214 41736 92270
rect 41672 92208 41678 92214
rect 41730 92208 41736 92214
rect 41672 92178 41736 92208
rect 42215 92276 42288 92296
rect 42215 92220 42223 92276
rect 42279 92220 42288 92276
rect 42215 92214 42225 92220
rect 42277 92214 42288 92220
rect 42215 92202 42288 92214
rect 42215 92196 42225 92202
rect 42277 92196 42288 92202
rect 41131 92117 41204 92137
rect 42215 92140 42223 92196
rect 42279 92140 42288 92196
rect 42215 92120 42288 92140
rect 42902 92105 42954 92409
rect 42895 92091 42959 92105
rect 42895 92035 42899 92091
rect 42955 92035 42959 92091
rect 42895 92021 42959 92035
rect 42902 92018 42954 92021
rect 40517 91631 40581 91645
rect 40517 91575 40521 91631
rect 40577 91575 40581 91631
rect 40517 91561 40581 91575
rect 41672 91625 41736 91639
rect 41672 91569 41676 91625
rect 41732 91569 41736 91625
rect 41672 91555 41736 91569
rect 42790 91636 42854 91650
rect 42790 91580 42794 91636
rect 42850 91580 42854 91636
rect 42790 91566 42854 91580
rect 74524 88760 74590 88775
rect 74524 88746 74531 88760
rect 74583 88746 74590 88760
rect 74524 88690 74529 88746
rect 74585 88690 74590 88746
rect 74524 88666 74531 88690
rect 74583 88666 74590 88690
rect 74524 88610 74529 88666
rect 74585 88610 74590 88666
rect 74524 88586 74531 88610
rect 74583 88586 74590 88610
rect 74524 88530 74529 88586
rect 74585 88530 74590 88586
rect 74524 88516 74531 88530
rect 74583 88516 74590 88530
rect 74524 88506 74590 88516
rect 74524 88450 74529 88506
rect 74585 88450 74590 88506
rect 74524 88440 74590 88450
rect 74524 88426 74531 88440
rect 74583 88426 74590 88440
rect 74524 88370 74529 88426
rect 74585 88370 74590 88426
rect 74524 88346 74531 88370
rect 74583 88346 74590 88370
rect 74524 88290 74529 88346
rect 74585 88290 74590 88346
rect 74524 88266 74531 88290
rect 74583 88266 74590 88290
rect 74524 88210 74529 88266
rect 74585 88210 74590 88266
rect 74524 88196 74531 88210
rect 74583 88196 74590 88210
rect 74524 88181 74590 88196
rect 81052 88760 81118 88775
rect 81052 88746 81059 88760
rect 81111 88746 81118 88760
rect 81052 88690 81057 88746
rect 81113 88690 81118 88746
rect 81052 88666 81059 88690
rect 81111 88666 81118 88690
rect 81052 88610 81057 88666
rect 81113 88610 81118 88666
rect 81052 88586 81059 88610
rect 81111 88586 81118 88610
rect 81052 88530 81057 88586
rect 81113 88530 81118 88586
rect 81052 88516 81059 88530
rect 81111 88516 81118 88530
rect 81052 88506 81118 88516
rect 81052 88450 81057 88506
rect 81113 88450 81118 88506
rect 81052 88440 81118 88450
rect 81052 88426 81059 88440
rect 81111 88426 81118 88440
rect 81052 88370 81057 88426
rect 81113 88370 81118 88426
rect 81052 88346 81059 88370
rect 81111 88346 81118 88370
rect 81052 88290 81057 88346
rect 81113 88290 81118 88346
rect 81052 88266 81059 88290
rect 81111 88266 81118 88290
rect 81052 88210 81057 88266
rect 81113 88210 81118 88266
rect 81052 88196 81059 88210
rect 81111 88196 81118 88210
rect 81052 88181 81118 88196
rect 88668 88760 88734 88775
rect 88668 88746 88675 88760
rect 88727 88746 88734 88760
rect 88668 88690 88673 88746
rect 88729 88690 88734 88746
rect 88668 88666 88675 88690
rect 88727 88666 88734 88690
rect 88668 88610 88673 88666
rect 88729 88610 88734 88666
rect 88668 88586 88675 88610
rect 88727 88586 88734 88610
rect 88668 88530 88673 88586
rect 88729 88530 88734 88586
rect 88668 88516 88675 88530
rect 88727 88516 88734 88530
rect 88668 88506 88734 88516
rect 88668 88450 88673 88506
rect 88729 88450 88734 88506
rect 88668 88440 88734 88450
rect 88668 88426 88675 88440
rect 88727 88426 88734 88440
rect 88668 88370 88673 88426
rect 88729 88370 88734 88426
rect 88668 88346 88675 88370
rect 88727 88346 88734 88370
rect 88668 88290 88673 88346
rect 88729 88290 88734 88346
rect 88668 88266 88675 88290
rect 88727 88266 88734 88290
rect 88668 88210 88673 88266
rect 88729 88210 88734 88266
rect 88668 88196 88675 88210
rect 88727 88196 88734 88210
rect 88668 88181 88734 88196
rect 47210 87420 47652 87434
rect 47210 87418 47243 87420
rect 47299 87418 47323 87420
rect 47379 87418 47403 87420
rect 47459 87418 47483 87420
rect 47539 87418 47563 87420
rect 47619 87418 47652 87420
rect 47210 87366 47213 87418
rect 47393 87366 47403 87418
rect 47459 87366 47469 87418
rect 47649 87366 47652 87418
rect 47210 87364 47243 87366
rect 47299 87364 47323 87366
rect 47379 87364 47403 87366
rect 47459 87364 47483 87366
rect 47539 87364 47563 87366
rect 47619 87364 47652 87366
rect 47210 87350 47652 87364
rect 49021 87422 49463 87436
rect 49021 87420 49054 87422
rect 49110 87420 49134 87422
rect 49190 87420 49214 87422
rect 49270 87420 49294 87422
rect 49350 87420 49374 87422
rect 49430 87420 49463 87422
rect 49021 87368 49024 87420
rect 49204 87368 49214 87420
rect 49270 87368 49280 87420
rect 49460 87368 49463 87420
rect 49021 87366 49054 87368
rect 49110 87366 49134 87368
rect 49190 87366 49214 87368
rect 49270 87366 49294 87368
rect 49350 87366 49374 87368
rect 49430 87366 49463 87368
rect 49021 87352 49463 87366
rect 50816 87418 51258 87432
rect 50816 87416 50849 87418
rect 50905 87416 50929 87418
rect 50985 87416 51009 87418
rect 51065 87416 51089 87418
rect 51145 87416 51169 87418
rect 51225 87416 51258 87418
rect 50816 87364 50819 87416
rect 50999 87364 51009 87416
rect 51065 87364 51075 87416
rect 51255 87364 51258 87416
rect 50816 87362 50849 87364
rect 50905 87362 50929 87364
rect 50985 87362 51009 87364
rect 51065 87362 51089 87364
rect 51145 87362 51169 87364
rect 51225 87362 51258 87364
rect 50816 87348 51258 87362
rect 52615 87416 53057 87430
rect 52615 87414 52648 87416
rect 52704 87414 52728 87416
rect 52784 87414 52808 87416
rect 52864 87414 52888 87416
rect 52944 87414 52968 87416
rect 53024 87414 53057 87416
rect 52615 87362 52618 87414
rect 52798 87362 52808 87414
rect 52864 87362 52874 87414
rect 53054 87362 53057 87414
rect 52615 87360 52648 87362
rect 52704 87360 52728 87362
rect 52784 87360 52808 87362
rect 52864 87360 52888 87362
rect 52944 87360 52968 87362
rect 53024 87360 53057 87362
rect 52615 87346 53057 87360
rect 54406 87420 54848 87434
rect 54406 87418 54439 87420
rect 54495 87418 54519 87420
rect 54575 87418 54599 87420
rect 54655 87418 54679 87420
rect 54735 87418 54759 87420
rect 54815 87418 54848 87420
rect 54406 87366 54409 87418
rect 54589 87366 54599 87418
rect 54655 87366 54665 87418
rect 54845 87366 54848 87418
rect 54406 87364 54439 87366
rect 54495 87364 54519 87366
rect 54575 87364 54599 87366
rect 54655 87364 54679 87366
rect 54735 87364 54759 87366
rect 54815 87364 54848 87366
rect 54406 87350 54848 87364
rect 56208 87416 56650 87430
rect 56208 87414 56241 87416
rect 56297 87414 56321 87416
rect 56377 87414 56401 87416
rect 56457 87414 56481 87416
rect 56537 87414 56561 87416
rect 56617 87414 56650 87416
rect 56208 87362 56211 87414
rect 56391 87362 56401 87414
rect 56457 87362 56467 87414
rect 56647 87362 56650 87414
rect 56208 87360 56241 87362
rect 56297 87360 56321 87362
rect 56377 87360 56401 87362
rect 56457 87360 56481 87362
rect 56537 87360 56561 87362
rect 56617 87360 56650 87362
rect 56208 87346 56650 87360
rect 57851 87242 58381 87264
rect 50155 87216 50395 87238
rect 50155 87000 50167 87216
rect 50383 87000 50395 87216
rect 57851 87224 57888 87242
rect 58344 87224 58381 87242
rect 57851 87044 57866 87224
rect 58366 87044 58381 87224
rect 57851 87026 57888 87044
rect 58344 87026 58381 87044
rect 57851 87004 58381 87026
rect 50155 86978 50395 87000
rect 75069 86757 75135 86772
rect 75069 86743 75076 86757
rect 75128 86743 75135 86757
rect 75069 86687 75074 86743
rect 75130 86687 75135 86743
rect 75069 86663 75076 86687
rect 75128 86663 75135 86687
rect 75069 86607 75074 86663
rect 75130 86607 75135 86663
rect 75069 86583 75076 86607
rect 75128 86583 75135 86607
rect 75069 86527 75074 86583
rect 75130 86527 75135 86583
rect 75069 86513 75076 86527
rect 75128 86513 75135 86527
rect 75069 86503 75135 86513
rect 75069 86447 75074 86503
rect 75130 86447 75135 86503
rect 75069 86437 75135 86447
rect 75069 86423 75076 86437
rect 75128 86423 75135 86437
rect 75069 86367 75074 86423
rect 75130 86367 75135 86423
rect 75069 86343 75076 86367
rect 75128 86343 75135 86367
rect 75069 86287 75074 86343
rect 75130 86287 75135 86343
rect 75069 86263 75076 86287
rect 75128 86263 75135 86287
rect 75069 86207 75074 86263
rect 75130 86207 75135 86263
rect 75069 86193 75076 86207
rect 75128 86193 75135 86207
rect 75069 86178 75135 86193
rect 76157 86757 76223 86772
rect 76157 86743 76164 86757
rect 76216 86743 76223 86757
rect 76157 86687 76162 86743
rect 76218 86687 76223 86743
rect 76157 86663 76164 86687
rect 76216 86663 76223 86687
rect 76157 86607 76162 86663
rect 76218 86607 76223 86663
rect 76157 86583 76164 86607
rect 76216 86583 76223 86607
rect 76157 86527 76162 86583
rect 76218 86527 76223 86583
rect 76157 86513 76164 86527
rect 76216 86513 76223 86527
rect 76157 86503 76223 86513
rect 76157 86447 76162 86503
rect 76218 86447 76223 86503
rect 76157 86437 76223 86447
rect 76157 86423 76164 86437
rect 76216 86423 76223 86437
rect 76157 86367 76162 86423
rect 76218 86367 76223 86423
rect 76157 86343 76164 86367
rect 76216 86343 76223 86367
rect 76157 86287 76162 86343
rect 76218 86287 76223 86343
rect 76157 86263 76164 86287
rect 76216 86263 76223 86287
rect 76157 86207 76162 86263
rect 76218 86207 76223 86263
rect 76157 86193 76164 86207
rect 76216 86193 76223 86207
rect 76157 86178 76223 86193
rect 78333 86757 78399 86772
rect 78333 86743 78340 86757
rect 78392 86743 78399 86757
rect 78333 86687 78338 86743
rect 78394 86687 78399 86743
rect 78333 86663 78340 86687
rect 78392 86663 78399 86687
rect 78333 86607 78338 86663
rect 78394 86607 78399 86663
rect 78333 86583 78340 86607
rect 78392 86583 78399 86607
rect 78333 86527 78338 86583
rect 78394 86527 78399 86583
rect 78333 86513 78340 86527
rect 78392 86513 78399 86527
rect 78333 86503 78399 86513
rect 78333 86447 78338 86503
rect 78394 86447 78399 86503
rect 78333 86437 78399 86447
rect 78333 86423 78340 86437
rect 78392 86423 78399 86437
rect 78333 86367 78338 86423
rect 78394 86367 78399 86423
rect 78333 86343 78340 86367
rect 78392 86343 78399 86367
rect 78333 86287 78338 86343
rect 78394 86287 78399 86343
rect 78333 86263 78340 86287
rect 78392 86263 78399 86287
rect 78333 86207 78338 86263
rect 78394 86207 78399 86263
rect 78333 86193 78340 86207
rect 78392 86193 78399 86207
rect 78333 86178 78399 86193
rect 79421 86757 79487 86772
rect 79421 86743 79428 86757
rect 79480 86743 79487 86757
rect 79421 86687 79426 86743
rect 79482 86687 79487 86743
rect 79421 86663 79428 86687
rect 79480 86663 79487 86687
rect 79421 86607 79426 86663
rect 79482 86607 79487 86663
rect 79421 86583 79428 86607
rect 79480 86583 79487 86607
rect 79421 86527 79426 86583
rect 79482 86527 79487 86583
rect 79421 86513 79428 86527
rect 79480 86513 79487 86527
rect 79421 86503 79487 86513
rect 79421 86447 79426 86503
rect 79482 86447 79487 86503
rect 79421 86437 79487 86447
rect 79421 86423 79428 86437
rect 79480 86423 79487 86437
rect 79421 86367 79426 86423
rect 79482 86367 79487 86423
rect 79421 86343 79428 86367
rect 79480 86343 79487 86367
rect 79421 86287 79426 86343
rect 79482 86287 79487 86343
rect 79421 86263 79428 86287
rect 79480 86263 79487 86287
rect 79421 86207 79426 86263
rect 79482 86207 79487 86263
rect 79421 86193 79428 86207
rect 79480 86193 79487 86207
rect 79421 86178 79487 86193
rect 80509 86757 80575 86772
rect 80509 86743 80516 86757
rect 80568 86743 80575 86757
rect 80509 86687 80514 86743
rect 80570 86687 80575 86743
rect 80509 86663 80516 86687
rect 80568 86663 80575 86687
rect 80509 86607 80514 86663
rect 80570 86607 80575 86663
rect 80509 86583 80516 86607
rect 80568 86583 80575 86607
rect 80509 86527 80514 86583
rect 80570 86527 80575 86583
rect 80509 86513 80516 86527
rect 80568 86513 80575 86527
rect 80509 86503 80575 86513
rect 80509 86447 80514 86503
rect 80570 86447 80575 86503
rect 80509 86437 80575 86447
rect 80509 86423 80516 86437
rect 80568 86423 80575 86437
rect 80509 86367 80514 86423
rect 80570 86367 80575 86423
rect 80509 86343 80516 86367
rect 80568 86343 80575 86367
rect 80509 86287 80514 86343
rect 80570 86287 80575 86343
rect 80509 86263 80516 86287
rect 80568 86263 80575 86287
rect 80509 86207 80514 86263
rect 80570 86207 80575 86263
rect 80509 86193 80516 86207
rect 80568 86193 80575 86207
rect 80509 86178 80575 86193
rect 81597 86757 81663 86772
rect 81597 86743 81604 86757
rect 81656 86743 81663 86757
rect 81597 86687 81602 86743
rect 81658 86687 81663 86743
rect 81597 86663 81604 86687
rect 81656 86663 81663 86687
rect 81597 86607 81602 86663
rect 81658 86607 81663 86663
rect 81597 86583 81604 86607
rect 81656 86583 81663 86607
rect 81597 86527 81602 86583
rect 81658 86527 81663 86583
rect 81597 86513 81604 86527
rect 81656 86513 81663 86527
rect 81597 86503 81663 86513
rect 81597 86447 81602 86503
rect 81658 86447 81663 86503
rect 81597 86437 81663 86447
rect 81597 86423 81604 86437
rect 81656 86423 81663 86437
rect 81597 86367 81602 86423
rect 81658 86367 81663 86423
rect 81597 86343 81604 86367
rect 81656 86343 81663 86367
rect 81597 86287 81602 86343
rect 81658 86287 81663 86343
rect 81597 86263 81604 86287
rect 81656 86263 81663 86287
rect 81597 86207 81602 86263
rect 81658 86207 81663 86263
rect 81597 86193 81604 86207
rect 81656 86193 81663 86207
rect 81597 86178 81663 86193
rect 82685 86757 82751 86772
rect 82685 86743 82692 86757
rect 82744 86743 82751 86757
rect 82685 86687 82690 86743
rect 82746 86687 82751 86743
rect 82685 86663 82692 86687
rect 82744 86663 82751 86687
rect 82685 86607 82690 86663
rect 82746 86607 82751 86663
rect 82685 86583 82692 86607
rect 82744 86583 82751 86607
rect 82685 86527 82690 86583
rect 82746 86527 82751 86583
rect 82685 86513 82692 86527
rect 82744 86513 82751 86527
rect 82685 86503 82751 86513
rect 82685 86447 82690 86503
rect 82746 86447 82751 86503
rect 82685 86437 82751 86447
rect 82685 86423 82692 86437
rect 82744 86423 82751 86437
rect 82685 86367 82690 86423
rect 82746 86367 82751 86423
rect 82685 86343 82692 86367
rect 82744 86343 82751 86367
rect 82685 86287 82690 86343
rect 82746 86287 82751 86343
rect 82685 86263 82692 86287
rect 82744 86263 82751 86287
rect 82685 86207 82690 86263
rect 82746 86207 82751 86263
rect 82685 86193 82692 86207
rect 82744 86193 82751 86207
rect 82685 86178 82751 86193
rect 83773 86757 83839 86772
rect 83773 86743 83780 86757
rect 83832 86743 83839 86757
rect 83773 86687 83778 86743
rect 83834 86687 83839 86743
rect 83773 86663 83780 86687
rect 83832 86663 83839 86687
rect 83773 86607 83778 86663
rect 83834 86607 83839 86663
rect 83773 86583 83780 86607
rect 83832 86583 83839 86607
rect 83773 86527 83778 86583
rect 83834 86527 83839 86583
rect 83773 86513 83780 86527
rect 83832 86513 83839 86527
rect 83773 86503 83839 86513
rect 83773 86447 83778 86503
rect 83834 86447 83839 86503
rect 83773 86437 83839 86447
rect 83773 86423 83780 86437
rect 83832 86423 83839 86437
rect 83773 86367 83778 86423
rect 83834 86367 83839 86423
rect 83773 86343 83780 86367
rect 83832 86343 83839 86367
rect 83773 86287 83778 86343
rect 83834 86287 83839 86343
rect 83773 86263 83780 86287
rect 83832 86263 83839 86287
rect 83773 86207 83778 86263
rect 83834 86207 83839 86263
rect 83773 86193 83780 86207
rect 83832 86193 83839 86207
rect 83773 86178 83839 86193
rect 85949 86757 86015 86772
rect 85949 86743 85956 86757
rect 86008 86743 86015 86757
rect 85949 86687 85954 86743
rect 86010 86687 86015 86743
rect 85949 86663 85956 86687
rect 86008 86663 86015 86687
rect 85949 86607 85954 86663
rect 86010 86607 86015 86663
rect 85949 86583 85956 86607
rect 86008 86583 86015 86607
rect 85949 86527 85954 86583
rect 86010 86527 86015 86583
rect 85949 86513 85956 86527
rect 86008 86513 86015 86527
rect 85949 86503 86015 86513
rect 85949 86447 85954 86503
rect 86010 86447 86015 86503
rect 85949 86437 86015 86447
rect 85949 86423 85956 86437
rect 86008 86423 86015 86437
rect 85949 86367 85954 86423
rect 86010 86367 86015 86423
rect 85949 86343 85956 86367
rect 86008 86343 86015 86367
rect 85949 86287 85954 86343
rect 86010 86287 86015 86343
rect 85949 86263 85956 86287
rect 86008 86263 86015 86287
rect 85949 86207 85954 86263
rect 86010 86207 86015 86263
rect 85949 86193 85956 86207
rect 86008 86193 86015 86207
rect 85949 86178 86015 86193
rect 87037 86757 87103 86772
rect 87037 86743 87044 86757
rect 87096 86743 87103 86757
rect 87037 86687 87042 86743
rect 87098 86687 87103 86743
rect 87037 86663 87044 86687
rect 87096 86663 87103 86687
rect 87037 86607 87042 86663
rect 87098 86607 87103 86663
rect 87037 86583 87044 86607
rect 87096 86583 87103 86607
rect 87037 86527 87042 86583
rect 87098 86527 87103 86583
rect 87037 86513 87044 86527
rect 87096 86513 87103 86527
rect 87037 86503 87103 86513
rect 87037 86447 87042 86503
rect 87098 86447 87103 86503
rect 87037 86437 87103 86447
rect 87037 86423 87044 86437
rect 87096 86423 87103 86437
rect 87037 86367 87042 86423
rect 87098 86367 87103 86423
rect 87037 86343 87044 86367
rect 87096 86343 87103 86367
rect 87037 86287 87042 86343
rect 87098 86287 87103 86343
rect 87037 86263 87044 86287
rect 87096 86263 87103 86287
rect 87037 86207 87042 86263
rect 87098 86207 87103 86263
rect 87037 86193 87044 86207
rect 87096 86193 87103 86207
rect 87037 86178 87103 86193
rect 88125 86757 88191 86772
rect 88125 86743 88132 86757
rect 88184 86743 88191 86757
rect 88125 86687 88130 86743
rect 88186 86687 88191 86743
rect 88125 86663 88132 86687
rect 88184 86663 88191 86687
rect 88125 86607 88130 86663
rect 88186 86607 88191 86663
rect 88125 86583 88132 86607
rect 88184 86583 88191 86607
rect 88125 86527 88130 86583
rect 88186 86527 88191 86583
rect 88125 86513 88132 86527
rect 88184 86513 88191 86527
rect 88125 86503 88191 86513
rect 88125 86447 88130 86503
rect 88186 86447 88191 86503
rect 88125 86437 88191 86447
rect 88125 86423 88132 86437
rect 88184 86423 88191 86437
rect 88125 86367 88130 86423
rect 88186 86367 88191 86423
rect 88125 86343 88132 86367
rect 88184 86343 88191 86367
rect 88125 86287 88130 86343
rect 88186 86287 88191 86343
rect 88125 86263 88132 86287
rect 88184 86263 88191 86287
rect 88125 86207 88130 86263
rect 88186 86207 88191 86263
rect 88125 86193 88132 86207
rect 88184 86193 88191 86207
rect 88125 86178 88191 86193
rect 57441 84830 57613 84859
rect 57441 84824 57469 84830
rect 57585 84824 57613 84830
rect 48537 78613 48601 78627
rect 48537 78557 48541 78613
rect 48597 78557 48601 78613
rect 48537 78543 48601 78557
rect 50228 78614 50292 78628
rect 50228 78558 50232 78614
rect 50288 78558 50292 78614
rect 50228 78544 50292 78558
rect 51933 78613 51997 78627
rect 51933 78557 51937 78613
rect 51993 78557 51997 78613
rect 51933 78543 51997 78557
rect 53729 78613 53793 78627
rect 53729 78557 53733 78613
rect 53789 78557 53793 78613
rect 53729 78543 53793 78557
rect 55558 78613 55622 78627
rect 55558 78557 55562 78613
rect 55618 78557 55622 78613
rect 55558 78543 55622 78557
rect 47390 78421 47632 78435
rect 47390 78365 47403 78421
rect 47459 78419 47483 78421
rect 47539 78419 47563 78421
rect 47473 78367 47483 78419
rect 47539 78367 47549 78419
rect 47459 78365 47483 78367
rect 47539 78365 47563 78367
rect 47619 78365 47632 78421
rect 47390 78351 47632 78365
rect 49185 78420 49427 78434
rect 49185 78364 49198 78420
rect 49254 78418 49278 78420
rect 49334 78418 49358 78420
rect 49268 78366 49278 78418
rect 49334 78366 49344 78418
rect 49254 78364 49278 78366
rect 49334 78364 49358 78366
rect 49414 78364 49427 78420
rect 49185 78350 49427 78364
rect 50985 78422 51227 78436
rect 50985 78366 50998 78422
rect 51054 78420 51078 78422
rect 51134 78420 51158 78422
rect 51068 78368 51078 78420
rect 51134 78368 51144 78420
rect 51054 78366 51078 78368
rect 51134 78366 51158 78368
rect 51214 78366 51227 78422
rect 50985 78352 51227 78366
rect 52783 78421 53025 78435
rect 52783 78365 52796 78421
rect 52852 78419 52876 78421
rect 52932 78419 52956 78421
rect 52866 78367 52876 78419
rect 52932 78367 52942 78419
rect 52852 78365 52876 78367
rect 52932 78365 52956 78367
rect 53012 78365 53025 78421
rect 52783 78351 53025 78365
rect 54581 78422 54823 78436
rect 54581 78366 54594 78422
rect 54650 78420 54674 78422
rect 54730 78420 54754 78422
rect 54664 78368 54674 78420
rect 54730 78368 54740 78420
rect 54650 78366 54674 78368
rect 54730 78366 54754 78368
rect 54810 78366 54823 78422
rect 54581 78352 54823 78366
rect 56384 78421 56626 78435
rect 56384 78365 56397 78421
rect 56453 78419 56477 78421
rect 56533 78419 56557 78421
rect 56467 78367 56477 78419
rect 56533 78367 56543 78419
rect 56453 78365 56477 78367
rect 56533 78365 56557 78367
rect 56613 78365 56626 78421
rect 56384 78351 56626 78365
rect 57270 78422 57334 78436
rect 57270 78366 57274 78422
rect 57330 78366 57334 78422
rect 57270 78352 57334 78366
rect 42311 77622 42439 77632
rect 49544 77622 49608 77632
rect 42311 77616 49608 77622
rect 42311 77564 42317 77616
rect 42369 77564 42381 77616
rect 42433 77564 49550 77616
rect 49602 77564 49608 77616
rect 42311 77558 49608 77564
rect 42311 77548 42439 77558
rect 49544 77548 49608 77558
rect 50105 77616 50233 77632
rect 50105 77564 50111 77616
rect 50163 77564 50175 77616
rect 50227 77564 50233 77616
rect 47696 77008 47824 77024
rect 47696 76956 47702 77008
rect 47754 76956 47766 77008
rect 47818 76956 47824 77008
rect 47696 74953 47824 76956
rect 48240 75261 48324 75281
rect 48240 75205 48254 75261
rect 48310 75205 48324 75261
rect 48240 75191 48256 75205
rect 48308 75191 48324 75205
rect 49372 75265 49436 75279
rect 49372 75209 49376 75265
rect 49432 75209 49436 75265
rect 49372 75195 49436 75209
rect 48240 75181 48324 75191
rect 48240 75125 48254 75181
rect 48310 75125 48324 75181
rect 48240 75115 48324 75125
rect 48240 75101 48256 75115
rect 48308 75101 48324 75115
rect 48240 75045 48254 75101
rect 48310 75045 48324 75101
rect 48240 75026 48324 75045
rect 47696 74901 47702 74953
rect 47754 74901 47766 74953
rect 47818 74901 47824 74953
rect 30024 73738 30368 73752
rect 30024 73736 30048 73738
rect 30104 73736 30128 73738
rect 30184 73736 30208 73738
rect 30264 73736 30288 73738
rect 30344 73736 30368 73738
rect 30024 73684 30042 73736
rect 30104 73684 30106 73736
rect 30286 73684 30288 73736
rect 30350 73684 30368 73736
rect 30024 73682 30048 73684
rect 30104 73682 30128 73684
rect 30184 73682 30208 73684
rect 30264 73682 30288 73684
rect 30344 73682 30368 73684
rect 30024 73668 30368 73682
rect 30686 73431 30937 73445
rect 30686 73429 30703 73431
rect 30759 73429 30783 73431
rect 30839 73429 30863 73431
rect 30919 73429 30937 73431
rect 30686 73377 30689 73429
rect 30933 73377 30937 73429
rect 30686 73375 30703 73377
rect 30759 73375 30783 73377
rect 30839 73375 30863 73377
rect 30919 73375 30937 73377
rect 30686 73361 30937 73375
rect 31034 73442 31098 73456
rect 31034 73386 31038 73442
rect 31094 73386 31098 73442
rect 31034 73372 31098 73386
rect 31110 73196 31454 73210
rect 31110 73194 31134 73196
rect 31190 73194 31214 73196
rect 31270 73194 31294 73196
rect 31350 73194 31374 73196
rect 31430 73194 31454 73196
rect 31110 73142 31128 73194
rect 31190 73142 31192 73194
rect 31372 73142 31374 73194
rect 31436 73142 31454 73194
rect 31110 73140 31134 73142
rect 31190 73140 31214 73142
rect 31270 73140 31294 73142
rect 31350 73140 31374 73142
rect 31430 73140 31454 73142
rect 31110 73126 31454 73140
rect 30007 67318 30104 67345
rect 30007 67296 30029 67318
rect 30081 67296 30104 67318
rect 30007 67240 30027 67296
rect 30083 67240 30104 67296
rect 30007 67216 30029 67240
rect 30081 67216 30104 67240
rect 30007 67160 30027 67216
rect 30083 67160 30104 67216
rect 30007 67138 30029 67160
rect 30081 67138 30104 67160
rect 30007 67136 30104 67138
rect 30007 67080 30027 67136
rect 30083 67080 30104 67136
rect 30007 67074 30029 67080
rect 30081 67074 30104 67080
rect 30007 67062 30104 67074
rect 30007 67056 30029 67062
rect 30081 67056 30104 67062
rect 30007 67000 30027 67056
rect 30083 67000 30104 67056
rect 43625 67079 43689 67093
rect 43625 67023 43629 67079
rect 43685 67023 43689 67079
rect 43625 67009 43689 67023
rect 30007 66998 30104 67000
rect 30007 66976 30029 66998
rect 30081 66976 30104 66998
rect 30007 66920 30027 66976
rect 30083 66920 30104 66976
rect 30007 66896 30029 66920
rect 30081 66896 30104 66920
rect 30007 66840 30027 66896
rect 30083 66840 30104 66896
rect 30007 66818 30029 66840
rect 30081 66818 30104 66840
rect 30007 66791 30104 66818
rect 44401 66416 44465 66430
rect 44401 66360 44405 66416
rect 44461 66360 44465 66416
rect 44401 66346 44465 66360
rect 30012 66177 30099 66201
rect 30012 66155 30029 66177
rect 30081 66155 30099 66177
rect 30012 66099 30027 66155
rect 30083 66099 30099 66155
rect 35619 66181 35683 66195
rect 35619 66125 35623 66181
rect 35679 66125 35683 66181
rect 35619 66111 35683 66125
rect 30012 66075 30029 66099
rect 30081 66075 30099 66099
rect 30012 66019 30027 66075
rect 30083 66019 30099 66075
rect 30012 65997 30029 66019
rect 30081 65997 30099 66019
rect 30012 65995 30099 65997
rect 30012 65939 30027 65995
rect 30083 65939 30099 65995
rect 30012 65933 30029 65939
rect 30081 65933 30099 65939
rect 30012 65921 30099 65933
rect 30012 65915 30029 65921
rect 30081 65915 30099 65921
rect 30012 65859 30027 65915
rect 30083 65859 30099 65915
rect 30012 65857 30099 65859
rect 30012 65835 30029 65857
rect 30081 65835 30099 65857
rect 30012 65779 30027 65835
rect 30083 65779 30099 65835
rect 30012 65755 30029 65779
rect 30081 65755 30099 65779
rect 30012 65699 30027 65755
rect 30083 65699 30099 65755
rect 30012 65677 30029 65699
rect 30081 65677 30099 65699
rect 30012 65675 30099 65677
rect 30012 65619 30027 65675
rect 30083 65619 30099 65675
rect 30012 65613 30029 65619
rect 30081 65613 30099 65619
rect 30012 65601 30099 65613
rect 30012 65595 30029 65601
rect 30081 65595 30099 65601
rect 30012 65539 30027 65595
rect 30083 65539 30099 65595
rect 30012 65537 30099 65539
rect 30012 65515 30029 65537
rect 30081 65515 30099 65537
rect 30012 65459 30027 65515
rect 30083 65459 30099 65515
rect 30012 65435 30029 65459
rect 30081 65435 30099 65459
rect 30012 65379 30027 65435
rect 30083 65379 30099 65435
rect 30012 65357 30029 65379
rect 30081 65357 30099 65379
rect 30012 65355 30099 65357
rect 30012 65299 30027 65355
rect 30083 65299 30099 65355
rect 30012 65293 30029 65299
rect 30081 65293 30099 65299
rect 30012 65281 30099 65293
rect 30012 65275 30029 65281
rect 30081 65275 30099 65281
rect 30012 65219 30027 65275
rect 30083 65219 30099 65275
rect 30012 65217 30099 65219
rect 30012 65195 30029 65217
rect 30081 65195 30099 65217
rect 30012 65139 30027 65195
rect 30083 65139 30099 65195
rect 30012 65115 30029 65139
rect 30081 65115 30099 65139
rect 30012 65059 30027 65115
rect 30083 65059 30099 65115
rect 30012 65037 30029 65059
rect 30081 65037 30099 65059
rect 30012 65014 30099 65037
rect 30017 64651 30104 64675
rect 30017 64629 30034 64651
rect 30086 64629 30104 64651
rect 30017 64573 30032 64629
rect 30088 64573 30104 64629
rect 30017 64549 30034 64573
rect 30086 64549 30104 64573
rect 30017 64493 30032 64549
rect 30088 64493 30104 64549
rect 30017 64471 30034 64493
rect 30086 64471 30104 64493
rect 30017 64469 30104 64471
rect 30017 64413 30032 64469
rect 30088 64413 30104 64469
rect 30017 64407 30034 64413
rect 30086 64407 30104 64413
rect 30017 64395 30104 64407
rect 30017 64389 30034 64395
rect 30086 64389 30104 64395
rect 30017 64333 30032 64389
rect 30088 64333 30104 64389
rect 30017 64331 30104 64333
rect 30017 64309 30034 64331
rect 30086 64309 30104 64331
rect 30017 64253 30032 64309
rect 30088 64253 30104 64309
rect 30017 64229 30034 64253
rect 30086 64229 30104 64253
rect 30017 64173 30032 64229
rect 30088 64173 30104 64229
rect 30017 64151 30034 64173
rect 30086 64151 30104 64173
rect 30017 64149 30104 64151
rect 30017 64093 30032 64149
rect 30088 64093 30104 64149
rect 30017 64087 30034 64093
rect 30086 64087 30104 64093
rect 30017 64075 30104 64087
rect 30017 64069 30034 64075
rect 30086 64069 30104 64075
rect 30017 64013 30032 64069
rect 30088 64013 30104 64069
rect 30017 64011 30104 64013
rect 30017 63989 30034 64011
rect 30086 63989 30104 64011
rect 30017 63933 30032 63989
rect 30088 63933 30104 63989
rect 30017 63909 30034 63933
rect 30086 63909 30104 63933
rect 30017 63853 30032 63909
rect 30088 63853 30104 63909
rect 30017 63831 30034 63853
rect 30086 63831 30104 63853
rect 30017 63829 30104 63831
rect 30017 63773 30032 63829
rect 30088 63773 30104 63829
rect 30017 63767 30034 63773
rect 30086 63767 30104 63773
rect 30017 63755 30104 63767
rect 30017 63749 30034 63755
rect 30086 63749 30104 63755
rect 47696 63821 47824 74901
rect 50105 74951 50233 77564
rect 57441 77168 57459 84824
rect 57595 77168 57613 84824
rect 57441 77162 57469 77168
rect 57585 77162 57613 77168
rect 57441 77133 57613 77162
rect 67271 84836 67645 84868
rect 67271 84834 67310 84836
rect 67606 84834 67645 84836
rect 50105 74899 50111 74951
rect 50163 74899 50175 74951
rect 50227 74899 50233 74951
rect 48220 74794 48314 74823
rect 48220 74738 48239 74794
rect 48295 74738 48314 74794
rect 48220 74728 48314 74738
rect 48220 74714 48241 74728
rect 48293 74714 48314 74728
rect 48220 74658 48239 74714
rect 48295 74658 48314 74714
rect 48220 74634 48241 74658
rect 48293 74634 48314 74658
rect 48220 74578 48239 74634
rect 48295 74578 48314 74634
rect 48220 74554 48241 74578
rect 48293 74554 48314 74578
rect 48220 74498 48239 74554
rect 48295 74498 48314 74554
rect 48220 74484 48241 74498
rect 48293 74484 48314 74498
rect 48220 74474 48314 74484
rect 48220 74418 48239 74474
rect 48295 74418 48314 74474
rect 48220 74390 48314 74418
rect 48614 74459 48678 74473
rect 48614 74403 48618 74459
rect 48674 74403 48678 74459
rect 48614 74389 48678 74403
rect 47696 63769 47702 63821
rect 47754 63769 47766 63821
rect 47818 63769 47824 63821
rect 47696 63750 47824 63769
rect 50105 63821 50233 74899
rect 51406 75086 53206 75098
rect 51406 74906 51416 75086
rect 53196 74906 53206 75086
rect 53732 75075 54558 75106
rect 53732 75065 53757 75075
rect 54533 75065 54558 75075
rect 53732 74949 53735 75065
rect 54555 74949 54558 75065
rect 53732 74939 53757 74949
rect 54533 74939 54558 74949
rect 53732 74908 54558 74939
rect 55439 75065 56329 75096
rect 55439 75055 55456 75065
rect 56312 75055 56329 75065
rect 55439 74939 55442 75055
rect 56326 74939 56329 75055
rect 55439 74929 55456 74939
rect 56312 74929 56329 74939
rect 51406 74895 53206 74906
rect 55439 74898 56329 74929
rect 57016 74793 57215 74806
rect 57016 74783 57047 74793
rect 57183 74783 57215 74793
rect 51162 74738 51346 74752
rect 51162 74736 51186 74738
rect 51322 74736 51346 74738
rect 51162 71804 51164 74736
rect 51344 71804 51346 74736
rect 51162 71802 51186 71804
rect 51322 71802 51346 71804
rect 51162 71788 51346 71802
rect 57016 71787 57025 74783
rect 57205 71787 57215 74783
rect 57016 71777 57047 71787
rect 57183 71777 57215 71787
rect 57016 71764 57215 71777
rect 67271 71662 67272 84834
rect 67644 71662 67645 84834
rect 74524 84760 74590 84775
rect 74524 84746 74531 84760
rect 74583 84746 74590 84760
rect 74524 84690 74529 84746
rect 74585 84690 74590 84746
rect 74524 84666 74531 84690
rect 74583 84666 74590 84690
rect 74524 84610 74529 84666
rect 74585 84610 74590 84666
rect 74524 84586 74531 84610
rect 74583 84586 74590 84610
rect 74524 84530 74529 84586
rect 74585 84530 74590 84586
rect 74524 84516 74531 84530
rect 74583 84516 74590 84530
rect 74524 84506 74590 84516
rect 74524 84450 74529 84506
rect 74585 84450 74590 84506
rect 74524 84440 74590 84450
rect 74524 84426 74531 84440
rect 74583 84426 74590 84440
rect 74524 84370 74529 84426
rect 74585 84370 74590 84426
rect 74524 84346 74531 84370
rect 74583 84346 74590 84370
rect 74524 84290 74529 84346
rect 74585 84290 74590 84346
rect 74524 84266 74531 84290
rect 74583 84266 74590 84290
rect 74524 84210 74529 84266
rect 74585 84210 74590 84266
rect 74524 84196 74531 84210
rect 74583 84196 74590 84210
rect 74524 84181 74590 84196
rect 75612 84760 75678 84775
rect 75612 84746 75619 84760
rect 75671 84746 75678 84760
rect 75612 84690 75617 84746
rect 75673 84690 75678 84746
rect 75612 84666 75619 84690
rect 75671 84666 75678 84690
rect 75612 84610 75617 84666
rect 75673 84610 75678 84666
rect 75612 84586 75619 84610
rect 75671 84586 75678 84610
rect 75612 84530 75617 84586
rect 75673 84530 75678 84586
rect 75612 84516 75619 84530
rect 75671 84516 75678 84530
rect 75612 84506 75678 84516
rect 75612 84450 75617 84506
rect 75673 84450 75678 84506
rect 75612 84440 75678 84450
rect 75612 84426 75619 84440
rect 75671 84426 75678 84440
rect 75612 84370 75617 84426
rect 75673 84370 75678 84426
rect 75612 84346 75619 84370
rect 75671 84346 75678 84370
rect 75612 84290 75617 84346
rect 75673 84290 75678 84346
rect 75612 84266 75619 84290
rect 75671 84266 75678 84290
rect 75612 84210 75617 84266
rect 75673 84210 75678 84266
rect 75612 84196 75619 84210
rect 75671 84196 75678 84210
rect 75612 84181 75678 84196
rect 76700 84760 76766 84775
rect 76700 84746 76707 84760
rect 76759 84746 76766 84760
rect 76700 84690 76705 84746
rect 76761 84690 76766 84746
rect 76700 84666 76707 84690
rect 76759 84666 76766 84690
rect 76700 84610 76705 84666
rect 76761 84610 76766 84666
rect 76700 84586 76707 84610
rect 76759 84586 76766 84610
rect 76700 84530 76705 84586
rect 76761 84530 76766 84586
rect 76700 84516 76707 84530
rect 76759 84516 76766 84530
rect 76700 84506 76766 84516
rect 76700 84450 76705 84506
rect 76761 84450 76766 84506
rect 76700 84440 76766 84450
rect 76700 84426 76707 84440
rect 76759 84426 76766 84440
rect 76700 84370 76705 84426
rect 76761 84370 76766 84426
rect 76700 84346 76707 84370
rect 76759 84346 76766 84370
rect 76700 84290 76705 84346
rect 76761 84290 76766 84346
rect 76700 84266 76707 84290
rect 76759 84266 76766 84290
rect 76700 84210 76705 84266
rect 76761 84210 76766 84266
rect 76700 84196 76707 84210
rect 76759 84196 76766 84210
rect 76700 84181 76766 84196
rect 77788 84760 77854 84775
rect 77788 84746 77795 84760
rect 77847 84746 77854 84760
rect 77788 84690 77793 84746
rect 77849 84690 77854 84746
rect 77788 84666 77795 84690
rect 77847 84666 77854 84690
rect 77788 84610 77793 84666
rect 77849 84610 77854 84666
rect 77788 84586 77795 84610
rect 77847 84586 77854 84610
rect 77788 84530 77793 84586
rect 77849 84530 77854 84586
rect 77788 84516 77795 84530
rect 77847 84516 77854 84530
rect 77788 84506 77854 84516
rect 77788 84450 77793 84506
rect 77849 84450 77854 84506
rect 77788 84440 77854 84450
rect 77788 84426 77795 84440
rect 77847 84426 77854 84440
rect 77788 84370 77793 84426
rect 77849 84370 77854 84426
rect 77788 84346 77795 84370
rect 77847 84346 77854 84370
rect 77788 84290 77793 84346
rect 77849 84290 77854 84346
rect 77788 84266 77795 84290
rect 77847 84266 77854 84290
rect 77788 84210 77793 84266
rect 77849 84210 77854 84266
rect 77788 84196 77795 84210
rect 77847 84196 77854 84210
rect 77788 84181 77854 84196
rect 78876 84760 78942 84775
rect 78876 84746 78883 84760
rect 78935 84746 78942 84760
rect 78876 84690 78881 84746
rect 78937 84690 78942 84746
rect 78876 84666 78883 84690
rect 78935 84666 78942 84690
rect 78876 84610 78881 84666
rect 78937 84610 78942 84666
rect 78876 84586 78883 84610
rect 78935 84586 78942 84610
rect 78876 84530 78881 84586
rect 78937 84530 78942 84586
rect 78876 84516 78883 84530
rect 78935 84516 78942 84530
rect 78876 84506 78942 84516
rect 78876 84450 78881 84506
rect 78937 84450 78942 84506
rect 78876 84440 78942 84450
rect 78876 84426 78883 84440
rect 78935 84426 78942 84440
rect 78876 84370 78881 84426
rect 78937 84370 78942 84426
rect 78876 84346 78883 84370
rect 78935 84346 78942 84370
rect 78876 84290 78881 84346
rect 78937 84290 78942 84346
rect 78876 84266 78883 84290
rect 78935 84266 78942 84290
rect 78876 84210 78881 84266
rect 78937 84210 78942 84266
rect 78876 84196 78883 84210
rect 78935 84196 78942 84210
rect 78876 84181 78942 84196
rect 79964 84760 80030 84775
rect 79964 84746 79971 84760
rect 80023 84746 80030 84760
rect 79964 84690 79969 84746
rect 80025 84690 80030 84746
rect 79964 84666 79971 84690
rect 80023 84666 80030 84690
rect 79964 84610 79969 84666
rect 80025 84610 80030 84666
rect 79964 84586 79971 84610
rect 80023 84586 80030 84610
rect 79964 84530 79969 84586
rect 80025 84530 80030 84586
rect 79964 84516 79971 84530
rect 80023 84516 80030 84530
rect 79964 84506 80030 84516
rect 79964 84450 79969 84506
rect 80025 84450 80030 84506
rect 79964 84440 80030 84450
rect 79964 84426 79971 84440
rect 80023 84426 80030 84440
rect 79964 84370 79969 84426
rect 80025 84370 80030 84426
rect 79964 84346 79971 84370
rect 80023 84346 80030 84370
rect 79964 84290 79969 84346
rect 80025 84290 80030 84346
rect 79964 84266 79971 84290
rect 80023 84266 80030 84290
rect 79964 84210 79969 84266
rect 80025 84210 80030 84266
rect 79964 84196 79971 84210
rect 80023 84196 80030 84210
rect 79964 84181 80030 84196
rect 81052 84760 81118 84775
rect 81052 84746 81059 84760
rect 81111 84746 81118 84760
rect 81052 84690 81057 84746
rect 81113 84690 81118 84746
rect 81052 84666 81059 84690
rect 81111 84666 81118 84690
rect 81052 84610 81057 84666
rect 81113 84610 81118 84666
rect 81052 84586 81059 84610
rect 81111 84586 81118 84610
rect 81052 84530 81057 84586
rect 81113 84530 81118 84586
rect 81052 84516 81059 84530
rect 81111 84516 81118 84530
rect 81052 84506 81118 84516
rect 81052 84450 81057 84506
rect 81113 84450 81118 84506
rect 81052 84440 81118 84450
rect 81052 84426 81059 84440
rect 81111 84426 81118 84440
rect 81052 84370 81057 84426
rect 81113 84370 81118 84426
rect 81052 84346 81059 84370
rect 81111 84346 81118 84370
rect 81052 84290 81057 84346
rect 81113 84290 81118 84346
rect 81052 84266 81059 84290
rect 81111 84266 81118 84290
rect 81052 84210 81057 84266
rect 81113 84210 81118 84266
rect 81052 84196 81059 84210
rect 81111 84196 81118 84210
rect 81052 84181 81118 84196
rect 82140 84760 82206 84775
rect 82140 84746 82147 84760
rect 82199 84746 82206 84760
rect 82140 84690 82145 84746
rect 82201 84690 82206 84746
rect 82140 84666 82147 84690
rect 82199 84666 82206 84690
rect 82140 84610 82145 84666
rect 82201 84610 82206 84666
rect 82140 84586 82147 84610
rect 82199 84586 82206 84610
rect 82140 84530 82145 84586
rect 82201 84530 82206 84586
rect 82140 84516 82147 84530
rect 82199 84516 82206 84530
rect 82140 84506 82206 84516
rect 82140 84450 82145 84506
rect 82201 84450 82206 84506
rect 82140 84440 82206 84450
rect 82140 84426 82147 84440
rect 82199 84426 82206 84440
rect 82140 84370 82145 84426
rect 82201 84370 82206 84426
rect 82140 84346 82147 84370
rect 82199 84346 82206 84370
rect 82140 84290 82145 84346
rect 82201 84290 82206 84346
rect 82140 84266 82147 84290
rect 82199 84266 82206 84290
rect 82140 84210 82145 84266
rect 82201 84210 82206 84266
rect 82140 84196 82147 84210
rect 82199 84196 82206 84210
rect 82140 84181 82206 84196
rect 83228 84760 83294 84775
rect 83228 84746 83235 84760
rect 83287 84746 83294 84760
rect 83228 84690 83233 84746
rect 83289 84690 83294 84746
rect 83228 84666 83235 84690
rect 83287 84666 83294 84690
rect 83228 84610 83233 84666
rect 83289 84610 83294 84666
rect 83228 84586 83235 84610
rect 83287 84586 83294 84610
rect 83228 84530 83233 84586
rect 83289 84530 83294 84586
rect 83228 84516 83235 84530
rect 83287 84516 83294 84530
rect 83228 84506 83294 84516
rect 83228 84450 83233 84506
rect 83289 84450 83294 84506
rect 83228 84440 83294 84450
rect 83228 84426 83235 84440
rect 83287 84426 83294 84440
rect 83228 84370 83233 84426
rect 83289 84370 83294 84426
rect 83228 84346 83235 84370
rect 83287 84346 83294 84370
rect 83228 84290 83233 84346
rect 83289 84290 83294 84346
rect 83228 84266 83235 84290
rect 83287 84266 83294 84290
rect 83228 84210 83233 84266
rect 83289 84210 83294 84266
rect 83228 84196 83235 84210
rect 83287 84196 83294 84210
rect 83228 84181 83294 84196
rect 84316 84760 84382 84775
rect 84316 84746 84323 84760
rect 84375 84746 84382 84760
rect 84316 84690 84321 84746
rect 84377 84690 84382 84746
rect 84316 84666 84323 84690
rect 84375 84666 84382 84690
rect 84316 84610 84321 84666
rect 84377 84610 84382 84666
rect 84316 84586 84323 84610
rect 84375 84586 84382 84610
rect 84316 84530 84321 84586
rect 84377 84530 84382 84586
rect 84316 84516 84323 84530
rect 84375 84516 84382 84530
rect 84316 84506 84382 84516
rect 84316 84450 84321 84506
rect 84377 84450 84382 84506
rect 84316 84440 84382 84450
rect 84316 84426 84323 84440
rect 84375 84426 84382 84440
rect 84316 84370 84321 84426
rect 84377 84370 84382 84426
rect 84316 84346 84323 84370
rect 84375 84346 84382 84370
rect 84316 84290 84321 84346
rect 84377 84290 84382 84346
rect 84316 84266 84323 84290
rect 84375 84266 84382 84290
rect 84316 84210 84321 84266
rect 84377 84210 84382 84266
rect 84316 84196 84323 84210
rect 84375 84196 84382 84210
rect 84316 84181 84382 84196
rect 85404 84760 85470 84775
rect 85404 84746 85411 84760
rect 85463 84746 85470 84760
rect 85404 84690 85409 84746
rect 85465 84690 85470 84746
rect 85404 84666 85411 84690
rect 85463 84666 85470 84690
rect 85404 84610 85409 84666
rect 85465 84610 85470 84666
rect 85404 84586 85411 84610
rect 85463 84586 85470 84610
rect 85404 84530 85409 84586
rect 85465 84530 85470 84586
rect 85404 84516 85411 84530
rect 85463 84516 85470 84530
rect 85404 84506 85470 84516
rect 85404 84450 85409 84506
rect 85465 84450 85470 84506
rect 85404 84440 85470 84450
rect 85404 84426 85411 84440
rect 85463 84426 85470 84440
rect 85404 84370 85409 84426
rect 85465 84370 85470 84426
rect 85404 84346 85411 84370
rect 85463 84346 85470 84370
rect 85404 84290 85409 84346
rect 85465 84290 85470 84346
rect 85404 84266 85411 84290
rect 85463 84266 85470 84290
rect 85404 84210 85409 84266
rect 85465 84210 85470 84266
rect 85404 84196 85411 84210
rect 85463 84196 85470 84210
rect 85404 84181 85470 84196
rect 86492 84760 86558 84775
rect 86492 84746 86499 84760
rect 86551 84746 86558 84760
rect 86492 84690 86497 84746
rect 86553 84690 86558 84746
rect 86492 84666 86499 84690
rect 86551 84666 86558 84690
rect 86492 84610 86497 84666
rect 86553 84610 86558 84666
rect 86492 84586 86499 84610
rect 86551 84586 86558 84610
rect 86492 84530 86497 84586
rect 86553 84530 86558 84586
rect 86492 84516 86499 84530
rect 86551 84516 86558 84530
rect 86492 84506 86558 84516
rect 86492 84450 86497 84506
rect 86553 84450 86558 84506
rect 86492 84440 86558 84450
rect 86492 84426 86499 84440
rect 86551 84426 86558 84440
rect 86492 84370 86497 84426
rect 86553 84370 86558 84426
rect 86492 84346 86499 84370
rect 86551 84346 86558 84370
rect 86492 84290 86497 84346
rect 86553 84290 86558 84346
rect 86492 84266 86499 84290
rect 86551 84266 86558 84290
rect 86492 84210 86497 84266
rect 86553 84210 86558 84266
rect 86492 84196 86499 84210
rect 86551 84196 86558 84210
rect 86492 84181 86558 84196
rect 87580 84760 87646 84775
rect 87580 84746 87587 84760
rect 87639 84746 87646 84760
rect 87580 84690 87585 84746
rect 87641 84690 87646 84746
rect 87580 84666 87587 84690
rect 87639 84666 87646 84690
rect 87580 84610 87585 84666
rect 87641 84610 87646 84666
rect 87580 84586 87587 84610
rect 87639 84586 87646 84610
rect 87580 84530 87585 84586
rect 87641 84530 87646 84586
rect 87580 84516 87587 84530
rect 87639 84516 87646 84530
rect 87580 84506 87646 84516
rect 87580 84450 87585 84506
rect 87641 84450 87646 84506
rect 87580 84440 87646 84450
rect 87580 84426 87587 84440
rect 87639 84426 87646 84440
rect 87580 84370 87585 84426
rect 87641 84370 87646 84426
rect 87580 84346 87587 84370
rect 87639 84346 87646 84370
rect 87580 84290 87585 84346
rect 87641 84290 87646 84346
rect 87580 84266 87587 84290
rect 87639 84266 87646 84290
rect 87580 84210 87585 84266
rect 87641 84210 87646 84266
rect 87580 84196 87587 84210
rect 87639 84196 87646 84210
rect 87580 84181 87646 84196
rect 88668 84760 88734 84775
rect 88668 84746 88675 84760
rect 88727 84746 88734 84760
rect 88668 84690 88673 84746
rect 88729 84690 88734 84746
rect 88668 84666 88675 84690
rect 88727 84666 88734 84690
rect 88668 84610 88673 84666
rect 88729 84610 88734 84666
rect 88668 84586 88675 84610
rect 88727 84586 88734 84610
rect 88668 84530 88673 84586
rect 88729 84530 88734 84586
rect 88668 84516 88675 84530
rect 88727 84516 88734 84530
rect 88668 84506 88734 84516
rect 88668 84450 88673 84506
rect 88729 84450 88734 84506
rect 88668 84440 88734 84450
rect 88668 84426 88675 84440
rect 88727 84426 88734 84440
rect 88668 84370 88673 84426
rect 88729 84370 88734 84426
rect 88668 84346 88675 84370
rect 88727 84346 88734 84370
rect 88668 84290 88673 84346
rect 88729 84290 88734 84346
rect 88668 84266 88675 84290
rect 88727 84266 88734 84290
rect 88668 84210 88673 84266
rect 88729 84210 88734 84266
rect 88668 84196 88675 84210
rect 88727 84196 88734 84210
rect 88668 84181 88734 84196
rect 75069 82757 75135 82772
rect 75069 82743 75076 82757
rect 75128 82743 75135 82757
rect 75069 82687 75074 82743
rect 75130 82687 75135 82743
rect 75069 82663 75076 82687
rect 75128 82663 75135 82687
rect 75069 82607 75074 82663
rect 75130 82607 75135 82663
rect 75069 82583 75076 82607
rect 75128 82583 75135 82607
rect 75069 82527 75074 82583
rect 75130 82527 75135 82583
rect 75069 82513 75076 82527
rect 75128 82513 75135 82527
rect 75069 82503 75135 82513
rect 75069 82447 75074 82503
rect 75130 82447 75135 82503
rect 75069 82437 75135 82447
rect 75069 82423 75076 82437
rect 75128 82423 75135 82437
rect 75069 82367 75074 82423
rect 75130 82367 75135 82423
rect 75069 82343 75076 82367
rect 75128 82343 75135 82367
rect 75069 82287 75074 82343
rect 75130 82287 75135 82343
rect 75069 82263 75076 82287
rect 75128 82263 75135 82287
rect 75069 82207 75074 82263
rect 75130 82207 75135 82263
rect 75069 82193 75076 82207
rect 75128 82193 75135 82207
rect 75069 82178 75135 82193
rect 76157 82757 76223 82772
rect 76157 82743 76164 82757
rect 76216 82743 76223 82757
rect 76157 82687 76162 82743
rect 76218 82687 76223 82743
rect 76157 82663 76164 82687
rect 76216 82663 76223 82687
rect 76157 82607 76162 82663
rect 76218 82607 76223 82663
rect 76157 82583 76164 82607
rect 76216 82583 76223 82607
rect 76157 82527 76162 82583
rect 76218 82527 76223 82583
rect 76157 82513 76164 82527
rect 76216 82513 76223 82527
rect 76157 82503 76223 82513
rect 76157 82447 76162 82503
rect 76218 82447 76223 82503
rect 76157 82437 76223 82447
rect 76157 82423 76164 82437
rect 76216 82423 76223 82437
rect 76157 82367 76162 82423
rect 76218 82367 76223 82423
rect 76157 82343 76164 82367
rect 76216 82343 76223 82367
rect 76157 82287 76162 82343
rect 76218 82287 76223 82343
rect 76157 82263 76164 82287
rect 76216 82263 76223 82287
rect 76157 82207 76162 82263
rect 76218 82207 76223 82263
rect 76157 82193 76164 82207
rect 76216 82193 76223 82207
rect 76157 82178 76223 82193
rect 77245 82757 77311 82772
rect 77245 82743 77252 82757
rect 77304 82743 77311 82757
rect 77245 82687 77250 82743
rect 77306 82687 77311 82743
rect 77245 82663 77252 82687
rect 77304 82663 77311 82687
rect 77245 82607 77250 82663
rect 77306 82607 77311 82663
rect 77245 82583 77252 82607
rect 77304 82583 77311 82607
rect 77245 82527 77250 82583
rect 77306 82527 77311 82583
rect 77245 82513 77252 82527
rect 77304 82513 77311 82527
rect 77245 82503 77311 82513
rect 77245 82447 77250 82503
rect 77306 82447 77311 82503
rect 77245 82437 77311 82447
rect 77245 82423 77252 82437
rect 77304 82423 77311 82437
rect 77245 82367 77250 82423
rect 77306 82367 77311 82423
rect 77245 82343 77252 82367
rect 77304 82343 77311 82367
rect 77245 82287 77250 82343
rect 77306 82287 77311 82343
rect 77245 82263 77252 82287
rect 77304 82263 77311 82287
rect 77245 82207 77250 82263
rect 77306 82207 77311 82263
rect 77245 82193 77252 82207
rect 77304 82193 77311 82207
rect 77245 82178 77311 82193
rect 78333 82757 78399 82772
rect 78333 82743 78340 82757
rect 78392 82743 78399 82757
rect 78333 82687 78338 82743
rect 78394 82687 78399 82743
rect 78333 82663 78340 82687
rect 78392 82663 78399 82687
rect 78333 82607 78338 82663
rect 78394 82607 78399 82663
rect 78333 82583 78340 82607
rect 78392 82583 78399 82607
rect 78333 82527 78338 82583
rect 78394 82527 78399 82583
rect 78333 82513 78340 82527
rect 78392 82513 78399 82527
rect 78333 82503 78399 82513
rect 78333 82447 78338 82503
rect 78394 82447 78399 82503
rect 78333 82437 78399 82447
rect 78333 82423 78340 82437
rect 78392 82423 78399 82437
rect 78333 82367 78338 82423
rect 78394 82367 78399 82423
rect 78333 82343 78340 82367
rect 78392 82343 78399 82367
rect 78333 82287 78338 82343
rect 78394 82287 78399 82343
rect 78333 82263 78340 82287
rect 78392 82263 78399 82287
rect 78333 82207 78338 82263
rect 78394 82207 78399 82263
rect 78333 82193 78340 82207
rect 78392 82193 78399 82207
rect 78333 82178 78399 82193
rect 79421 82757 79487 82772
rect 79421 82743 79428 82757
rect 79480 82743 79487 82757
rect 79421 82687 79426 82743
rect 79482 82687 79487 82743
rect 79421 82663 79428 82687
rect 79480 82663 79487 82687
rect 79421 82607 79426 82663
rect 79482 82607 79487 82663
rect 79421 82583 79428 82607
rect 79480 82583 79487 82607
rect 79421 82527 79426 82583
rect 79482 82527 79487 82583
rect 79421 82513 79428 82527
rect 79480 82513 79487 82527
rect 79421 82503 79487 82513
rect 79421 82447 79426 82503
rect 79482 82447 79487 82503
rect 79421 82437 79487 82447
rect 79421 82423 79428 82437
rect 79480 82423 79487 82437
rect 79421 82367 79426 82423
rect 79482 82367 79487 82423
rect 79421 82343 79428 82367
rect 79480 82343 79487 82367
rect 79421 82287 79426 82343
rect 79482 82287 79487 82343
rect 79421 82263 79428 82287
rect 79480 82263 79487 82287
rect 79421 82207 79426 82263
rect 79482 82207 79487 82263
rect 79421 82193 79428 82207
rect 79480 82193 79487 82207
rect 79421 82178 79487 82193
rect 80509 82757 80575 82772
rect 80509 82743 80516 82757
rect 80568 82743 80575 82757
rect 80509 82687 80514 82743
rect 80570 82687 80575 82743
rect 80509 82663 80516 82687
rect 80568 82663 80575 82687
rect 80509 82607 80514 82663
rect 80570 82607 80575 82663
rect 80509 82583 80516 82607
rect 80568 82583 80575 82607
rect 80509 82527 80514 82583
rect 80570 82527 80575 82583
rect 80509 82513 80516 82527
rect 80568 82513 80575 82527
rect 80509 82503 80575 82513
rect 80509 82447 80514 82503
rect 80570 82447 80575 82503
rect 80509 82437 80575 82447
rect 80509 82423 80516 82437
rect 80568 82423 80575 82437
rect 80509 82367 80514 82423
rect 80570 82367 80575 82423
rect 80509 82343 80516 82367
rect 80568 82343 80575 82367
rect 80509 82287 80514 82343
rect 80570 82287 80575 82343
rect 80509 82263 80516 82287
rect 80568 82263 80575 82287
rect 80509 82207 80514 82263
rect 80570 82207 80575 82263
rect 80509 82193 80516 82207
rect 80568 82193 80575 82207
rect 80509 82178 80575 82193
rect 81597 82757 81663 82772
rect 81597 82743 81604 82757
rect 81656 82743 81663 82757
rect 81597 82687 81602 82743
rect 81658 82687 81663 82743
rect 81597 82663 81604 82687
rect 81656 82663 81663 82687
rect 81597 82607 81602 82663
rect 81658 82607 81663 82663
rect 81597 82583 81604 82607
rect 81656 82583 81663 82607
rect 81597 82527 81602 82583
rect 81658 82527 81663 82583
rect 81597 82513 81604 82527
rect 81656 82513 81663 82527
rect 81597 82503 81663 82513
rect 81597 82447 81602 82503
rect 81658 82447 81663 82503
rect 81597 82437 81663 82447
rect 81597 82423 81604 82437
rect 81656 82423 81663 82437
rect 81597 82367 81602 82423
rect 81658 82367 81663 82423
rect 81597 82343 81604 82367
rect 81656 82343 81663 82367
rect 81597 82287 81602 82343
rect 81658 82287 81663 82343
rect 81597 82263 81604 82287
rect 81656 82263 81663 82287
rect 81597 82207 81602 82263
rect 81658 82207 81663 82263
rect 81597 82193 81604 82207
rect 81656 82193 81663 82207
rect 81597 82178 81663 82193
rect 82685 82757 82751 82772
rect 82685 82743 82692 82757
rect 82744 82743 82751 82757
rect 82685 82687 82690 82743
rect 82746 82687 82751 82743
rect 82685 82663 82692 82687
rect 82744 82663 82751 82687
rect 82685 82607 82690 82663
rect 82746 82607 82751 82663
rect 82685 82583 82692 82607
rect 82744 82583 82751 82607
rect 82685 82527 82690 82583
rect 82746 82527 82751 82583
rect 82685 82513 82692 82527
rect 82744 82513 82751 82527
rect 82685 82503 82751 82513
rect 82685 82447 82690 82503
rect 82746 82447 82751 82503
rect 82685 82437 82751 82447
rect 82685 82423 82692 82437
rect 82744 82423 82751 82437
rect 82685 82367 82690 82423
rect 82746 82367 82751 82423
rect 82685 82343 82692 82367
rect 82744 82343 82751 82367
rect 82685 82287 82690 82343
rect 82746 82287 82751 82343
rect 82685 82263 82692 82287
rect 82744 82263 82751 82287
rect 82685 82207 82690 82263
rect 82746 82207 82751 82263
rect 82685 82193 82692 82207
rect 82744 82193 82751 82207
rect 82685 82178 82751 82193
rect 83773 82757 83839 82772
rect 83773 82743 83780 82757
rect 83832 82743 83839 82757
rect 83773 82687 83778 82743
rect 83834 82687 83839 82743
rect 83773 82663 83780 82687
rect 83832 82663 83839 82687
rect 83773 82607 83778 82663
rect 83834 82607 83839 82663
rect 83773 82583 83780 82607
rect 83832 82583 83839 82607
rect 83773 82527 83778 82583
rect 83834 82527 83839 82583
rect 83773 82513 83780 82527
rect 83832 82513 83839 82527
rect 83773 82503 83839 82513
rect 83773 82447 83778 82503
rect 83834 82447 83839 82503
rect 83773 82437 83839 82447
rect 83773 82423 83780 82437
rect 83832 82423 83839 82437
rect 83773 82367 83778 82423
rect 83834 82367 83839 82423
rect 83773 82343 83780 82367
rect 83832 82343 83839 82367
rect 83773 82287 83778 82343
rect 83834 82287 83839 82343
rect 83773 82263 83780 82287
rect 83832 82263 83839 82287
rect 83773 82207 83778 82263
rect 83834 82207 83839 82263
rect 83773 82193 83780 82207
rect 83832 82193 83839 82207
rect 83773 82178 83839 82193
rect 84861 82757 84927 82772
rect 84861 82743 84868 82757
rect 84920 82743 84927 82757
rect 84861 82687 84866 82743
rect 84922 82687 84927 82743
rect 84861 82663 84868 82687
rect 84920 82663 84927 82687
rect 84861 82607 84866 82663
rect 84922 82607 84927 82663
rect 84861 82583 84868 82607
rect 84920 82583 84927 82607
rect 84861 82527 84866 82583
rect 84922 82527 84927 82583
rect 84861 82513 84868 82527
rect 84920 82513 84927 82527
rect 84861 82503 84927 82513
rect 84861 82447 84866 82503
rect 84922 82447 84927 82503
rect 84861 82437 84927 82447
rect 84861 82423 84868 82437
rect 84920 82423 84927 82437
rect 84861 82367 84866 82423
rect 84922 82367 84927 82423
rect 84861 82343 84868 82367
rect 84920 82343 84927 82367
rect 84861 82287 84866 82343
rect 84922 82287 84927 82343
rect 84861 82263 84868 82287
rect 84920 82263 84927 82287
rect 84861 82207 84866 82263
rect 84922 82207 84927 82263
rect 84861 82193 84868 82207
rect 84920 82193 84927 82207
rect 84861 82178 84927 82193
rect 85949 82757 86015 82772
rect 85949 82743 85956 82757
rect 86008 82743 86015 82757
rect 85949 82687 85954 82743
rect 86010 82687 86015 82743
rect 85949 82663 85956 82687
rect 86008 82663 86015 82687
rect 85949 82607 85954 82663
rect 86010 82607 86015 82663
rect 85949 82583 85956 82607
rect 86008 82583 86015 82607
rect 85949 82527 85954 82583
rect 86010 82527 86015 82583
rect 85949 82513 85956 82527
rect 86008 82513 86015 82527
rect 85949 82503 86015 82513
rect 85949 82447 85954 82503
rect 86010 82447 86015 82503
rect 85949 82437 86015 82447
rect 85949 82423 85956 82437
rect 86008 82423 86015 82437
rect 85949 82367 85954 82423
rect 86010 82367 86015 82423
rect 85949 82343 85956 82367
rect 86008 82343 86015 82367
rect 85949 82287 85954 82343
rect 86010 82287 86015 82343
rect 85949 82263 85956 82287
rect 86008 82263 86015 82287
rect 85949 82207 85954 82263
rect 86010 82207 86015 82263
rect 85949 82193 85956 82207
rect 86008 82193 86015 82207
rect 85949 82178 86015 82193
rect 87037 82757 87103 82772
rect 87037 82743 87044 82757
rect 87096 82743 87103 82757
rect 87037 82687 87042 82743
rect 87098 82687 87103 82743
rect 87037 82663 87044 82687
rect 87096 82663 87103 82687
rect 87037 82607 87042 82663
rect 87098 82607 87103 82663
rect 87037 82583 87044 82607
rect 87096 82583 87103 82607
rect 87037 82527 87042 82583
rect 87098 82527 87103 82583
rect 87037 82513 87044 82527
rect 87096 82513 87103 82527
rect 87037 82503 87103 82513
rect 87037 82447 87042 82503
rect 87098 82447 87103 82503
rect 87037 82437 87103 82447
rect 87037 82423 87044 82437
rect 87096 82423 87103 82437
rect 87037 82367 87042 82423
rect 87098 82367 87103 82423
rect 87037 82343 87044 82367
rect 87096 82343 87103 82367
rect 87037 82287 87042 82343
rect 87098 82287 87103 82343
rect 87037 82263 87044 82287
rect 87096 82263 87103 82287
rect 87037 82207 87042 82263
rect 87098 82207 87103 82263
rect 87037 82193 87044 82207
rect 87096 82193 87103 82207
rect 87037 82178 87103 82193
rect 88125 82757 88191 82772
rect 88125 82743 88132 82757
rect 88184 82743 88191 82757
rect 88125 82687 88130 82743
rect 88186 82687 88191 82743
rect 88125 82663 88132 82687
rect 88184 82663 88191 82687
rect 88125 82607 88130 82663
rect 88186 82607 88191 82663
rect 88125 82583 88132 82607
rect 88184 82583 88191 82607
rect 88125 82527 88130 82583
rect 88186 82527 88191 82583
rect 88125 82513 88132 82527
rect 88184 82513 88191 82527
rect 88125 82503 88191 82513
rect 88125 82447 88130 82503
rect 88186 82447 88191 82503
rect 88125 82437 88191 82447
rect 88125 82423 88132 82437
rect 88184 82423 88191 82437
rect 88125 82367 88130 82423
rect 88186 82367 88191 82423
rect 88125 82343 88132 82367
rect 88184 82343 88191 82367
rect 88125 82287 88130 82343
rect 88186 82287 88191 82343
rect 88125 82263 88132 82287
rect 88184 82263 88191 82287
rect 88125 82207 88130 82263
rect 88186 82207 88191 82263
rect 88125 82193 88132 82207
rect 88184 82193 88191 82207
rect 88125 82178 88191 82193
rect 74524 80760 74590 80775
rect 74524 80746 74531 80760
rect 74583 80746 74590 80760
rect 74524 80690 74529 80746
rect 74585 80690 74590 80746
rect 74524 80666 74531 80690
rect 74583 80666 74590 80690
rect 74524 80610 74529 80666
rect 74585 80610 74590 80666
rect 74524 80586 74531 80610
rect 74583 80586 74590 80610
rect 74524 80530 74529 80586
rect 74585 80530 74590 80586
rect 74524 80516 74531 80530
rect 74583 80516 74590 80530
rect 74524 80506 74590 80516
rect 74524 80450 74529 80506
rect 74585 80450 74590 80506
rect 74524 80440 74590 80450
rect 74524 80426 74531 80440
rect 74583 80426 74590 80440
rect 74524 80370 74529 80426
rect 74585 80370 74590 80426
rect 74524 80346 74531 80370
rect 74583 80346 74590 80370
rect 74524 80290 74529 80346
rect 74585 80290 74590 80346
rect 74524 80266 74531 80290
rect 74583 80266 74590 80290
rect 74524 80210 74529 80266
rect 74585 80210 74590 80266
rect 74524 80196 74531 80210
rect 74583 80196 74590 80210
rect 74524 80181 74590 80196
rect 75612 80760 75678 80775
rect 75612 80746 75619 80760
rect 75671 80746 75678 80760
rect 75612 80690 75617 80746
rect 75673 80690 75678 80746
rect 75612 80666 75619 80690
rect 75671 80666 75678 80690
rect 75612 80610 75617 80666
rect 75673 80610 75678 80666
rect 75612 80586 75619 80610
rect 75671 80586 75678 80610
rect 75612 80530 75617 80586
rect 75673 80530 75678 80586
rect 75612 80516 75619 80530
rect 75671 80516 75678 80530
rect 75612 80506 75678 80516
rect 75612 80450 75617 80506
rect 75673 80450 75678 80506
rect 75612 80440 75678 80450
rect 75612 80426 75619 80440
rect 75671 80426 75678 80440
rect 75612 80370 75617 80426
rect 75673 80370 75678 80426
rect 75612 80346 75619 80370
rect 75671 80346 75678 80370
rect 75612 80290 75617 80346
rect 75673 80290 75678 80346
rect 75612 80266 75619 80290
rect 75671 80266 75678 80290
rect 75612 80210 75617 80266
rect 75673 80210 75678 80266
rect 75612 80196 75619 80210
rect 75671 80196 75678 80210
rect 75612 80181 75678 80196
rect 76700 80760 76766 80775
rect 76700 80746 76707 80760
rect 76759 80746 76766 80760
rect 76700 80690 76705 80746
rect 76761 80690 76766 80746
rect 76700 80666 76707 80690
rect 76759 80666 76766 80690
rect 76700 80610 76705 80666
rect 76761 80610 76766 80666
rect 76700 80586 76707 80610
rect 76759 80586 76766 80610
rect 76700 80530 76705 80586
rect 76761 80530 76766 80586
rect 76700 80516 76707 80530
rect 76759 80516 76766 80530
rect 76700 80506 76766 80516
rect 76700 80450 76705 80506
rect 76761 80450 76766 80506
rect 76700 80440 76766 80450
rect 76700 80426 76707 80440
rect 76759 80426 76766 80440
rect 76700 80370 76705 80426
rect 76761 80370 76766 80426
rect 76700 80346 76707 80370
rect 76759 80346 76766 80370
rect 76700 80290 76705 80346
rect 76761 80290 76766 80346
rect 76700 80266 76707 80290
rect 76759 80266 76766 80290
rect 76700 80210 76705 80266
rect 76761 80210 76766 80266
rect 76700 80196 76707 80210
rect 76759 80196 76766 80210
rect 76700 80181 76766 80196
rect 77788 80760 77854 80775
rect 77788 80746 77795 80760
rect 77847 80746 77854 80760
rect 77788 80690 77793 80746
rect 77849 80690 77854 80746
rect 77788 80666 77795 80690
rect 77847 80666 77854 80690
rect 77788 80610 77793 80666
rect 77849 80610 77854 80666
rect 77788 80586 77795 80610
rect 77847 80586 77854 80610
rect 77788 80530 77793 80586
rect 77849 80530 77854 80586
rect 77788 80516 77795 80530
rect 77847 80516 77854 80530
rect 77788 80506 77854 80516
rect 77788 80450 77793 80506
rect 77849 80450 77854 80506
rect 77788 80440 77854 80450
rect 77788 80426 77795 80440
rect 77847 80426 77854 80440
rect 77788 80370 77793 80426
rect 77849 80370 77854 80426
rect 77788 80346 77795 80370
rect 77847 80346 77854 80370
rect 77788 80290 77793 80346
rect 77849 80290 77854 80346
rect 77788 80266 77795 80290
rect 77847 80266 77854 80290
rect 77788 80210 77793 80266
rect 77849 80210 77854 80266
rect 77788 80196 77795 80210
rect 77847 80196 77854 80210
rect 77788 80181 77854 80196
rect 78876 80760 78942 80775
rect 78876 80746 78883 80760
rect 78935 80746 78942 80760
rect 78876 80690 78881 80746
rect 78937 80690 78942 80746
rect 78876 80666 78883 80690
rect 78935 80666 78942 80690
rect 78876 80610 78881 80666
rect 78937 80610 78942 80666
rect 78876 80586 78883 80610
rect 78935 80586 78942 80610
rect 78876 80530 78881 80586
rect 78937 80530 78942 80586
rect 78876 80516 78883 80530
rect 78935 80516 78942 80530
rect 78876 80506 78942 80516
rect 78876 80450 78881 80506
rect 78937 80450 78942 80506
rect 78876 80440 78942 80450
rect 78876 80426 78883 80440
rect 78935 80426 78942 80440
rect 78876 80370 78881 80426
rect 78937 80370 78942 80426
rect 78876 80346 78883 80370
rect 78935 80346 78942 80370
rect 78876 80290 78881 80346
rect 78937 80290 78942 80346
rect 78876 80266 78883 80290
rect 78935 80266 78942 80290
rect 78876 80210 78881 80266
rect 78937 80210 78942 80266
rect 78876 80196 78883 80210
rect 78935 80196 78942 80210
rect 78876 80181 78942 80196
rect 79964 80760 80030 80775
rect 79964 80746 79971 80760
rect 80023 80746 80030 80760
rect 79964 80690 79969 80746
rect 80025 80690 80030 80746
rect 79964 80666 79971 80690
rect 80023 80666 80030 80690
rect 79964 80610 79969 80666
rect 80025 80610 80030 80666
rect 79964 80586 79971 80610
rect 80023 80586 80030 80610
rect 79964 80530 79969 80586
rect 80025 80530 80030 80586
rect 79964 80516 79971 80530
rect 80023 80516 80030 80530
rect 79964 80506 80030 80516
rect 79964 80450 79969 80506
rect 80025 80450 80030 80506
rect 79964 80440 80030 80450
rect 79964 80426 79971 80440
rect 80023 80426 80030 80440
rect 79964 80370 79969 80426
rect 80025 80370 80030 80426
rect 79964 80346 79971 80370
rect 80023 80346 80030 80370
rect 79964 80290 79969 80346
rect 80025 80290 80030 80346
rect 79964 80266 79971 80290
rect 80023 80266 80030 80290
rect 79964 80210 79969 80266
rect 80025 80210 80030 80266
rect 79964 80196 79971 80210
rect 80023 80196 80030 80210
rect 79964 80181 80030 80196
rect 81052 80760 81118 80775
rect 81052 80746 81059 80760
rect 81111 80746 81118 80760
rect 81052 80690 81057 80746
rect 81113 80690 81118 80746
rect 81052 80666 81059 80690
rect 81111 80666 81118 80690
rect 81052 80610 81057 80666
rect 81113 80610 81118 80666
rect 81052 80586 81059 80610
rect 81111 80586 81118 80610
rect 81052 80530 81057 80586
rect 81113 80530 81118 80586
rect 81052 80516 81059 80530
rect 81111 80516 81118 80530
rect 81052 80506 81118 80516
rect 81052 80450 81057 80506
rect 81113 80450 81118 80506
rect 81052 80440 81118 80450
rect 81052 80426 81059 80440
rect 81111 80426 81118 80440
rect 81052 80370 81057 80426
rect 81113 80370 81118 80426
rect 81052 80346 81059 80370
rect 81111 80346 81118 80370
rect 81052 80290 81057 80346
rect 81113 80290 81118 80346
rect 81052 80266 81059 80290
rect 81111 80266 81118 80290
rect 81052 80210 81057 80266
rect 81113 80210 81118 80266
rect 81052 80196 81059 80210
rect 81111 80196 81118 80210
rect 81052 80181 81118 80196
rect 82140 80760 82206 80775
rect 82140 80746 82147 80760
rect 82199 80746 82206 80760
rect 82140 80690 82145 80746
rect 82201 80690 82206 80746
rect 82140 80666 82147 80690
rect 82199 80666 82206 80690
rect 82140 80610 82145 80666
rect 82201 80610 82206 80666
rect 82140 80586 82147 80610
rect 82199 80586 82206 80610
rect 82140 80530 82145 80586
rect 82201 80530 82206 80586
rect 82140 80516 82147 80530
rect 82199 80516 82206 80530
rect 82140 80506 82206 80516
rect 82140 80450 82145 80506
rect 82201 80450 82206 80506
rect 82140 80440 82206 80450
rect 82140 80426 82147 80440
rect 82199 80426 82206 80440
rect 82140 80370 82145 80426
rect 82201 80370 82206 80426
rect 82140 80346 82147 80370
rect 82199 80346 82206 80370
rect 82140 80290 82145 80346
rect 82201 80290 82206 80346
rect 82140 80266 82147 80290
rect 82199 80266 82206 80290
rect 82140 80210 82145 80266
rect 82201 80210 82206 80266
rect 82140 80196 82147 80210
rect 82199 80196 82206 80210
rect 82140 80181 82206 80196
rect 83228 80760 83294 80775
rect 83228 80746 83235 80760
rect 83287 80746 83294 80760
rect 83228 80690 83233 80746
rect 83289 80690 83294 80746
rect 83228 80666 83235 80690
rect 83287 80666 83294 80690
rect 83228 80610 83233 80666
rect 83289 80610 83294 80666
rect 83228 80586 83235 80610
rect 83287 80586 83294 80610
rect 83228 80530 83233 80586
rect 83289 80530 83294 80586
rect 83228 80516 83235 80530
rect 83287 80516 83294 80530
rect 83228 80506 83294 80516
rect 83228 80450 83233 80506
rect 83289 80450 83294 80506
rect 83228 80440 83294 80450
rect 83228 80426 83235 80440
rect 83287 80426 83294 80440
rect 83228 80370 83233 80426
rect 83289 80370 83294 80426
rect 83228 80346 83235 80370
rect 83287 80346 83294 80370
rect 83228 80290 83233 80346
rect 83289 80290 83294 80346
rect 83228 80266 83235 80290
rect 83287 80266 83294 80290
rect 83228 80210 83233 80266
rect 83289 80210 83294 80266
rect 83228 80196 83235 80210
rect 83287 80196 83294 80210
rect 83228 80181 83294 80196
rect 84316 80760 84382 80775
rect 84316 80746 84323 80760
rect 84375 80746 84382 80760
rect 84316 80690 84321 80746
rect 84377 80690 84382 80746
rect 84316 80666 84323 80690
rect 84375 80666 84382 80690
rect 84316 80610 84321 80666
rect 84377 80610 84382 80666
rect 84316 80586 84323 80610
rect 84375 80586 84382 80610
rect 84316 80530 84321 80586
rect 84377 80530 84382 80586
rect 84316 80516 84323 80530
rect 84375 80516 84382 80530
rect 84316 80506 84382 80516
rect 84316 80450 84321 80506
rect 84377 80450 84382 80506
rect 84316 80440 84382 80450
rect 84316 80426 84323 80440
rect 84375 80426 84382 80440
rect 84316 80370 84321 80426
rect 84377 80370 84382 80426
rect 84316 80346 84323 80370
rect 84375 80346 84382 80370
rect 84316 80290 84321 80346
rect 84377 80290 84382 80346
rect 84316 80266 84323 80290
rect 84375 80266 84382 80290
rect 84316 80210 84321 80266
rect 84377 80210 84382 80266
rect 84316 80196 84323 80210
rect 84375 80196 84382 80210
rect 84316 80181 84382 80196
rect 85404 80760 85470 80775
rect 85404 80746 85411 80760
rect 85463 80746 85470 80760
rect 85404 80690 85409 80746
rect 85465 80690 85470 80746
rect 85404 80666 85411 80690
rect 85463 80666 85470 80690
rect 85404 80610 85409 80666
rect 85465 80610 85470 80666
rect 85404 80586 85411 80610
rect 85463 80586 85470 80610
rect 85404 80530 85409 80586
rect 85465 80530 85470 80586
rect 85404 80516 85411 80530
rect 85463 80516 85470 80530
rect 85404 80506 85470 80516
rect 85404 80450 85409 80506
rect 85465 80450 85470 80506
rect 85404 80440 85470 80450
rect 85404 80426 85411 80440
rect 85463 80426 85470 80440
rect 85404 80370 85409 80426
rect 85465 80370 85470 80426
rect 85404 80346 85411 80370
rect 85463 80346 85470 80370
rect 85404 80290 85409 80346
rect 85465 80290 85470 80346
rect 85404 80266 85411 80290
rect 85463 80266 85470 80290
rect 85404 80210 85409 80266
rect 85465 80210 85470 80266
rect 85404 80196 85411 80210
rect 85463 80196 85470 80210
rect 85404 80181 85470 80196
rect 86492 80760 86558 80775
rect 86492 80746 86499 80760
rect 86551 80746 86558 80760
rect 86492 80690 86497 80746
rect 86553 80690 86558 80746
rect 86492 80666 86499 80690
rect 86551 80666 86558 80690
rect 86492 80610 86497 80666
rect 86553 80610 86558 80666
rect 86492 80586 86499 80610
rect 86551 80586 86558 80610
rect 86492 80530 86497 80586
rect 86553 80530 86558 80586
rect 86492 80516 86499 80530
rect 86551 80516 86558 80530
rect 86492 80506 86558 80516
rect 86492 80450 86497 80506
rect 86553 80450 86558 80506
rect 86492 80440 86558 80450
rect 86492 80426 86499 80440
rect 86551 80426 86558 80440
rect 86492 80370 86497 80426
rect 86553 80370 86558 80426
rect 86492 80346 86499 80370
rect 86551 80346 86558 80370
rect 86492 80290 86497 80346
rect 86553 80290 86558 80346
rect 86492 80266 86499 80290
rect 86551 80266 86558 80290
rect 86492 80210 86497 80266
rect 86553 80210 86558 80266
rect 86492 80196 86499 80210
rect 86551 80196 86558 80210
rect 86492 80181 86558 80196
rect 87580 80760 87646 80775
rect 87580 80746 87587 80760
rect 87639 80746 87646 80760
rect 87580 80690 87585 80746
rect 87641 80690 87646 80746
rect 87580 80666 87587 80690
rect 87639 80666 87646 80690
rect 87580 80610 87585 80666
rect 87641 80610 87646 80666
rect 87580 80586 87587 80610
rect 87639 80586 87646 80610
rect 87580 80530 87585 80586
rect 87641 80530 87646 80586
rect 87580 80516 87587 80530
rect 87639 80516 87646 80530
rect 87580 80506 87646 80516
rect 87580 80450 87585 80506
rect 87641 80450 87646 80506
rect 87580 80440 87646 80450
rect 87580 80426 87587 80440
rect 87639 80426 87646 80440
rect 87580 80370 87585 80426
rect 87641 80370 87646 80426
rect 87580 80346 87587 80370
rect 87639 80346 87646 80370
rect 87580 80290 87585 80346
rect 87641 80290 87646 80346
rect 87580 80266 87587 80290
rect 87639 80266 87646 80290
rect 87580 80210 87585 80266
rect 87641 80210 87646 80266
rect 87580 80196 87587 80210
rect 87639 80196 87646 80210
rect 87580 80181 87646 80196
rect 88668 80760 88734 80775
rect 88668 80746 88675 80760
rect 88727 80746 88734 80760
rect 88668 80690 88673 80746
rect 88729 80690 88734 80746
rect 88668 80666 88675 80690
rect 88727 80666 88734 80690
rect 88668 80610 88673 80666
rect 88729 80610 88734 80666
rect 88668 80586 88675 80610
rect 88727 80586 88734 80610
rect 88668 80530 88673 80586
rect 88729 80530 88734 80586
rect 88668 80516 88675 80530
rect 88727 80516 88734 80530
rect 88668 80506 88734 80516
rect 88668 80450 88673 80506
rect 88729 80450 88734 80506
rect 88668 80440 88734 80450
rect 88668 80426 88675 80440
rect 88727 80426 88734 80440
rect 88668 80370 88673 80426
rect 88729 80370 88734 80426
rect 88668 80346 88675 80370
rect 88727 80346 88734 80370
rect 88668 80290 88673 80346
rect 88729 80290 88734 80346
rect 88668 80266 88675 80290
rect 88727 80266 88734 80290
rect 88668 80210 88673 80266
rect 88729 80210 88734 80266
rect 88668 80196 88675 80210
rect 88727 80196 88734 80210
rect 88668 80181 88734 80196
rect 75069 78757 75135 78772
rect 75069 78743 75076 78757
rect 75128 78743 75135 78757
rect 75069 78687 75074 78743
rect 75130 78687 75135 78743
rect 75069 78663 75076 78687
rect 75128 78663 75135 78687
rect 75069 78607 75074 78663
rect 75130 78607 75135 78663
rect 75069 78583 75076 78607
rect 75128 78583 75135 78607
rect 75069 78527 75074 78583
rect 75130 78527 75135 78583
rect 75069 78513 75076 78527
rect 75128 78513 75135 78527
rect 75069 78503 75135 78513
rect 75069 78447 75074 78503
rect 75130 78447 75135 78503
rect 75069 78437 75135 78447
rect 75069 78423 75076 78437
rect 75128 78423 75135 78437
rect 75069 78367 75074 78423
rect 75130 78367 75135 78423
rect 75069 78343 75076 78367
rect 75128 78343 75135 78367
rect 75069 78287 75074 78343
rect 75130 78287 75135 78343
rect 75069 78263 75076 78287
rect 75128 78263 75135 78287
rect 75069 78207 75074 78263
rect 75130 78207 75135 78263
rect 75069 78193 75076 78207
rect 75128 78193 75135 78207
rect 75069 78178 75135 78193
rect 76157 78757 76223 78772
rect 76157 78743 76164 78757
rect 76216 78743 76223 78757
rect 76157 78687 76162 78743
rect 76218 78687 76223 78743
rect 76157 78663 76164 78687
rect 76216 78663 76223 78687
rect 76157 78607 76162 78663
rect 76218 78607 76223 78663
rect 76157 78583 76164 78607
rect 76216 78583 76223 78607
rect 76157 78527 76162 78583
rect 76218 78527 76223 78583
rect 76157 78513 76164 78527
rect 76216 78513 76223 78527
rect 76157 78503 76223 78513
rect 76157 78447 76162 78503
rect 76218 78447 76223 78503
rect 76157 78437 76223 78447
rect 76157 78423 76164 78437
rect 76216 78423 76223 78437
rect 76157 78367 76162 78423
rect 76218 78367 76223 78423
rect 76157 78343 76164 78367
rect 76216 78343 76223 78367
rect 76157 78287 76162 78343
rect 76218 78287 76223 78343
rect 76157 78263 76164 78287
rect 76216 78263 76223 78287
rect 76157 78207 76162 78263
rect 76218 78207 76223 78263
rect 76157 78193 76164 78207
rect 76216 78193 76223 78207
rect 76157 78178 76223 78193
rect 77245 78757 77311 78772
rect 77245 78743 77252 78757
rect 77304 78743 77311 78757
rect 77245 78687 77250 78743
rect 77306 78687 77311 78743
rect 77245 78663 77252 78687
rect 77304 78663 77311 78687
rect 77245 78607 77250 78663
rect 77306 78607 77311 78663
rect 77245 78583 77252 78607
rect 77304 78583 77311 78607
rect 77245 78527 77250 78583
rect 77306 78527 77311 78583
rect 77245 78513 77252 78527
rect 77304 78513 77311 78527
rect 77245 78503 77311 78513
rect 77245 78447 77250 78503
rect 77306 78447 77311 78503
rect 77245 78437 77311 78447
rect 77245 78423 77252 78437
rect 77304 78423 77311 78437
rect 77245 78367 77250 78423
rect 77306 78367 77311 78423
rect 77245 78343 77252 78367
rect 77304 78343 77311 78367
rect 77245 78287 77250 78343
rect 77306 78287 77311 78343
rect 77245 78263 77252 78287
rect 77304 78263 77311 78287
rect 77245 78207 77250 78263
rect 77306 78207 77311 78263
rect 77245 78193 77252 78207
rect 77304 78193 77311 78207
rect 77245 78178 77311 78193
rect 78333 78757 78399 78772
rect 78333 78743 78340 78757
rect 78392 78743 78399 78757
rect 78333 78687 78338 78743
rect 78394 78687 78399 78743
rect 78333 78663 78340 78687
rect 78392 78663 78399 78687
rect 78333 78607 78338 78663
rect 78394 78607 78399 78663
rect 78333 78583 78340 78607
rect 78392 78583 78399 78607
rect 78333 78527 78338 78583
rect 78394 78527 78399 78583
rect 78333 78513 78340 78527
rect 78392 78513 78399 78527
rect 78333 78503 78399 78513
rect 78333 78447 78338 78503
rect 78394 78447 78399 78503
rect 78333 78437 78399 78447
rect 78333 78423 78340 78437
rect 78392 78423 78399 78437
rect 78333 78367 78338 78423
rect 78394 78367 78399 78423
rect 78333 78343 78340 78367
rect 78392 78343 78399 78367
rect 78333 78287 78338 78343
rect 78394 78287 78399 78343
rect 78333 78263 78340 78287
rect 78392 78263 78399 78287
rect 78333 78207 78338 78263
rect 78394 78207 78399 78263
rect 78333 78193 78340 78207
rect 78392 78193 78399 78207
rect 78333 78178 78399 78193
rect 79421 78757 79487 78772
rect 79421 78743 79428 78757
rect 79480 78743 79487 78757
rect 79421 78687 79426 78743
rect 79482 78687 79487 78743
rect 79421 78663 79428 78687
rect 79480 78663 79487 78687
rect 79421 78607 79426 78663
rect 79482 78607 79487 78663
rect 79421 78583 79428 78607
rect 79480 78583 79487 78607
rect 79421 78527 79426 78583
rect 79482 78527 79487 78583
rect 79421 78513 79428 78527
rect 79480 78513 79487 78527
rect 79421 78503 79487 78513
rect 79421 78447 79426 78503
rect 79482 78447 79487 78503
rect 79421 78437 79487 78447
rect 79421 78423 79428 78437
rect 79480 78423 79487 78437
rect 79421 78367 79426 78423
rect 79482 78367 79487 78423
rect 79421 78343 79428 78367
rect 79480 78343 79487 78367
rect 79421 78287 79426 78343
rect 79482 78287 79487 78343
rect 79421 78263 79428 78287
rect 79480 78263 79487 78287
rect 79421 78207 79426 78263
rect 79482 78207 79487 78263
rect 79421 78193 79428 78207
rect 79480 78193 79487 78207
rect 79421 78178 79487 78193
rect 80509 78757 80575 78772
rect 80509 78743 80516 78757
rect 80568 78743 80575 78757
rect 80509 78687 80514 78743
rect 80570 78687 80575 78743
rect 80509 78663 80516 78687
rect 80568 78663 80575 78687
rect 80509 78607 80514 78663
rect 80570 78607 80575 78663
rect 80509 78583 80516 78607
rect 80568 78583 80575 78607
rect 80509 78527 80514 78583
rect 80570 78527 80575 78583
rect 80509 78513 80516 78527
rect 80568 78513 80575 78527
rect 80509 78503 80575 78513
rect 80509 78447 80514 78503
rect 80570 78447 80575 78503
rect 80509 78437 80575 78447
rect 80509 78423 80516 78437
rect 80568 78423 80575 78437
rect 80509 78367 80514 78423
rect 80570 78367 80575 78423
rect 80509 78343 80516 78367
rect 80568 78343 80575 78367
rect 80509 78287 80514 78343
rect 80570 78287 80575 78343
rect 80509 78263 80516 78287
rect 80568 78263 80575 78287
rect 80509 78207 80514 78263
rect 80570 78207 80575 78263
rect 80509 78193 80516 78207
rect 80568 78193 80575 78207
rect 80509 78178 80575 78193
rect 81597 78757 81663 78772
rect 81597 78743 81604 78757
rect 81656 78743 81663 78757
rect 81597 78687 81602 78743
rect 81658 78687 81663 78743
rect 81597 78663 81604 78687
rect 81656 78663 81663 78687
rect 81597 78607 81602 78663
rect 81658 78607 81663 78663
rect 81597 78583 81604 78607
rect 81656 78583 81663 78607
rect 81597 78527 81602 78583
rect 81658 78527 81663 78583
rect 81597 78513 81604 78527
rect 81656 78513 81663 78527
rect 81597 78503 81663 78513
rect 81597 78447 81602 78503
rect 81658 78447 81663 78503
rect 81597 78437 81663 78447
rect 81597 78423 81604 78437
rect 81656 78423 81663 78437
rect 81597 78367 81602 78423
rect 81658 78367 81663 78423
rect 81597 78343 81604 78367
rect 81656 78343 81663 78367
rect 81597 78287 81602 78343
rect 81658 78287 81663 78343
rect 81597 78263 81604 78287
rect 81656 78263 81663 78287
rect 81597 78207 81602 78263
rect 81658 78207 81663 78263
rect 81597 78193 81604 78207
rect 81656 78193 81663 78207
rect 81597 78178 81663 78193
rect 82685 78757 82751 78772
rect 82685 78743 82692 78757
rect 82744 78743 82751 78757
rect 82685 78687 82690 78743
rect 82746 78687 82751 78743
rect 82685 78663 82692 78687
rect 82744 78663 82751 78687
rect 82685 78607 82690 78663
rect 82746 78607 82751 78663
rect 82685 78583 82692 78607
rect 82744 78583 82751 78607
rect 82685 78527 82690 78583
rect 82746 78527 82751 78583
rect 82685 78513 82692 78527
rect 82744 78513 82751 78527
rect 82685 78503 82751 78513
rect 82685 78447 82690 78503
rect 82746 78447 82751 78503
rect 82685 78437 82751 78447
rect 82685 78423 82692 78437
rect 82744 78423 82751 78437
rect 82685 78367 82690 78423
rect 82746 78367 82751 78423
rect 82685 78343 82692 78367
rect 82744 78343 82751 78367
rect 82685 78287 82690 78343
rect 82746 78287 82751 78343
rect 82685 78263 82692 78287
rect 82744 78263 82751 78287
rect 82685 78207 82690 78263
rect 82746 78207 82751 78263
rect 82685 78193 82692 78207
rect 82744 78193 82751 78207
rect 82685 78178 82751 78193
rect 83773 78757 83839 78772
rect 83773 78743 83780 78757
rect 83832 78743 83839 78757
rect 83773 78687 83778 78743
rect 83834 78687 83839 78743
rect 83773 78663 83780 78687
rect 83832 78663 83839 78687
rect 83773 78607 83778 78663
rect 83834 78607 83839 78663
rect 83773 78583 83780 78607
rect 83832 78583 83839 78607
rect 83773 78527 83778 78583
rect 83834 78527 83839 78583
rect 83773 78513 83780 78527
rect 83832 78513 83839 78527
rect 83773 78503 83839 78513
rect 83773 78447 83778 78503
rect 83834 78447 83839 78503
rect 83773 78437 83839 78447
rect 83773 78423 83780 78437
rect 83832 78423 83839 78437
rect 83773 78367 83778 78423
rect 83834 78367 83839 78423
rect 83773 78343 83780 78367
rect 83832 78343 83839 78367
rect 83773 78287 83778 78343
rect 83834 78287 83839 78343
rect 83773 78263 83780 78287
rect 83832 78263 83839 78287
rect 83773 78207 83778 78263
rect 83834 78207 83839 78263
rect 83773 78193 83780 78207
rect 83832 78193 83839 78207
rect 83773 78178 83839 78193
rect 84861 78757 84927 78772
rect 84861 78743 84868 78757
rect 84920 78743 84927 78757
rect 84861 78687 84866 78743
rect 84922 78687 84927 78743
rect 84861 78663 84868 78687
rect 84920 78663 84927 78687
rect 84861 78607 84866 78663
rect 84922 78607 84927 78663
rect 84861 78583 84868 78607
rect 84920 78583 84927 78607
rect 84861 78527 84866 78583
rect 84922 78527 84927 78583
rect 84861 78513 84868 78527
rect 84920 78513 84927 78527
rect 84861 78503 84927 78513
rect 84861 78447 84866 78503
rect 84922 78447 84927 78503
rect 84861 78437 84927 78447
rect 84861 78423 84868 78437
rect 84920 78423 84927 78437
rect 84861 78367 84866 78423
rect 84922 78367 84927 78423
rect 84861 78343 84868 78367
rect 84920 78343 84927 78367
rect 84861 78287 84866 78343
rect 84922 78287 84927 78343
rect 84861 78263 84868 78287
rect 84920 78263 84927 78287
rect 84861 78207 84866 78263
rect 84922 78207 84927 78263
rect 84861 78193 84868 78207
rect 84920 78193 84927 78207
rect 84861 78178 84927 78193
rect 85949 78757 86015 78772
rect 85949 78743 85956 78757
rect 86008 78743 86015 78757
rect 85949 78687 85954 78743
rect 86010 78687 86015 78743
rect 85949 78663 85956 78687
rect 86008 78663 86015 78687
rect 85949 78607 85954 78663
rect 86010 78607 86015 78663
rect 85949 78583 85956 78607
rect 86008 78583 86015 78607
rect 85949 78527 85954 78583
rect 86010 78527 86015 78583
rect 85949 78513 85956 78527
rect 86008 78513 86015 78527
rect 85949 78503 86015 78513
rect 85949 78447 85954 78503
rect 86010 78447 86015 78503
rect 85949 78437 86015 78447
rect 85949 78423 85956 78437
rect 86008 78423 86015 78437
rect 85949 78367 85954 78423
rect 86010 78367 86015 78423
rect 85949 78343 85956 78367
rect 86008 78343 86015 78367
rect 85949 78287 85954 78343
rect 86010 78287 86015 78343
rect 85949 78263 85956 78287
rect 86008 78263 86015 78287
rect 85949 78207 85954 78263
rect 86010 78207 86015 78263
rect 85949 78193 85956 78207
rect 86008 78193 86015 78207
rect 85949 78178 86015 78193
rect 87037 78757 87103 78772
rect 87037 78743 87044 78757
rect 87096 78743 87103 78757
rect 87037 78687 87042 78743
rect 87098 78687 87103 78743
rect 87037 78663 87044 78687
rect 87096 78663 87103 78687
rect 87037 78607 87042 78663
rect 87098 78607 87103 78663
rect 87037 78583 87044 78607
rect 87096 78583 87103 78607
rect 87037 78527 87042 78583
rect 87098 78527 87103 78583
rect 87037 78513 87044 78527
rect 87096 78513 87103 78527
rect 87037 78503 87103 78513
rect 87037 78447 87042 78503
rect 87098 78447 87103 78503
rect 87037 78437 87103 78447
rect 87037 78423 87044 78437
rect 87096 78423 87103 78437
rect 87037 78367 87042 78423
rect 87098 78367 87103 78423
rect 87037 78343 87044 78367
rect 87096 78343 87103 78367
rect 87037 78287 87042 78343
rect 87098 78287 87103 78343
rect 87037 78263 87044 78287
rect 87096 78263 87103 78287
rect 87037 78207 87042 78263
rect 87098 78207 87103 78263
rect 87037 78193 87044 78207
rect 87096 78193 87103 78207
rect 87037 78178 87103 78193
rect 88125 78757 88191 78772
rect 88125 78743 88132 78757
rect 88184 78743 88191 78757
rect 88125 78687 88130 78743
rect 88186 78687 88191 78743
rect 88125 78663 88132 78687
rect 88184 78663 88191 78687
rect 88125 78607 88130 78663
rect 88186 78607 88191 78663
rect 88125 78583 88132 78607
rect 88184 78583 88191 78607
rect 88125 78527 88130 78583
rect 88186 78527 88191 78583
rect 88125 78513 88132 78527
rect 88184 78513 88191 78527
rect 88125 78503 88191 78513
rect 88125 78447 88130 78503
rect 88186 78447 88191 78503
rect 88125 78437 88191 78447
rect 88125 78423 88132 78437
rect 88184 78423 88191 78437
rect 88125 78367 88130 78423
rect 88186 78367 88191 78423
rect 88125 78343 88132 78367
rect 88184 78343 88191 78367
rect 88125 78287 88130 78343
rect 88186 78287 88191 78343
rect 88125 78263 88132 78287
rect 88184 78263 88191 78287
rect 88125 78207 88130 78263
rect 88186 78207 88191 78263
rect 88125 78193 88132 78207
rect 88184 78193 88191 78207
rect 88125 78178 88191 78193
rect 74524 76760 74590 76775
rect 74524 76746 74531 76760
rect 74583 76746 74590 76760
rect 74524 76690 74529 76746
rect 74585 76690 74590 76746
rect 74524 76666 74531 76690
rect 74583 76666 74590 76690
rect 74524 76610 74529 76666
rect 74585 76610 74590 76666
rect 74524 76586 74531 76610
rect 74583 76586 74590 76610
rect 74524 76530 74529 76586
rect 74585 76530 74590 76586
rect 74524 76516 74531 76530
rect 74583 76516 74590 76530
rect 74524 76506 74590 76516
rect 74524 76450 74529 76506
rect 74585 76450 74590 76506
rect 74524 76440 74590 76450
rect 74524 76426 74531 76440
rect 74583 76426 74590 76440
rect 74524 76370 74529 76426
rect 74585 76370 74590 76426
rect 74524 76346 74531 76370
rect 74583 76346 74590 76370
rect 74524 76290 74529 76346
rect 74585 76290 74590 76346
rect 74524 76266 74531 76290
rect 74583 76266 74590 76290
rect 74524 76210 74529 76266
rect 74585 76210 74590 76266
rect 74524 76196 74531 76210
rect 74583 76196 74590 76210
rect 74524 76181 74590 76196
rect 75612 76760 75678 76775
rect 75612 76746 75619 76760
rect 75671 76746 75678 76760
rect 75612 76690 75617 76746
rect 75673 76690 75678 76746
rect 75612 76666 75619 76690
rect 75671 76666 75678 76690
rect 75612 76610 75617 76666
rect 75673 76610 75678 76666
rect 75612 76586 75619 76610
rect 75671 76586 75678 76610
rect 75612 76530 75617 76586
rect 75673 76530 75678 76586
rect 75612 76516 75619 76530
rect 75671 76516 75678 76530
rect 75612 76506 75678 76516
rect 75612 76450 75617 76506
rect 75673 76450 75678 76506
rect 75612 76440 75678 76450
rect 75612 76426 75619 76440
rect 75671 76426 75678 76440
rect 75612 76370 75617 76426
rect 75673 76370 75678 76426
rect 75612 76346 75619 76370
rect 75671 76346 75678 76370
rect 75612 76290 75617 76346
rect 75673 76290 75678 76346
rect 75612 76266 75619 76290
rect 75671 76266 75678 76290
rect 75612 76210 75617 76266
rect 75673 76210 75678 76266
rect 75612 76196 75619 76210
rect 75671 76196 75678 76210
rect 75612 76181 75678 76196
rect 76700 76760 76766 76775
rect 76700 76746 76707 76760
rect 76759 76746 76766 76760
rect 76700 76690 76705 76746
rect 76761 76690 76766 76746
rect 76700 76666 76707 76690
rect 76759 76666 76766 76690
rect 76700 76610 76705 76666
rect 76761 76610 76766 76666
rect 76700 76586 76707 76610
rect 76759 76586 76766 76610
rect 76700 76530 76705 76586
rect 76761 76530 76766 76586
rect 76700 76516 76707 76530
rect 76759 76516 76766 76530
rect 76700 76506 76766 76516
rect 76700 76450 76705 76506
rect 76761 76450 76766 76506
rect 76700 76440 76766 76450
rect 76700 76426 76707 76440
rect 76759 76426 76766 76440
rect 76700 76370 76705 76426
rect 76761 76370 76766 76426
rect 76700 76346 76707 76370
rect 76759 76346 76766 76370
rect 76700 76290 76705 76346
rect 76761 76290 76766 76346
rect 76700 76266 76707 76290
rect 76759 76266 76766 76290
rect 76700 76210 76705 76266
rect 76761 76210 76766 76266
rect 76700 76196 76707 76210
rect 76759 76196 76766 76210
rect 76700 76181 76766 76196
rect 77788 76760 77854 76775
rect 77788 76746 77795 76760
rect 77847 76746 77854 76760
rect 77788 76690 77793 76746
rect 77849 76690 77854 76746
rect 77788 76666 77795 76690
rect 77847 76666 77854 76690
rect 77788 76610 77793 76666
rect 77849 76610 77854 76666
rect 77788 76586 77795 76610
rect 77847 76586 77854 76610
rect 77788 76530 77793 76586
rect 77849 76530 77854 76586
rect 77788 76516 77795 76530
rect 77847 76516 77854 76530
rect 77788 76506 77854 76516
rect 77788 76450 77793 76506
rect 77849 76450 77854 76506
rect 77788 76440 77854 76450
rect 77788 76426 77795 76440
rect 77847 76426 77854 76440
rect 77788 76370 77793 76426
rect 77849 76370 77854 76426
rect 77788 76346 77795 76370
rect 77847 76346 77854 76370
rect 77788 76290 77793 76346
rect 77849 76290 77854 76346
rect 77788 76266 77795 76290
rect 77847 76266 77854 76290
rect 77788 76210 77793 76266
rect 77849 76210 77854 76266
rect 77788 76196 77795 76210
rect 77847 76196 77854 76210
rect 77788 76181 77854 76196
rect 78876 76760 78942 76775
rect 78876 76746 78883 76760
rect 78935 76746 78942 76760
rect 78876 76690 78881 76746
rect 78937 76690 78942 76746
rect 78876 76666 78883 76690
rect 78935 76666 78942 76690
rect 78876 76610 78881 76666
rect 78937 76610 78942 76666
rect 78876 76586 78883 76610
rect 78935 76586 78942 76610
rect 78876 76530 78881 76586
rect 78937 76530 78942 76586
rect 78876 76516 78883 76530
rect 78935 76516 78942 76530
rect 78876 76506 78942 76516
rect 78876 76450 78881 76506
rect 78937 76450 78942 76506
rect 78876 76440 78942 76450
rect 78876 76426 78883 76440
rect 78935 76426 78942 76440
rect 78876 76370 78881 76426
rect 78937 76370 78942 76426
rect 78876 76346 78883 76370
rect 78935 76346 78942 76370
rect 78876 76290 78881 76346
rect 78937 76290 78942 76346
rect 78876 76266 78883 76290
rect 78935 76266 78942 76290
rect 78876 76210 78881 76266
rect 78937 76210 78942 76266
rect 78876 76196 78883 76210
rect 78935 76196 78942 76210
rect 78876 76181 78942 76196
rect 79964 76760 80030 76775
rect 79964 76746 79971 76760
rect 80023 76746 80030 76760
rect 79964 76690 79969 76746
rect 80025 76690 80030 76746
rect 79964 76666 79971 76690
rect 80023 76666 80030 76690
rect 79964 76610 79969 76666
rect 80025 76610 80030 76666
rect 79964 76586 79971 76610
rect 80023 76586 80030 76610
rect 79964 76530 79969 76586
rect 80025 76530 80030 76586
rect 79964 76516 79971 76530
rect 80023 76516 80030 76530
rect 79964 76506 80030 76516
rect 79964 76450 79969 76506
rect 80025 76450 80030 76506
rect 79964 76440 80030 76450
rect 79964 76426 79971 76440
rect 80023 76426 80030 76440
rect 79964 76370 79969 76426
rect 80025 76370 80030 76426
rect 79964 76346 79971 76370
rect 80023 76346 80030 76370
rect 79964 76290 79969 76346
rect 80025 76290 80030 76346
rect 79964 76266 79971 76290
rect 80023 76266 80030 76290
rect 79964 76210 79969 76266
rect 80025 76210 80030 76266
rect 79964 76196 79971 76210
rect 80023 76196 80030 76210
rect 79964 76181 80030 76196
rect 81052 76760 81118 76775
rect 81052 76746 81059 76760
rect 81111 76746 81118 76760
rect 81052 76690 81057 76746
rect 81113 76690 81118 76746
rect 81052 76666 81059 76690
rect 81111 76666 81118 76690
rect 81052 76610 81057 76666
rect 81113 76610 81118 76666
rect 81052 76586 81059 76610
rect 81111 76586 81118 76610
rect 81052 76530 81057 76586
rect 81113 76530 81118 76586
rect 81052 76516 81059 76530
rect 81111 76516 81118 76530
rect 81052 76506 81118 76516
rect 81052 76450 81057 76506
rect 81113 76450 81118 76506
rect 81052 76440 81118 76450
rect 81052 76426 81059 76440
rect 81111 76426 81118 76440
rect 81052 76370 81057 76426
rect 81113 76370 81118 76426
rect 81052 76346 81059 76370
rect 81111 76346 81118 76370
rect 81052 76290 81057 76346
rect 81113 76290 81118 76346
rect 81052 76266 81059 76290
rect 81111 76266 81118 76290
rect 81052 76210 81057 76266
rect 81113 76210 81118 76266
rect 81052 76196 81059 76210
rect 81111 76196 81118 76210
rect 81052 76181 81118 76196
rect 82140 76760 82206 76775
rect 82140 76746 82147 76760
rect 82199 76746 82206 76760
rect 82140 76690 82145 76746
rect 82201 76690 82206 76746
rect 82140 76666 82147 76690
rect 82199 76666 82206 76690
rect 82140 76610 82145 76666
rect 82201 76610 82206 76666
rect 82140 76586 82147 76610
rect 82199 76586 82206 76610
rect 82140 76530 82145 76586
rect 82201 76530 82206 76586
rect 82140 76516 82147 76530
rect 82199 76516 82206 76530
rect 82140 76506 82206 76516
rect 82140 76450 82145 76506
rect 82201 76450 82206 76506
rect 82140 76440 82206 76450
rect 82140 76426 82147 76440
rect 82199 76426 82206 76440
rect 82140 76370 82145 76426
rect 82201 76370 82206 76426
rect 82140 76346 82147 76370
rect 82199 76346 82206 76370
rect 82140 76290 82145 76346
rect 82201 76290 82206 76346
rect 82140 76266 82147 76290
rect 82199 76266 82206 76290
rect 82140 76210 82145 76266
rect 82201 76210 82206 76266
rect 82140 76196 82147 76210
rect 82199 76196 82206 76210
rect 82140 76181 82206 76196
rect 83228 76760 83294 76775
rect 83228 76746 83235 76760
rect 83287 76746 83294 76760
rect 83228 76690 83233 76746
rect 83289 76690 83294 76746
rect 83228 76666 83235 76690
rect 83287 76666 83294 76690
rect 83228 76610 83233 76666
rect 83289 76610 83294 76666
rect 83228 76586 83235 76610
rect 83287 76586 83294 76610
rect 83228 76530 83233 76586
rect 83289 76530 83294 76586
rect 83228 76516 83235 76530
rect 83287 76516 83294 76530
rect 83228 76506 83294 76516
rect 83228 76450 83233 76506
rect 83289 76450 83294 76506
rect 83228 76440 83294 76450
rect 83228 76426 83235 76440
rect 83287 76426 83294 76440
rect 83228 76370 83233 76426
rect 83289 76370 83294 76426
rect 83228 76346 83235 76370
rect 83287 76346 83294 76370
rect 83228 76290 83233 76346
rect 83289 76290 83294 76346
rect 83228 76266 83235 76290
rect 83287 76266 83294 76290
rect 83228 76210 83233 76266
rect 83289 76210 83294 76266
rect 83228 76196 83235 76210
rect 83287 76196 83294 76210
rect 83228 76181 83294 76196
rect 84316 76760 84382 76775
rect 84316 76746 84323 76760
rect 84375 76746 84382 76760
rect 84316 76690 84321 76746
rect 84377 76690 84382 76746
rect 84316 76666 84323 76690
rect 84375 76666 84382 76690
rect 84316 76610 84321 76666
rect 84377 76610 84382 76666
rect 84316 76586 84323 76610
rect 84375 76586 84382 76610
rect 84316 76530 84321 76586
rect 84377 76530 84382 76586
rect 84316 76516 84323 76530
rect 84375 76516 84382 76530
rect 84316 76506 84382 76516
rect 84316 76450 84321 76506
rect 84377 76450 84382 76506
rect 84316 76440 84382 76450
rect 84316 76426 84323 76440
rect 84375 76426 84382 76440
rect 84316 76370 84321 76426
rect 84377 76370 84382 76426
rect 84316 76346 84323 76370
rect 84375 76346 84382 76370
rect 84316 76290 84321 76346
rect 84377 76290 84382 76346
rect 84316 76266 84323 76290
rect 84375 76266 84382 76290
rect 84316 76210 84321 76266
rect 84377 76210 84382 76266
rect 84316 76196 84323 76210
rect 84375 76196 84382 76210
rect 84316 76181 84382 76196
rect 85404 76760 85470 76775
rect 85404 76746 85411 76760
rect 85463 76746 85470 76760
rect 85404 76690 85409 76746
rect 85465 76690 85470 76746
rect 85404 76666 85411 76690
rect 85463 76666 85470 76690
rect 85404 76610 85409 76666
rect 85465 76610 85470 76666
rect 85404 76586 85411 76610
rect 85463 76586 85470 76610
rect 85404 76530 85409 76586
rect 85465 76530 85470 76586
rect 85404 76516 85411 76530
rect 85463 76516 85470 76530
rect 85404 76506 85470 76516
rect 85404 76450 85409 76506
rect 85465 76450 85470 76506
rect 85404 76440 85470 76450
rect 85404 76426 85411 76440
rect 85463 76426 85470 76440
rect 85404 76370 85409 76426
rect 85465 76370 85470 76426
rect 85404 76346 85411 76370
rect 85463 76346 85470 76370
rect 85404 76290 85409 76346
rect 85465 76290 85470 76346
rect 85404 76266 85411 76290
rect 85463 76266 85470 76290
rect 85404 76210 85409 76266
rect 85465 76210 85470 76266
rect 85404 76196 85411 76210
rect 85463 76196 85470 76210
rect 85404 76181 85470 76196
rect 86492 76760 86558 76775
rect 86492 76746 86499 76760
rect 86551 76746 86558 76760
rect 86492 76690 86497 76746
rect 86553 76690 86558 76746
rect 86492 76666 86499 76690
rect 86551 76666 86558 76690
rect 86492 76610 86497 76666
rect 86553 76610 86558 76666
rect 86492 76586 86499 76610
rect 86551 76586 86558 76610
rect 86492 76530 86497 76586
rect 86553 76530 86558 76586
rect 86492 76516 86499 76530
rect 86551 76516 86558 76530
rect 86492 76506 86558 76516
rect 86492 76450 86497 76506
rect 86553 76450 86558 76506
rect 86492 76440 86558 76450
rect 86492 76426 86499 76440
rect 86551 76426 86558 76440
rect 86492 76370 86497 76426
rect 86553 76370 86558 76426
rect 86492 76346 86499 76370
rect 86551 76346 86558 76370
rect 86492 76290 86497 76346
rect 86553 76290 86558 76346
rect 86492 76266 86499 76290
rect 86551 76266 86558 76290
rect 86492 76210 86497 76266
rect 86553 76210 86558 76266
rect 86492 76196 86499 76210
rect 86551 76196 86558 76210
rect 86492 76181 86558 76196
rect 87580 76760 87646 76775
rect 87580 76746 87587 76760
rect 87639 76746 87646 76760
rect 87580 76690 87585 76746
rect 87641 76690 87646 76746
rect 87580 76666 87587 76690
rect 87639 76666 87646 76690
rect 87580 76610 87585 76666
rect 87641 76610 87646 76666
rect 87580 76586 87587 76610
rect 87639 76586 87646 76610
rect 87580 76530 87585 76586
rect 87641 76530 87646 76586
rect 87580 76516 87587 76530
rect 87639 76516 87646 76530
rect 87580 76506 87646 76516
rect 87580 76450 87585 76506
rect 87641 76450 87646 76506
rect 87580 76440 87646 76450
rect 87580 76426 87587 76440
rect 87639 76426 87646 76440
rect 87580 76370 87585 76426
rect 87641 76370 87646 76426
rect 87580 76346 87587 76370
rect 87639 76346 87646 76370
rect 87580 76290 87585 76346
rect 87641 76290 87646 76346
rect 87580 76266 87587 76290
rect 87639 76266 87646 76290
rect 87580 76210 87585 76266
rect 87641 76210 87646 76266
rect 87580 76196 87587 76210
rect 87639 76196 87646 76210
rect 87580 76181 87646 76196
rect 88668 76760 88734 76775
rect 88668 76746 88675 76760
rect 88727 76746 88734 76760
rect 88668 76690 88673 76746
rect 88729 76690 88734 76746
rect 88668 76666 88675 76690
rect 88727 76666 88734 76690
rect 88668 76610 88673 76666
rect 88729 76610 88734 76666
rect 88668 76586 88675 76610
rect 88727 76586 88734 76610
rect 88668 76530 88673 76586
rect 88729 76530 88734 76586
rect 88668 76516 88675 76530
rect 88727 76516 88734 76530
rect 88668 76506 88734 76516
rect 88668 76450 88673 76506
rect 88729 76450 88734 76506
rect 88668 76440 88734 76450
rect 88668 76426 88675 76440
rect 88727 76426 88734 76440
rect 88668 76370 88673 76426
rect 88729 76370 88734 76426
rect 88668 76346 88675 76370
rect 88727 76346 88734 76370
rect 88668 76290 88673 76346
rect 88729 76290 88734 76346
rect 88668 76266 88675 76290
rect 88727 76266 88734 76290
rect 88668 76210 88673 76266
rect 88729 76210 88734 76266
rect 88668 76196 88675 76210
rect 88727 76196 88734 76210
rect 88668 76181 88734 76196
rect 75069 74757 75135 74772
rect 75069 74743 75076 74757
rect 75128 74743 75135 74757
rect 75069 74687 75074 74743
rect 75130 74687 75135 74743
rect 75069 74663 75076 74687
rect 75128 74663 75135 74687
rect 75069 74607 75074 74663
rect 75130 74607 75135 74663
rect 75069 74583 75076 74607
rect 75128 74583 75135 74607
rect 75069 74527 75074 74583
rect 75130 74527 75135 74583
rect 75069 74513 75076 74527
rect 75128 74513 75135 74527
rect 75069 74503 75135 74513
rect 75069 74447 75074 74503
rect 75130 74447 75135 74503
rect 75069 74437 75135 74447
rect 75069 74423 75076 74437
rect 75128 74423 75135 74437
rect 75069 74367 75074 74423
rect 75130 74367 75135 74423
rect 75069 74343 75076 74367
rect 75128 74343 75135 74367
rect 75069 74287 75074 74343
rect 75130 74287 75135 74343
rect 75069 74263 75076 74287
rect 75128 74263 75135 74287
rect 75069 74207 75074 74263
rect 75130 74207 75135 74263
rect 75069 74193 75076 74207
rect 75128 74193 75135 74207
rect 75069 74178 75135 74193
rect 77245 74757 77311 74772
rect 77245 74743 77252 74757
rect 77304 74743 77311 74757
rect 77245 74687 77250 74743
rect 77306 74687 77311 74743
rect 77245 74663 77252 74687
rect 77304 74663 77311 74687
rect 77245 74607 77250 74663
rect 77306 74607 77311 74663
rect 77245 74583 77252 74607
rect 77304 74583 77311 74607
rect 77245 74527 77250 74583
rect 77306 74527 77311 74583
rect 77245 74513 77252 74527
rect 77304 74513 77311 74527
rect 77245 74503 77311 74513
rect 77245 74447 77250 74503
rect 77306 74447 77311 74503
rect 77245 74437 77311 74447
rect 77245 74423 77252 74437
rect 77304 74423 77311 74437
rect 77245 74367 77250 74423
rect 77306 74367 77311 74423
rect 77245 74343 77252 74367
rect 77304 74343 77311 74367
rect 77245 74287 77250 74343
rect 77306 74287 77311 74343
rect 77245 74263 77252 74287
rect 77304 74263 77311 74287
rect 77245 74207 77250 74263
rect 77306 74207 77311 74263
rect 77245 74193 77252 74207
rect 77304 74193 77311 74207
rect 77245 74178 77311 74193
rect 78333 74757 78399 74772
rect 78333 74743 78340 74757
rect 78392 74743 78399 74757
rect 78333 74687 78338 74743
rect 78394 74687 78399 74743
rect 78333 74663 78340 74687
rect 78392 74663 78399 74687
rect 78333 74607 78338 74663
rect 78394 74607 78399 74663
rect 78333 74583 78340 74607
rect 78392 74583 78399 74607
rect 78333 74527 78338 74583
rect 78394 74527 78399 74583
rect 78333 74513 78340 74527
rect 78392 74513 78399 74527
rect 78333 74503 78399 74513
rect 78333 74447 78338 74503
rect 78394 74447 78399 74503
rect 78333 74437 78399 74447
rect 78333 74423 78340 74437
rect 78392 74423 78399 74437
rect 78333 74367 78338 74423
rect 78394 74367 78399 74423
rect 78333 74343 78340 74367
rect 78392 74343 78399 74367
rect 78333 74287 78338 74343
rect 78394 74287 78399 74343
rect 78333 74263 78340 74287
rect 78392 74263 78399 74287
rect 78333 74207 78338 74263
rect 78394 74207 78399 74263
rect 78333 74193 78340 74207
rect 78392 74193 78399 74207
rect 78333 74178 78399 74193
rect 80509 74757 80575 74772
rect 80509 74743 80516 74757
rect 80568 74743 80575 74757
rect 80509 74687 80514 74743
rect 80570 74687 80575 74743
rect 80509 74663 80516 74687
rect 80568 74663 80575 74687
rect 80509 74607 80514 74663
rect 80570 74607 80575 74663
rect 80509 74583 80516 74607
rect 80568 74583 80575 74607
rect 80509 74527 80514 74583
rect 80570 74527 80575 74583
rect 80509 74513 80516 74527
rect 80568 74513 80575 74527
rect 80509 74503 80575 74513
rect 80509 74447 80514 74503
rect 80570 74447 80575 74503
rect 80509 74437 80575 74447
rect 80509 74423 80516 74437
rect 80568 74423 80575 74437
rect 80509 74367 80514 74423
rect 80570 74367 80575 74423
rect 80509 74343 80516 74367
rect 80568 74343 80575 74367
rect 80509 74287 80514 74343
rect 80570 74287 80575 74343
rect 80509 74263 80516 74287
rect 80568 74263 80575 74287
rect 80509 74207 80514 74263
rect 80570 74207 80575 74263
rect 80509 74193 80516 74207
rect 80568 74193 80575 74207
rect 80509 74178 80575 74193
rect 81597 74757 81663 74772
rect 81597 74743 81604 74757
rect 81656 74743 81663 74757
rect 81597 74687 81602 74743
rect 81658 74687 81663 74743
rect 81597 74663 81604 74687
rect 81656 74663 81663 74687
rect 81597 74607 81602 74663
rect 81658 74607 81663 74663
rect 81597 74583 81604 74607
rect 81656 74583 81663 74607
rect 81597 74527 81602 74583
rect 81658 74527 81663 74583
rect 81597 74513 81604 74527
rect 81656 74513 81663 74527
rect 81597 74503 81663 74513
rect 81597 74447 81602 74503
rect 81658 74447 81663 74503
rect 81597 74437 81663 74447
rect 81597 74423 81604 74437
rect 81656 74423 81663 74437
rect 81597 74367 81602 74423
rect 81658 74367 81663 74423
rect 81597 74343 81604 74367
rect 81656 74343 81663 74367
rect 81597 74287 81602 74343
rect 81658 74287 81663 74343
rect 81597 74263 81604 74287
rect 81656 74263 81663 74287
rect 81597 74207 81602 74263
rect 81658 74207 81663 74263
rect 81597 74193 81604 74207
rect 81656 74193 81663 74207
rect 81597 74178 81663 74193
rect 82685 74757 82751 74772
rect 82685 74743 82692 74757
rect 82744 74743 82751 74757
rect 82685 74687 82690 74743
rect 82746 74687 82751 74743
rect 82685 74663 82692 74687
rect 82744 74663 82751 74687
rect 82685 74607 82690 74663
rect 82746 74607 82751 74663
rect 82685 74583 82692 74607
rect 82744 74583 82751 74607
rect 82685 74527 82690 74583
rect 82746 74527 82751 74583
rect 82685 74513 82692 74527
rect 82744 74513 82751 74527
rect 82685 74503 82751 74513
rect 82685 74447 82690 74503
rect 82746 74447 82751 74503
rect 82685 74437 82751 74447
rect 82685 74423 82692 74437
rect 82744 74423 82751 74437
rect 82685 74367 82690 74423
rect 82746 74367 82751 74423
rect 82685 74343 82692 74367
rect 82744 74343 82751 74367
rect 82685 74287 82690 74343
rect 82746 74287 82751 74343
rect 82685 74263 82692 74287
rect 82744 74263 82751 74287
rect 82685 74207 82690 74263
rect 82746 74207 82751 74263
rect 82685 74193 82692 74207
rect 82744 74193 82751 74207
rect 82685 74178 82751 74193
rect 84861 74757 84927 74772
rect 84861 74743 84868 74757
rect 84920 74743 84927 74757
rect 84861 74687 84866 74743
rect 84922 74687 84927 74743
rect 84861 74663 84868 74687
rect 84920 74663 84927 74687
rect 84861 74607 84866 74663
rect 84922 74607 84927 74663
rect 84861 74583 84868 74607
rect 84920 74583 84927 74607
rect 84861 74527 84866 74583
rect 84922 74527 84927 74583
rect 84861 74513 84868 74527
rect 84920 74513 84927 74527
rect 84861 74503 84927 74513
rect 84861 74447 84866 74503
rect 84922 74447 84927 74503
rect 84861 74437 84927 74447
rect 84861 74423 84868 74437
rect 84920 74423 84927 74437
rect 84861 74367 84866 74423
rect 84922 74367 84927 74423
rect 84861 74343 84868 74367
rect 84920 74343 84927 74367
rect 84861 74287 84866 74343
rect 84922 74287 84927 74343
rect 84861 74263 84868 74287
rect 84920 74263 84927 74287
rect 84861 74207 84866 74263
rect 84922 74207 84927 74263
rect 84861 74193 84868 74207
rect 84920 74193 84927 74207
rect 84861 74178 84927 74193
rect 85949 74757 86015 74772
rect 85949 74743 85956 74757
rect 86008 74743 86015 74757
rect 85949 74687 85954 74743
rect 86010 74687 86015 74743
rect 85949 74663 85956 74687
rect 86008 74663 86015 74687
rect 85949 74607 85954 74663
rect 86010 74607 86015 74663
rect 85949 74583 85956 74607
rect 86008 74583 86015 74607
rect 85949 74527 85954 74583
rect 86010 74527 86015 74583
rect 85949 74513 85956 74527
rect 86008 74513 86015 74527
rect 85949 74503 86015 74513
rect 85949 74447 85954 74503
rect 86010 74447 86015 74503
rect 85949 74437 86015 74447
rect 85949 74423 85956 74437
rect 86008 74423 86015 74437
rect 85949 74367 85954 74423
rect 86010 74367 86015 74423
rect 85949 74343 85956 74367
rect 86008 74343 86015 74367
rect 85949 74287 85954 74343
rect 86010 74287 86015 74343
rect 85949 74263 85956 74287
rect 86008 74263 86015 74287
rect 85949 74207 85954 74263
rect 86010 74207 86015 74263
rect 85949 74193 85956 74207
rect 86008 74193 86015 74207
rect 85949 74178 86015 74193
rect 88125 74757 88191 74772
rect 88125 74743 88132 74757
rect 88184 74743 88191 74757
rect 88125 74687 88130 74743
rect 88186 74687 88191 74743
rect 88125 74663 88132 74687
rect 88184 74663 88191 74687
rect 88125 74607 88130 74663
rect 88186 74607 88191 74663
rect 88125 74583 88132 74607
rect 88184 74583 88191 74607
rect 88125 74527 88130 74583
rect 88186 74527 88191 74583
rect 88125 74513 88132 74527
rect 88184 74513 88191 74527
rect 88125 74503 88191 74513
rect 88125 74447 88130 74503
rect 88186 74447 88191 74503
rect 88125 74437 88191 74447
rect 88125 74423 88132 74437
rect 88184 74423 88191 74437
rect 88125 74367 88130 74423
rect 88186 74367 88191 74423
rect 88125 74343 88132 74367
rect 88184 74343 88191 74367
rect 88125 74287 88130 74343
rect 88186 74287 88191 74343
rect 88125 74263 88132 74287
rect 88184 74263 88191 74287
rect 88125 74207 88130 74263
rect 88186 74207 88191 74263
rect 88125 74193 88132 74207
rect 88184 74193 88191 74207
rect 88125 74178 88191 74193
rect 74524 72760 74590 72775
rect 74524 72746 74531 72760
rect 74583 72746 74590 72760
rect 74524 72690 74529 72746
rect 74585 72690 74590 72746
rect 74524 72666 74531 72690
rect 74583 72666 74590 72690
rect 74524 72610 74529 72666
rect 74585 72610 74590 72666
rect 74524 72586 74531 72610
rect 74583 72586 74590 72610
rect 74524 72530 74529 72586
rect 74585 72530 74590 72586
rect 74524 72516 74531 72530
rect 74583 72516 74590 72530
rect 74524 72506 74590 72516
rect 74524 72450 74529 72506
rect 74585 72450 74590 72506
rect 74524 72440 74590 72450
rect 74524 72426 74531 72440
rect 74583 72426 74590 72440
rect 74524 72370 74529 72426
rect 74585 72370 74590 72426
rect 74524 72346 74531 72370
rect 74583 72346 74590 72370
rect 74524 72290 74529 72346
rect 74585 72290 74590 72346
rect 74524 72266 74531 72290
rect 74583 72266 74590 72290
rect 74524 72210 74529 72266
rect 74585 72210 74590 72266
rect 74524 72196 74531 72210
rect 74583 72196 74590 72210
rect 74524 72181 74590 72196
rect 75612 72760 75678 72775
rect 75612 72746 75619 72760
rect 75671 72746 75678 72760
rect 75612 72690 75617 72746
rect 75673 72690 75678 72746
rect 75612 72666 75619 72690
rect 75671 72666 75678 72690
rect 75612 72610 75617 72666
rect 75673 72610 75678 72666
rect 75612 72586 75619 72610
rect 75671 72586 75678 72610
rect 75612 72530 75617 72586
rect 75673 72530 75678 72586
rect 75612 72516 75619 72530
rect 75671 72516 75678 72530
rect 75612 72506 75678 72516
rect 75612 72450 75617 72506
rect 75673 72450 75678 72506
rect 75612 72440 75678 72450
rect 75612 72426 75619 72440
rect 75671 72426 75678 72440
rect 75612 72370 75617 72426
rect 75673 72370 75678 72426
rect 75612 72346 75619 72370
rect 75671 72346 75678 72370
rect 75612 72290 75617 72346
rect 75673 72290 75678 72346
rect 75612 72266 75619 72290
rect 75671 72266 75678 72290
rect 75612 72210 75617 72266
rect 75673 72210 75678 72266
rect 75612 72196 75619 72210
rect 75671 72196 75678 72210
rect 75612 72181 75678 72196
rect 76700 72760 76766 72775
rect 76700 72746 76707 72760
rect 76759 72746 76766 72760
rect 76700 72690 76705 72746
rect 76761 72690 76766 72746
rect 76700 72666 76707 72690
rect 76759 72666 76766 72690
rect 76700 72610 76705 72666
rect 76761 72610 76766 72666
rect 76700 72586 76707 72610
rect 76759 72586 76766 72610
rect 76700 72530 76705 72586
rect 76761 72530 76766 72586
rect 76700 72516 76707 72530
rect 76759 72516 76766 72530
rect 76700 72506 76766 72516
rect 76700 72450 76705 72506
rect 76761 72450 76766 72506
rect 76700 72440 76766 72450
rect 76700 72426 76707 72440
rect 76759 72426 76766 72440
rect 76700 72370 76705 72426
rect 76761 72370 76766 72426
rect 76700 72346 76707 72370
rect 76759 72346 76766 72370
rect 76700 72290 76705 72346
rect 76761 72290 76766 72346
rect 76700 72266 76707 72290
rect 76759 72266 76766 72290
rect 76700 72210 76705 72266
rect 76761 72210 76766 72266
rect 76700 72196 76707 72210
rect 76759 72196 76766 72210
rect 76700 72181 76766 72196
rect 77788 72760 77854 72775
rect 77788 72746 77795 72760
rect 77847 72746 77854 72760
rect 77788 72690 77793 72746
rect 77849 72690 77854 72746
rect 77788 72666 77795 72690
rect 77847 72666 77854 72690
rect 77788 72610 77793 72666
rect 77849 72610 77854 72666
rect 77788 72586 77795 72610
rect 77847 72586 77854 72610
rect 77788 72530 77793 72586
rect 77849 72530 77854 72586
rect 77788 72516 77795 72530
rect 77847 72516 77854 72530
rect 77788 72506 77854 72516
rect 77788 72450 77793 72506
rect 77849 72450 77854 72506
rect 77788 72440 77854 72450
rect 77788 72426 77795 72440
rect 77847 72426 77854 72440
rect 77788 72370 77793 72426
rect 77849 72370 77854 72426
rect 77788 72346 77795 72370
rect 77847 72346 77854 72370
rect 77788 72290 77793 72346
rect 77849 72290 77854 72346
rect 77788 72266 77795 72290
rect 77847 72266 77854 72290
rect 77788 72210 77793 72266
rect 77849 72210 77854 72266
rect 77788 72196 77795 72210
rect 77847 72196 77854 72210
rect 77788 72181 77854 72196
rect 78876 72760 78942 72775
rect 78876 72746 78883 72760
rect 78935 72746 78942 72760
rect 78876 72690 78881 72746
rect 78937 72690 78942 72746
rect 78876 72666 78883 72690
rect 78935 72666 78942 72690
rect 78876 72610 78881 72666
rect 78937 72610 78942 72666
rect 78876 72586 78883 72610
rect 78935 72586 78942 72610
rect 78876 72530 78881 72586
rect 78937 72530 78942 72586
rect 78876 72516 78883 72530
rect 78935 72516 78942 72530
rect 78876 72506 78942 72516
rect 78876 72450 78881 72506
rect 78937 72450 78942 72506
rect 78876 72440 78942 72450
rect 78876 72426 78883 72440
rect 78935 72426 78942 72440
rect 78876 72370 78881 72426
rect 78937 72370 78942 72426
rect 78876 72346 78883 72370
rect 78935 72346 78942 72370
rect 78876 72290 78881 72346
rect 78937 72290 78942 72346
rect 78876 72266 78883 72290
rect 78935 72266 78942 72290
rect 78876 72210 78881 72266
rect 78937 72210 78942 72266
rect 78876 72196 78883 72210
rect 78935 72196 78942 72210
rect 78876 72181 78942 72196
rect 79964 72760 80030 72775
rect 79964 72746 79971 72760
rect 80023 72746 80030 72760
rect 79964 72690 79969 72746
rect 80025 72690 80030 72746
rect 79964 72666 79971 72690
rect 80023 72666 80030 72690
rect 79964 72610 79969 72666
rect 80025 72610 80030 72666
rect 79964 72586 79971 72610
rect 80023 72586 80030 72610
rect 79964 72530 79969 72586
rect 80025 72530 80030 72586
rect 79964 72516 79971 72530
rect 80023 72516 80030 72530
rect 79964 72506 80030 72516
rect 79964 72450 79969 72506
rect 80025 72450 80030 72506
rect 79964 72440 80030 72450
rect 79964 72426 79971 72440
rect 80023 72426 80030 72440
rect 79964 72370 79969 72426
rect 80025 72370 80030 72426
rect 79964 72346 79971 72370
rect 80023 72346 80030 72370
rect 79964 72290 79969 72346
rect 80025 72290 80030 72346
rect 79964 72266 79971 72290
rect 80023 72266 80030 72290
rect 79964 72210 79969 72266
rect 80025 72210 80030 72266
rect 79964 72196 79971 72210
rect 80023 72196 80030 72210
rect 79964 72181 80030 72196
rect 81052 72760 81118 72775
rect 81052 72746 81059 72760
rect 81111 72746 81118 72760
rect 81052 72690 81057 72746
rect 81113 72690 81118 72746
rect 81052 72666 81059 72690
rect 81111 72666 81118 72690
rect 81052 72610 81057 72666
rect 81113 72610 81118 72666
rect 81052 72586 81059 72610
rect 81111 72586 81118 72610
rect 81052 72530 81057 72586
rect 81113 72530 81118 72586
rect 81052 72516 81059 72530
rect 81111 72516 81118 72530
rect 81052 72506 81118 72516
rect 81052 72450 81057 72506
rect 81113 72450 81118 72506
rect 81052 72440 81118 72450
rect 81052 72426 81059 72440
rect 81111 72426 81118 72440
rect 81052 72370 81057 72426
rect 81113 72370 81118 72426
rect 81052 72346 81059 72370
rect 81111 72346 81118 72370
rect 81052 72290 81057 72346
rect 81113 72290 81118 72346
rect 81052 72266 81059 72290
rect 81111 72266 81118 72290
rect 81052 72210 81057 72266
rect 81113 72210 81118 72266
rect 81052 72196 81059 72210
rect 81111 72196 81118 72210
rect 81052 72181 81118 72196
rect 86492 72760 86558 72775
rect 86492 72746 86499 72760
rect 86551 72746 86558 72760
rect 86492 72690 86497 72746
rect 86553 72690 86558 72746
rect 86492 72666 86499 72690
rect 86551 72666 86558 72690
rect 86492 72610 86497 72666
rect 86553 72610 86558 72666
rect 86492 72586 86499 72610
rect 86551 72586 86558 72610
rect 86492 72530 86497 72586
rect 86553 72530 86558 72586
rect 86492 72516 86499 72530
rect 86551 72516 86558 72530
rect 86492 72506 86558 72516
rect 86492 72450 86497 72506
rect 86553 72450 86558 72506
rect 86492 72440 86558 72450
rect 86492 72426 86499 72440
rect 86551 72426 86558 72440
rect 86492 72370 86497 72426
rect 86553 72370 86558 72426
rect 86492 72346 86499 72370
rect 86551 72346 86558 72370
rect 86492 72290 86497 72346
rect 86553 72290 86558 72346
rect 86492 72266 86499 72290
rect 86551 72266 86558 72290
rect 86492 72210 86497 72266
rect 86553 72210 86558 72266
rect 86492 72196 86499 72210
rect 86551 72196 86558 72210
rect 86492 72181 86558 72196
rect 87580 72760 87646 72775
rect 87580 72746 87587 72760
rect 87639 72746 87646 72760
rect 87580 72690 87585 72746
rect 87641 72690 87646 72746
rect 87580 72666 87587 72690
rect 87639 72666 87646 72690
rect 87580 72610 87585 72666
rect 87641 72610 87646 72666
rect 87580 72586 87587 72610
rect 87639 72586 87646 72610
rect 87580 72530 87585 72586
rect 87641 72530 87646 72586
rect 87580 72516 87587 72530
rect 87639 72516 87646 72530
rect 87580 72506 87646 72516
rect 87580 72450 87585 72506
rect 87641 72450 87646 72506
rect 87580 72440 87646 72450
rect 87580 72426 87587 72440
rect 87639 72426 87646 72440
rect 87580 72370 87585 72426
rect 87641 72370 87646 72426
rect 87580 72346 87587 72370
rect 87639 72346 87646 72370
rect 87580 72290 87585 72346
rect 87641 72290 87646 72346
rect 87580 72266 87587 72290
rect 87639 72266 87646 72290
rect 87580 72210 87585 72266
rect 87641 72210 87646 72266
rect 87580 72196 87587 72210
rect 87639 72196 87646 72210
rect 87580 72181 87646 72196
rect 88668 72760 88734 72775
rect 88668 72746 88675 72760
rect 88727 72746 88734 72760
rect 88668 72690 88673 72746
rect 88729 72690 88734 72746
rect 88668 72666 88675 72690
rect 88727 72666 88734 72690
rect 88668 72610 88673 72666
rect 88729 72610 88734 72666
rect 88668 72586 88675 72610
rect 88727 72586 88734 72610
rect 88668 72530 88673 72586
rect 88729 72530 88734 72586
rect 88668 72516 88675 72530
rect 88727 72516 88734 72530
rect 88668 72506 88734 72516
rect 88668 72450 88673 72506
rect 88729 72450 88734 72506
rect 88668 72440 88734 72450
rect 88668 72426 88675 72440
rect 88727 72426 88734 72440
rect 88668 72370 88673 72426
rect 88729 72370 88734 72426
rect 88668 72346 88675 72370
rect 88727 72346 88734 72370
rect 88668 72290 88673 72346
rect 88729 72290 88734 72346
rect 88668 72266 88675 72290
rect 88727 72266 88734 72290
rect 88668 72210 88673 72266
rect 88729 72210 88734 72266
rect 88668 72196 88675 72210
rect 88727 72196 88734 72210
rect 88668 72181 88734 72196
rect 67271 71660 67310 71662
rect 67606 71660 67645 71662
rect 67271 71629 67645 71660
rect 75069 70757 75135 70772
rect 75069 70743 75076 70757
rect 75128 70743 75135 70757
rect 75069 70687 75074 70743
rect 75130 70687 75135 70743
rect 75069 70663 75076 70687
rect 75128 70663 75135 70687
rect 75069 70607 75074 70663
rect 75130 70607 75135 70663
rect 75069 70583 75076 70607
rect 75128 70583 75135 70607
rect 75069 70527 75074 70583
rect 75130 70527 75135 70583
rect 75069 70513 75076 70527
rect 75128 70513 75135 70527
rect 75069 70503 75135 70513
rect 75069 70447 75074 70503
rect 75130 70447 75135 70503
rect 75069 70437 75135 70447
rect 75069 70423 75076 70437
rect 75128 70423 75135 70437
rect 75069 70367 75074 70423
rect 75130 70367 75135 70423
rect 75069 70343 75076 70367
rect 75128 70343 75135 70367
rect 51170 70294 51372 70306
rect 51170 63842 51181 70294
rect 51361 63842 51372 70294
rect 75069 70287 75074 70343
rect 75130 70287 75135 70343
rect 75069 70263 75076 70287
rect 75128 70263 75135 70287
rect 75069 70207 75074 70263
rect 75130 70207 75135 70263
rect 75069 70193 75076 70207
rect 75128 70193 75135 70207
rect 75069 70178 75135 70193
rect 76157 70757 76223 70772
rect 76157 70743 76164 70757
rect 76216 70743 76223 70757
rect 76157 70687 76162 70743
rect 76218 70687 76223 70743
rect 76157 70663 76164 70687
rect 76216 70663 76223 70687
rect 76157 70607 76162 70663
rect 76218 70607 76223 70663
rect 76157 70583 76164 70607
rect 76216 70583 76223 70607
rect 76157 70527 76162 70583
rect 76218 70527 76223 70583
rect 76157 70513 76164 70527
rect 76216 70513 76223 70527
rect 76157 70503 76223 70513
rect 76157 70447 76162 70503
rect 76218 70447 76223 70503
rect 76157 70437 76223 70447
rect 76157 70423 76164 70437
rect 76216 70423 76223 70437
rect 76157 70367 76162 70423
rect 76218 70367 76223 70423
rect 76157 70343 76164 70367
rect 76216 70343 76223 70367
rect 76157 70287 76162 70343
rect 76218 70287 76223 70343
rect 76157 70263 76164 70287
rect 76216 70263 76223 70287
rect 76157 70207 76162 70263
rect 76218 70207 76223 70263
rect 76157 70193 76164 70207
rect 76216 70193 76223 70207
rect 76157 70178 76223 70193
rect 77245 70757 77311 70772
rect 77245 70743 77252 70757
rect 77304 70743 77311 70757
rect 77245 70687 77250 70743
rect 77306 70687 77311 70743
rect 77245 70663 77252 70687
rect 77304 70663 77311 70687
rect 77245 70607 77250 70663
rect 77306 70607 77311 70663
rect 77245 70583 77252 70607
rect 77304 70583 77311 70607
rect 77245 70527 77250 70583
rect 77306 70527 77311 70583
rect 77245 70513 77252 70527
rect 77304 70513 77311 70527
rect 77245 70503 77311 70513
rect 77245 70447 77250 70503
rect 77306 70447 77311 70503
rect 77245 70437 77311 70447
rect 77245 70423 77252 70437
rect 77304 70423 77311 70437
rect 77245 70367 77250 70423
rect 77306 70367 77311 70423
rect 77245 70343 77252 70367
rect 77304 70343 77311 70367
rect 77245 70287 77250 70343
rect 77306 70287 77311 70343
rect 77245 70263 77252 70287
rect 77304 70263 77311 70287
rect 77245 70207 77250 70263
rect 77306 70207 77311 70263
rect 77245 70193 77252 70207
rect 77304 70193 77311 70207
rect 77245 70178 77311 70193
rect 78333 70757 78399 70772
rect 78333 70743 78340 70757
rect 78392 70743 78399 70757
rect 78333 70687 78338 70743
rect 78394 70687 78399 70743
rect 78333 70663 78340 70687
rect 78392 70663 78399 70687
rect 78333 70607 78338 70663
rect 78394 70607 78399 70663
rect 78333 70583 78340 70607
rect 78392 70583 78399 70607
rect 78333 70527 78338 70583
rect 78394 70527 78399 70583
rect 78333 70513 78340 70527
rect 78392 70513 78399 70527
rect 78333 70503 78399 70513
rect 78333 70447 78338 70503
rect 78394 70447 78399 70503
rect 78333 70437 78399 70447
rect 78333 70423 78340 70437
rect 78392 70423 78399 70437
rect 78333 70367 78338 70423
rect 78394 70367 78399 70423
rect 78333 70343 78340 70367
rect 78392 70343 78399 70367
rect 78333 70287 78338 70343
rect 78394 70287 78399 70343
rect 78333 70263 78340 70287
rect 78392 70263 78399 70287
rect 78333 70207 78338 70263
rect 78394 70207 78399 70263
rect 78333 70193 78340 70207
rect 78392 70193 78399 70207
rect 78333 70178 78399 70193
rect 79421 70757 79487 70772
rect 79421 70743 79428 70757
rect 79480 70743 79487 70757
rect 79421 70687 79426 70743
rect 79482 70687 79487 70743
rect 79421 70663 79428 70687
rect 79480 70663 79487 70687
rect 79421 70607 79426 70663
rect 79482 70607 79487 70663
rect 79421 70583 79428 70607
rect 79480 70583 79487 70607
rect 79421 70527 79426 70583
rect 79482 70527 79487 70583
rect 79421 70513 79428 70527
rect 79480 70513 79487 70527
rect 79421 70503 79487 70513
rect 79421 70447 79426 70503
rect 79482 70447 79487 70503
rect 79421 70437 79487 70447
rect 79421 70423 79428 70437
rect 79480 70423 79487 70437
rect 79421 70367 79426 70423
rect 79482 70367 79487 70423
rect 79421 70343 79428 70367
rect 79480 70343 79487 70367
rect 79421 70287 79426 70343
rect 79482 70287 79487 70343
rect 79421 70263 79428 70287
rect 79480 70263 79487 70287
rect 79421 70207 79426 70263
rect 79482 70207 79487 70263
rect 79421 70193 79428 70207
rect 79480 70193 79487 70207
rect 79421 70178 79487 70193
rect 81597 70757 81663 70772
rect 81597 70743 81604 70757
rect 81656 70743 81663 70757
rect 81597 70687 81602 70743
rect 81658 70687 81663 70743
rect 81597 70663 81604 70687
rect 81656 70663 81663 70687
rect 81597 70607 81602 70663
rect 81658 70607 81663 70663
rect 81597 70583 81604 70607
rect 81656 70583 81663 70607
rect 81597 70527 81602 70583
rect 81658 70527 81663 70583
rect 81597 70513 81604 70527
rect 81656 70513 81663 70527
rect 81597 70503 81663 70513
rect 81597 70447 81602 70503
rect 81658 70447 81663 70503
rect 81597 70437 81663 70447
rect 81597 70423 81604 70437
rect 81656 70423 81663 70437
rect 81597 70367 81602 70423
rect 81658 70367 81663 70423
rect 81597 70343 81604 70367
rect 81656 70343 81663 70367
rect 81597 70287 81602 70343
rect 81658 70287 81663 70343
rect 81597 70263 81604 70287
rect 81656 70263 81663 70287
rect 81597 70207 81602 70263
rect 81658 70207 81663 70263
rect 81597 70193 81604 70207
rect 81656 70193 81663 70207
rect 81597 70178 81663 70193
rect 82685 70757 82751 70772
rect 82685 70743 82692 70757
rect 82744 70743 82751 70757
rect 82685 70687 82690 70743
rect 82746 70687 82751 70743
rect 82685 70663 82692 70687
rect 82744 70663 82751 70687
rect 82685 70607 82690 70663
rect 82746 70607 82751 70663
rect 82685 70583 82692 70607
rect 82744 70583 82751 70607
rect 82685 70527 82690 70583
rect 82746 70527 82751 70583
rect 82685 70513 82692 70527
rect 82744 70513 82751 70527
rect 82685 70503 82751 70513
rect 82685 70447 82690 70503
rect 82746 70447 82751 70503
rect 82685 70437 82751 70447
rect 82685 70423 82692 70437
rect 82744 70423 82751 70437
rect 82685 70367 82690 70423
rect 82746 70367 82751 70423
rect 82685 70343 82692 70367
rect 82744 70343 82751 70367
rect 82685 70287 82690 70343
rect 82746 70287 82751 70343
rect 82685 70263 82692 70287
rect 82744 70263 82751 70287
rect 82685 70207 82690 70263
rect 82746 70207 82751 70263
rect 82685 70193 82692 70207
rect 82744 70193 82751 70207
rect 82685 70178 82751 70193
rect 83773 70757 83839 70772
rect 83773 70743 83780 70757
rect 83832 70743 83839 70757
rect 83773 70687 83778 70743
rect 83834 70687 83839 70743
rect 83773 70663 83780 70687
rect 83832 70663 83839 70687
rect 83773 70607 83778 70663
rect 83834 70607 83839 70663
rect 83773 70583 83780 70607
rect 83832 70583 83839 70607
rect 83773 70527 83778 70583
rect 83834 70527 83839 70583
rect 83773 70513 83780 70527
rect 83832 70513 83839 70527
rect 83773 70503 83839 70513
rect 83773 70447 83778 70503
rect 83834 70447 83839 70503
rect 83773 70437 83839 70447
rect 83773 70423 83780 70437
rect 83832 70423 83839 70437
rect 83773 70367 83778 70423
rect 83834 70367 83839 70423
rect 83773 70343 83780 70367
rect 83832 70343 83839 70367
rect 83773 70287 83778 70343
rect 83834 70287 83839 70343
rect 83773 70263 83780 70287
rect 83832 70263 83839 70287
rect 83773 70207 83778 70263
rect 83834 70207 83839 70263
rect 83773 70193 83780 70207
rect 83832 70193 83839 70207
rect 83773 70178 83839 70193
rect 84861 70757 84927 70772
rect 84861 70743 84868 70757
rect 84920 70743 84927 70757
rect 84861 70687 84866 70743
rect 84922 70687 84927 70743
rect 84861 70663 84868 70687
rect 84920 70663 84927 70687
rect 84861 70607 84866 70663
rect 84922 70607 84927 70663
rect 84861 70583 84868 70607
rect 84920 70583 84927 70607
rect 84861 70527 84866 70583
rect 84922 70527 84927 70583
rect 84861 70513 84868 70527
rect 84920 70513 84927 70527
rect 84861 70503 84927 70513
rect 84861 70447 84866 70503
rect 84922 70447 84927 70503
rect 84861 70437 84927 70447
rect 84861 70423 84868 70437
rect 84920 70423 84927 70437
rect 84861 70367 84866 70423
rect 84922 70367 84927 70423
rect 84861 70343 84868 70367
rect 84920 70343 84927 70367
rect 84861 70287 84866 70343
rect 84922 70287 84927 70343
rect 84861 70263 84868 70287
rect 84920 70263 84927 70287
rect 84861 70207 84866 70263
rect 84922 70207 84927 70263
rect 84861 70193 84868 70207
rect 84920 70193 84927 70207
rect 84861 70178 84927 70193
rect 85949 70757 86015 70772
rect 85949 70743 85956 70757
rect 86008 70743 86015 70757
rect 85949 70687 85954 70743
rect 86010 70687 86015 70743
rect 85949 70663 85956 70687
rect 86008 70663 86015 70687
rect 85949 70607 85954 70663
rect 86010 70607 86015 70663
rect 85949 70583 85956 70607
rect 86008 70583 86015 70607
rect 85949 70527 85954 70583
rect 86010 70527 86015 70583
rect 85949 70513 85956 70527
rect 86008 70513 86015 70527
rect 85949 70503 86015 70513
rect 85949 70447 85954 70503
rect 86010 70447 86015 70503
rect 85949 70437 86015 70447
rect 85949 70423 85956 70437
rect 86008 70423 86015 70437
rect 85949 70367 85954 70423
rect 86010 70367 86015 70423
rect 85949 70343 85956 70367
rect 86008 70343 86015 70367
rect 85949 70287 85954 70343
rect 86010 70287 86015 70343
rect 85949 70263 85956 70287
rect 86008 70263 86015 70287
rect 85949 70207 85954 70263
rect 86010 70207 86015 70263
rect 85949 70193 85956 70207
rect 86008 70193 86015 70207
rect 85949 70178 86015 70193
rect 87037 70757 87103 70772
rect 87037 70743 87044 70757
rect 87096 70743 87103 70757
rect 87037 70687 87042 70743
rect 87098 70687 87103 70743
rect 87037 70663 87044 70687
rect 87096 70663 87103 70687
rect 87037 70607 87042 70663
rect 87098 70607 87103 70663
rect 87037 70583 87044 70607
rect 87096 70583 87103 70607
rect 87037 70527 87042 70583
rect 87098 70527 87103 70583
rect 87037 70513 87044 70527
rect 87096 70513 87103 70527
rect 87037 70503 87103 70513
rect 87037 70447 87042 70503
rect 87098 70447 87103 70503
rect 87037 70437 87103 70447
rect 87037 70423 87044 70437
rect 87096 70423 87103 70437
rect 87037 70367 87042 70423
rect 87098 70367 87103 70423
rect 87037 70343 87044 70367
rect 87096 70343 87103 70367
rect 87037 70287 87042 70343
rect 87098 70287 87103 70343
rect 87037 70263 87044 70287
rect 87096 70263 87103 70287
rect 87037 70207 87042 70263
rect 87098 70207 87103 70263
rect 87037 70193 87044 70207
rect 87096 70193 87103 70207
rect 87037 70178 87103 70193
rect 88125 70757 88191 70772
rect 88125 70743 88132 70757
rect 88184 70743 88191 70757
rect 88125 70687 88130 70743
rect 88186 70687 88191 70743
rect 88125 70663 88132 70687
rect 88184 70663 88191 70687
rect 88125 70607 88130 70663
rect 88186 70607 88191 70663
rect 88125 70583 88132 70607
rect 88184 70583 88191 70607
rect 88125 70527 88130 70583
rect 88186 70527 88191 70583
rect 88125 70513 88132 70527
rect 88184 70513 88191 70527
rect 88125 70503 88191 70513
rect 88125 70447 88130 70503
rect 88186 70447 88191 70503
rect 88125 70437 88191 70447
rect 88125 70423 88132 70437
rect 88184 70423 88191 70437
rect 88125 70367 88130 70423
rect 88186 70367 88191 70423
rect 88125 70343 88132 70367
rect 88184 70343 88191 70367
rect 88125 70287 88130 70343
rect 88186 70287 88191 70343
rect 97683 70393 97747 70407
rect 97683 70337 97687 70393
rect 97743 70337 97747 70393
rect 97683 70323 97747 70337
rect 88125 70263 88132 70287
rect 88184 70263 88191 70287
rect 88125 70207 88130 70263
rect 88186 70207 88191 70263
rect 88125 70193 88132 70207
rect 88184 70193 88191 70207
rect 88125 70178 88191 70193
rect 67274 70149 67645 70160
rect 57438 69865 57652 69876
rect 57438 68341 57455 69865
rect 57635 68341 57652 69865
rect 57438 68330 57652 68341
rect 57446 65403 57606 65415
rect 57446 65389 57468 65403
rect 57584 65389 57606 65403
rect 57446 63893 57458 65389
rect 57594 63893 57606 65389
rect 57446 63879 57468 63893
rect 57584 63879 57606 63893
rect 67274 63889 67305 70149
rect 67613 63889 67645 70149
rect 75339 69766 75403 69780
rect 75339 69710 75343 69766
rect 75399 69710 75403 69766
rect 75339 69696 75403 69710
rect 75885 69766 75949 69780
rect 75885 69710 75889 69766
rect 75945 69710 75949 69766
rect 75885 69696 75949 69710
rect 76431 69757 76495 69771
rect 76431 69701 76435 69757
rect 76491 69701 76495 69757
rect 76431 69687 76495 69701
rect 76976 69756 77040 69770
rect 76976 69700 76980 69756
rect 77036 69700 77040 69756
rect 76976 69686 77040 69700
rect 78607 69744 78671 69758
rect 78607 69688 78611 69744
rect 78667 69688 78671 69744
rect 78607 69674 78671 69688
rect 79150 69741 79214 69755
rect 79150 69685 79154 69741
rect 79210 69685 79214 69741
rect 79150 69671 79214 69685
rect 79692 69740 79756 69754
rect 79692 69684 79696 69740
rect 79752 69684 79756 69740
rect 79692 69670 79756 69684
rect 80239 69745 80303 69759
rect 80239 69689 80243 69745
rect 80299 69689 80303 69745
rect 80239 69675 80303 69689
rect 82957 69756 83021 69770
rect 82957 69700 82961 69756
rect 83017 69700 83021 69756
rect 82957 69686 83021 69700
rect 83500 69760 83564 69774
rect 83500 69704 83504 69760
rect 83560 69704 83564 69760
rect 83500 69690 83564 69704
rect 84042 69754 84106 69768
rect 84042 69698 84046 69754
rect 84102 69698 84106 69754
rect 84042 69684 84106 69698
rect 84599 69745 84663 69759
rect 84599 69689 84603 69745
rect 84659 69689 84663 69745
rect 84599 69675 84663 69689
rect 86223 69756 86287 69770
rect 86223 69700 86227 69756
rect 86283 69700 86287 69756
rect 86223 69686 86287 69700
rect 86767 69749 86831 69763
rect 86767 69693 86771 69749
rect 86827 69693 86831 69749
rect 86767 69679 86831 69693
rect 87317 69753 87381 69767
rect 87317 69697 87321 69753
rect 87377 69697 87381 69753
rect 87317 69683 87381 69697
rect 87850 69753 87914 69767
rect 87850 69697 87854 69753
rect 87910 69697 87914 69753
rect 87850 69683 87914 69697
rect 96651 68909 96715 68923
rect 96651 68853 96655 68909
rect 96711 68853 96715 68909
rect 96651 68839 96715 68853
rect 97689 68852 97741 70323
rect 98240 69837 98304 69851
rect 98240 69781 98244 69837
rect 98300 69781 98304 69837
rect 98240 69767 98304 69781
rect 98082 69009 98146 69023
rect 98082 68953 98086 69009
rect 98142 68953 98146 69009
rect 98082 68939 98146 68953
rect 96651 68719 96715 68733
rect 96651 68663 96655 68719
rect 96711 68663 96715 68719
rect 96651 68649 96715 68663
rect 96651 67759 96715 67773
rect 96651 67703 96655 67759
rect 96711 67703 96715 67759
rect 96651 67689 96715 67703
rect 97689 67702 97741 68800
rect 98089 68841 98141 68939
rect 97988 68784 98040 68794
rect 98089 68779 98141 68789
rect 98246 68845 98298 69767
rect 101848 69090 102400 69106
rect 101848 69034 101856 69090
rect 101912 69088 101936 69090
rect 101992 69088 102016 69090
rect 102072 69088 102096 69090
rect 102152 69088 102176 69090
rect 102232 69088 102256 69090
rect 102312 69088 102336 69090
rect 101926 69036 101936 69088
rect 101992 69036 102002 69088
rect 102246 69036 102256 69088
rect 102312 69036 102322 69088
rect 101912 69034 101936 69036
rect 101992 69034 102016 69036
rect 102072 69034 102096 69036
rect 102152 69034 102176 69036
rect 102232 69034 102256 69036
rect 102312 69034 102336 69036
rect 102392 69034 102400 69090
rect 101848 69019 102400 69034
rect 97988 68639 98040 68732
rect 97982 68625 98046 68639
rect 97982 68569 97986 68625
rect 98042 68569 98046 68625
rect 97982 68555 98046 68569
rect 98082 67859 98146 67873
rect 98082 67803 98086 67859
rect 98142 67803 98146 67859
rect 98082 67789 98146 67803
rect 97689 67640 97741 67650
rect 98089 67691 98141 67789
rect 97988 67634 98040 67644
rect 96651 67569 96715 67583
rect 96651 67513 96655 67569
rect 96711 67513 96715 67569
rect 96651 67499 96715 67513
rect 98089 67629 98141 67639
rect 98246 67695 98298 68793
rect 103388 68951 103624 68971
rect 103388 68735 103398 68951
rect 103614 68735 103624 68951
rect 103388 68715 103624 68735
rect 98610 68544 98968 68559
rect 98610 68542 98641 68544
rect 98697 68542 98721 68544
rect 98777 68542 98801 68544
rect 98857 68542 98881 68544
rect 98937 68542 98968 68544
rect 98610 68490 98635 68542
rect 98697 68490 98699 68542
rect 98879 68490 98881 68542
rect 98943 68490 98968 68542
rect 98610 68488 98641 68490
rect 98697 68488 98721 68490
rect 98777 68488 98801 68490
rect 98857 68488 98881 68490
rect 98937 68488 98968 68490
rect 98610 68474 98968 68488
rect 101860 67939 102387 67957
rect 101860 67937 101895 67939
rect 101951 67937 101975 67939
rect 102031 67937 102055 67939
rect 102111 67937 102135 67939
rect 102191 67937 102215 67939
rect 102271 67937 102295 67939
rect 102351 67937 102387 67939
rect 101860 67885 101873 67937
rect 102053 67885 102055 67937
rect 102117 67885 102129 67937
rect 102191 67885 102193 67937
rect 102373 67885 102387 67937
rect 101860 67883 101895 67885
rect 101951 67883 101975 67885
rect 102031 67883 102055 67885
rect 102111 67883 102135 67885
rect 102191 67883 102215 67885
rect 102271 67883 102295 67885
rect 102351 67883 102387 67885
rect 101860 67866 102387 67883
rect 98246 67633 98298 67643
rect 103376 67800 103612 67820
rect 97988 67489 98040 67582
rect 103376 67584 103386 67800
rect 103602 67584 103612 67800
rect 103376 67564 103612 67584
rect 97982 67475 98046 67489
rect 97982 67419 97986 67475
rect 98042 67419 98046 67475
rect 97982 67405 98046 67419
rect 98608 67394 98966 67409
rect 98608 67392 98639 67394
rect 98695 67392 98719 67394
rect 98775 67392 98799 67394
rect 98855 67392 98879 67394
rect 98935 67392 98966 67394
rect 98608 67340 98633 67392
rect 98695 67340 98697 67392
rect 98877 67340 98879 67392
rect 98941 67340 98966 67392
rect 98608 67338 98639 67340
rect 98695 67338 98719 67340
rect 98775 67338 98799 67340
rect 98855 67338 98879 67340
rect 98935 67338 98966 67340
rect 98608 67324 98966 67338
rect 97683 66703 97747 66717
rect 97683 66647 97687 66703
rect 97743 66647 97747 66703
rect 97683 66633 97747 66647
rect 96651 65219 96715 65233
rect 96651 65163 96655 65219
rect 96711 65163 96715 65219
rect 96651 65149 96715 65163
rect 97689 65162 97741 66633
rect 98240 66147 98304 66161
rect 98240 66091 98244 66147
rect 98300 66091 98304 66147
rect 98240 66077 98304 66091
rect 98082 65319 98146 65333
rect 98082 65263 98086 65319
rect 98142 65263 98146 65319
rect 98082 65249 98146 65263
rect 96651 65029 96715 65043
rect 96651 64973 96655 65029
rect 96711 64973 96715 65029
rect 96651 64959 96715 64973
rect 67274 63879 67645 63889
rect 96651 63949 96715 63963
rect 96651 63893 96655 63949
rect 96711 63893 96715 63949
rect 96651 63879 96715 63893
rect 97689 63892 97741 65110
rect 98089 65151 98141 65249
rect 97988 65094 98040 65104
rect 98089 65089 98141 65099
rect 98246 65155 98298 66077
rect 101850 65397 102377 65415
rect 101850 65395 101885 65397
rect 101941 65395 101965 65397
rect 102021 65395 102045 65397
rect 102101 65395 102125 65397
rect 102181 65395 102205 65397
rect 102261 65395 102285 65397
rect 102341 65395 102377 65397
rect 101850 65343 101863 65395
rect 102043 65343 102045 65395
rect 102107 65343 102119 65395
rect 102181 65343 102183 65395
rect 102363 65343 102377 65395
rect 101850 65341 101885 65343
rect 101941 65341 101965 65343
rect 102021 65341 102045 65343
rect 102101 65341 102125 65343
rect 102181 65341 102205 65343
rect 102261 65341 102285 65343
rect 102341 65341 102377 65343
rect 101850 65324 102377 65341
rect 97988 64949 98040 65042
rect 97982 64935 98046 64949
rect 97982 64879 97986 64935
rect 98042 64879 98046 64935
rect 97982 64865 98046 64879
rect 98082 64049 98146 64063
rect 98082 63993 98086 64049
rect 98142 63993 98146 64049
rect 98082 63979 98146 63993
rect 51170 63831 51372 63842
rect 51410 63868 56946 63878
rect 51410 63846 51432 63868
rect 56924 63846 56946 63868
rect 57446 63867 57606 63879
rect 50105 63769 50111 63821
rect 50163 63769 50175 63821
rect 50227 63769 50233 63821
rect 50105 63753 50233 63769
rect 30017 63693 30032 63749
rect 30088 63693 30104 63749
rect 30017 63691 30104 63693
rect 30017 63669 30034 63691
rect 30086 63669 30104 63691
rect 51410 63710 51430 63846
rect 56926 63710 56946 63846
rect 97689 63830 97741 63840
rect 98089 63881 98141 63979
rect 97988 63824 98040 63834
rect 51410 63688 51432 63710
rect 56924 63688 56946 63710
rect 96651 63759 96715 63773
rect 96651 63703 96655 63759
rect 96711 63703 96715 63759
rect 96651 63689 96715 63703
rect 98089 63819 98141 63829
rect 98246 63885 98298 65103
rect 103234 65268 103470 65288
rect 103234 65052 103244 65268
rect 103460 65052 103470 65268
rect 103234 65032 103470 65052
rect 98526 64853 98884 64868
rect 98526 64851 98557 64853
rect 98613 64851 98637 64853
rect 98693 64851 98717 64853
rect 98773 64851 98797 64853
rect 98853 64851 98884 64853
rect 98526 64799 98551 64851
rect 98613 64799 98615 64851
rect 98795 64799 98797 64851
rect 98859 64799 98884 64851
rect 98526 64797 98557 64799
rect 98613 64797 98637 64799
rect 98693 64797 98717 64799
rect 98773 64797 98797 64799
rect 98853 64797 98884 64799
rect 98526 64783 98884 64797
rect 101850 64127 102377 64145
rect 101850 64125 101885 64127
rect 101941 64125 101965 64127
rect 102021 64125 102045 64127
rect 102101 64125 102125 64127
rect 102181 64125 102205 64127
rect 102261 64125 102285 64127
rect 102341 64125 102377 64127
rect 101850 64073 101863 64125
rect 102043 64073 102045 64125
rect 102107 64073 102119 64125
rect 102181 64073 102183 64125
rect 102363 64073 102377 64125
rect 101850 64071 101885 64073
rect 101941 64071 101965 64073
rect 102021 64071 102045 64073
rect 102101 64071 102125 64073
rect 102181 64071 102205 64073
rect 102261 64071 102285 64073
rect 102341 64071 102377 64073
rect 101850 64054 102377 64071
rect 98246 63823 98298 63833
rect 103205 63978 103441 63998
rect 51410 63678 56946 63688
rect 97988 63679 98040 63772
rect 103205 63762 103215 63978
rect 103431 63762 103441 63978
rect 103205 63742 103441 63762
rect 30017 63613 30032 63669
rect 30088 63613 30104 63669
rect 30017 63589 30034 63613
rect 30086 63589 30104 63613
rect 97982 63665 98046 63679
rect 97982 63609 97986 63665
rect 98042 63609 98046 63665
rect 97982 63595 98046 63609
rect 30017 63533 30032 63589
rect 30088 63533 30104 63589
rect 98524 63584 98882 63599
rect 98524 63582 98555 63584
rect 98611 63582 98635 63584
rect 98691 63582 98715 63584
rect 98771 63582 98795 63584
rect 98851 63582 98882 63584
rect 30017 63511 30034 63533
rect 30086 63511 30104 63533
rect 30017 63488 30104 63511
rect 38211 63542 38287 63569
rect 38211 63520 38223 63542
rect 38275 63520 38287 63542
rect 38211 63464 38221 63520
rect 38277 63464 38287 63520
rect 98524 63530 98549 63582
rect 98611 63530 98613 63582
rect 98793 63530 98795 63582
rect 98857 63530 98882 63582
rect 98524 63528 98555 63530
rect 98611 63528 98635 63530
rect 98691 63528 98715 63530
rect 98771 63528 98795 63530
rect 98851 63528 98882 63530
rect 98524 63514 98882 63528
rect 38211 63440 38223 63464
rect 38275 63440 38287 63464
rect 38211 63384 38221 63440
rect 38277 63384 38287 63440
rect 38211 63362 38223 63384
rect 38275 63362 38287 63384
rect 38211 63360 38287 63362
rect 38211 63304 38221 63360
rect 38277 63304 38287 63360
rect 38211 63298 38223 63304
rect 38275 63298 38287 63304
rect 38211 63286 38287 63298
rect 38211 63280 38223 63286
rect 38275 63280 38287 63286
rect 38211 63224 38221 63280
rect 38277 63224 38287 63280
rect 38211 63222 38287 63224
rect 38211 63200 38223 63222
rect 38275 63200 38287 63222
rect 25282 63172 25346 63198
rect 25282 63166 25288 63172
rect 25340 63166 25346 63172
rect 25282 63110 25286 63166
rect 25342 63110 25346 63166
rect 25282 63108 25346 63110
rect 25282 63086 25288 63108
rect 25340 63086 25346 63108
rect 25282 63030 25286 63086
rect 25342 63030 25346 63086
rect 25282 63006 25288 63030
rect 25340 63006 25346 63030
rect 25282 62950 25286 63006
rect 25342 62950 25346 63006
rect 25282 62928 25288 62950
rect 25340 62928 25346 62950
rect 25282 62926 25346 62928
rect 25282 62870 25286 62926
rect 25342 62870 25346 62926
rect 25282 62864 25288 62870
rect 25340 62864 25346 62870
rect 25282 62839 25346 62864
rect 30012 63140 30096 63152
rect 30012 63126 30028 63140
rect 30080 63126 30096 63140
rect 30012 63070 30026 63126
rect 30082 63070 30096 63126
rect 30012 63046 30028 63070
rect 30080 63046 30096 63070
rect 30012 62990 30026 63046
rect 30082 62990 30096 63046
rect 30012 62966 30028 62990
rect 30080 62966 30096 62990
rect 30012 62910 30026 62966
rect 30082 62910 30096 62966
rect 30012 62896 30028 62910
rect 30080 62896 30096 62910
rect 30012 62886 30096 62896
rect 30012 62830 30026 62886
rect 30082 62830 30096 62886
rect 30012 62820 30096 62830
rect 30012 62806 30028 62820
rect 30080 62806 30096 62820
rect 30012 62750 30026 62806
rect 30082 62750 30096 62806
rect 30012 62726 30028 62750
rect 30080 62726 30096 62750
rect 30012 62670 30026 62726
rect 30082 62670 30096 62726
rect 30012 62646 30028 62670
rect 30080 62646 30096 62670
rect 25283 62627 25347 62645
rect 25283 62571 25287 62627
rect 25343 62571 25347 62627
rect 25283 62565 25289 62571
rect 25341 62565 25347 62571
rect 25283 62553 25347 62565
rect 25283 62547 25289 62553
rect 25341 62547 25347 62553
rect 25283 62491 25287 62547
rect 25343 62491 25347 62547
rect 25283 62489 25347 62491
rect 25283 62467 25289 62489
rect 25341 62467 25347 62489
rect 25283 62411 25287 62467
rect 25343 62411 25347 62467
rect 30012 62590 30026 62646
rect 30082 62590 30096 62646
rect 30012 62576 30028 62590
rect 30080 62576 30096 62590
rect 30012 62566 30096 62576
rect 30012 62510 30026 62566
rect 30082 62510 30096 62566
rect 30012 62500 30096 62510
rect 30012 62486 30028 62500
rect 30080 62486 30096 62500
rect 25283 62387 25289 62411
rect 25341 62387 25347 62411
rect 25283 62331 25287 62387
rect 25343 62331 25347 62387
rect 27480 62431 27944 62445
rect 27480 62375 27484 62431
rect 27540 62429 27564 62431
rect 27620 62429 27644 62431
rect 27700 62429 27724 62431
rect 27780 62429 27804 62431
rect 27860 62429 27884 62431
rect 27546 62377 27558 62429
rect 27620 62377 27622 62429
rect 27802 62377 27804 62429
rect 27866 62377 27878 62429
rect 27540 62375 27564 62377
rect 27620 62375 27644 62377
rect 27700 62375 27724 62377
rect 27780 62375 27804 62377
rect 27860 62375 27884 62377
rect 27940 62375 27944 62431
rect 27480 62361 27944 62375
rect 30012 62430 30026 62486
rect 30082 62430 30096 62486
rect 30012 62406 30028 62430
rect 30080 62406 30096 62430
rect 25283 62309 25289 62331
rect 25341 62309 25347 62331
rect 25283 62307 25347 62309
rect 25283 62251 25287 62307
rect 25343 62251 25347 62307
rect 30012 62350 30026 62406
rect 30082 62350 30096 62406
rect 30012 62326 30028 62350
rect 30080 62326 30096 62350
rect 26064 62278 26193 62288
rect 25283 62245 25289 62251
rect 25341 62245 25347 62251
rect 25283 62233 25347 62245
rect 25283 62227 25289 62233
rect 25341 62227 25347 62233
rect 25283 62171 25287 62227
rect 25343 62171 25347 62227
rect 26047 62272 26209 62278
rect 26047 62220 26070 62272
rect 26122 62220 26134 62272
rect 26186 62220 26209 62272
rect 30012 62270 30026 62326
rect 30082 62270 30096 62326
rect 30012 62256 30028 62270
rect 30080 62256 30096 62270
rect 30012 62244 30096 62256
rect 38211 63144 38221 63200
rect 38277 63144 38287 63200
rect 38211 63120 38223 63144
rect 38275 63120 38287 63144
rect 38211 63064 38221 63120
rect 38277 63064 38287 63120
rect 38211 63042 38223 63064
rect 38275 63042 38287 63064
rect 38211 63040 38287 63042
rect 38211 62984 38221 63040
rect 38277 62984 38287 63040
rect 64176 63232 64412 63242
rect 69636 63232 69872 63242
rect 64176 63204 69872 63232
rect 64176 63024 64204 63204
rect 64384 63024 69664 63204
rect 69844 63024 69872 63204
rect 64176 62996 69872 63024
rect 64176 62986 64412 62996
rect 69636 62986 69872 62996
rect 38211 62978 38223 62984
rect 38275 62978 38287 62984
rect 38211 62966 38287 62978
rect 38211 62960 38223 62966
rect 38275 62960 38287 62966
rect 38211 62904 38221 62960
rect 38277 62904 38287 62960
rect 38211 62902 38287 62904
rect 38211 62880 38223 62902
rect 38275 62880 38287 62902
rect 38211 62824 38221 62880
rect 38277 62824 38287 62880
rect 58567 62896 58631 62910
rect 58567 62840 58571 62896
rect 58627 62840 58631 62896
rect 58567 62826 58631 62840
rect 59607 62891 59689 62913
rect 59607 62835 59620 62891
rect 59676 62835 59689 62891
rect 38211 62800 38223 62824
rect 38275 62800 38287 62824
rect 38211 62744 38221 62800
rect 38277 62744 38287 62800
rect 38211 62722 38223 62744
rect 38275 62722 38287 62744
rect 38211 62720 38287 62722
rect 38211 62664 38221 62720
rect 38277 62664 38287 62720
rect 38211 62658 38223 62664
rect 38275 62658 38287 62664
rect 38211 62646 38287 62658
rect 59607 62821 59622 62835
rect 59674 62821 59689 62835
rect 59607 62811 59689 62821
rect 59607 62755 59620 62811
rect 59676 62755 59689 62811
rect 59607 62745 59689 62755
rect 59607 62731 59622 62745
rect 59674 62731 59689 62745
rect 59607 62675 59620 62731
rect 59676 62675 59689 62731
rect 59607 62654 59689 62675
rect 38211 62640 38223 62646
rect 38275 62640 38287 62646
rect 38211 62584 38221 62640
rect 38277 62584 38287 62640
rect 57187 62588 57251 62598
rect 58324 62588 58388 62598
rect 38211 62582 38287 62584
rect 38211 62560 38223 62582
rect 38275 62560 38287 62582
rect 38211 62504 38221 62560
rect 38277 62504 38287 62560
rect 57181 62582 58388 62588
rect 57181 62530 57193 62582
rect 57245 62530 58330 62582
rect 58382 62530 58388 62582
rect 57181 62524 58388 62530
rect 57187 62514 57251 62524
rect 58324 62514 58388 62524
rect 59720 62590 59784 62600
rect 62455 62590 62519 62600
rect 59720 62584 62519 62590
rect 59720 62532 59726 62584
rect 59778 62532 62461 62584
rect 62513 62532 62519 62584
rect 59720 62526 62519 62532
rect 59720 62516 59784 62526
rect 62455 62516 62519 62526
rect 38211 62480 38223 62504
rect 38275 62480 38287 62504
rect 38211 62424 38221 62480
rect 38277 62424 38287 62480
rect 38211 62402 38223 62424
rect 38275 62402 38287 62424
rect 38211 62400 38287 62402
rect 38211 62344 38221 62400
rect 38277 62344 38287 62400
rect 38211 62338 38223 62344
rect 38275 62338 38287 62344
rect 38211 62326 38287 62338
rect 38211 62320 38223 62326
rect 38275 62320 38287 62326
rect 38211 62264 38221 62320
rect 38277 62264 38287 62320
rect 38211 62262 38287 62264
rect 26047 62214 26209 62220
rect 38211 62240 38223 62262
rect 38275 62240 38287 62262
rect 25283 62153 25347 62171
rect 21576 61580 21812 61600
rect 21576 61364 21586 61580
rect 21802 61364 21812 61580
rect 21576 61344 21812 61364
rect 26064 51945 26193 62214
rect 38211 62184 38221 62240
rect 38277 62184 38287 62240
rect 38211 62160 38223 62184
rect 38275 62160 38287 62184
rect 38211 62104 38221 62160
rect 38277 62104 38287 62160
rect 38211 62082 38223 62104
rect 38275 62082 38287 62104
rect 59609 62418 59708 62452
rect 59609 62362 59630 62418
rect 59686 62362 59708 62418
rect 59609 62352 59708 62362
rect 59609 62338 59632 62352
rect 59684 62338 59708 62352
rect 59609 62282 59630 62338
rect 59686 62282 59708 62338
rect 59609 62258 59632 62282
rect 59684 62258 59708 62282
rect 59609 62202 59630 62258
rect 59686 62202 59708 62258
rect 59609 62178 59632 62202
rect 59684 62178 59708 62202
rect 59609 62122 59630 62178
rect 59686 62122 59708 62178
rect 59609 62108 59632 62122
rect 59684 62108 59708 62122
rect 38211 62080 38287 62082
rect 38211 62024 38221 62080
rect 38277 62024 38287 62080
rect 38211 62018 38223 62024
rect 38275 62018 38287 62024
rect 38211 62006 38287 62018
rect 59090 62087 59154 62101
rect 59090 62031 59094 62087
rect 59150 62031 59154 62087
rect 59090 62017 59154 62031
rect 59609 62098 59708 62108
rect 62455 62177 62519 62187
rect 64330 62177 64394 62187
rect 62455 62171 64394 62177
rect 62455 62119 62461 62171
rect 62513 62119 64336 62171
rect 64388 62119 64394 62171
rect 62455 62113 64394 62119
rect 62455 62103 62519 62113
rect 64330 62103 64394 62113
rect 59609 62042 59630 62098
rect 59686 62042 59708 62098
rect 59609 62008 59708 62042
rect 38211 62000 38223 62006
rect 38275 62000 38287 62006
rect 38211 61944 38221 62000
rect 38277 61944 38287 62000
rect 38211 61942 38287 61944
rect 38211 61920 38223 61942
rect 38275 61920 38287 61942
rect 38211 61864 38221 61920
rect 38277 61864 38287 61920
rect 38211 61840 38223 61864
rect 38275 61840 38287 61864
rect 38211 61784 38221 61840
rect 38277 61784 38287 61840
rect 38211 61762 38223 61784
rect 38275 61762 38287 61784
rect 38211 61760 38287 61762
rect 38211 61704 38221 61760
rect 38277 61704 38287 61760
rect 38211 61698 38223 61704
rect 38275 61698 38287 61704
rect 38211 61686 38287 61698
rect 38211 61680 38223 61686
rect 38275 61680 38287 61686
rect 38211 61624 38221 61680
rect 38277 61624 38287 61680
rect 38211 61622 38287 61624
rect 38211 61600 38223 61622
rect 38275 61600 38287 61622
rect 38211 61544 38221 61600
rect 38277 61544 38287 61600
rect 57187 61673 57251 61683
rect 60521 61673 60585 61683
rect 66522 61673 66586 61683
rect 57187 61667 66586 61673
rect 57187 61615 57193 61667
rect 57245 61615 60527 61667
rect 60579 61615 66528 61667
rect 66580 61615 66586 61667
rect 57187 61609 66586 61615
rect 57187 61599 57251 61609
rect 60521 61599 60585 61609
rect 66522 61599 66586 61609
rect 38211 61520 38223 61544
rect 38275 61520 38287 61544
rect 26895 61497 27024 61518
rect 26877 61491 27039 61497
rect 26877 61439 26901 61491
rect 26953 61439 26965 61491
rect 27017 61439 27039 61491
rect 26877 61433 27039 61439
rect 38211 61464 38221 61520
rect 38277 61464 38287 61520
rect 38211 61442 38223 61464
rect 38275 61442 38287 61464
rect 38211 61440 38287 61442
rect 26895 53303 27024 61433
rect 30015 61373 30099 61385
rect 30015 61359 30031 61373
rect 30083 61359 30099 61373
rect 27442 61341 27951 61355
rect 27442 61339 27468 61341
rect 27524 61339 27548 61341
rect 27604 61339 27628 61341
rect 27684 61339 27708 61341
rect 27764 61339 27788 61341
rect 27844 61339 27868 61341
rect 27924 61339 27951 61341
rect 27442 61287 27446 61339
rect 27626 61287 27628 61339
rect 27690 61287 27702 61339
rect 27764 61287 27766 61339
rect 27946 61287 27951 61339
rect 27442 61285 27468 61287
rect 27524 61285 27548 61287
rect 27604 61285 27628 61287
rect 27684 61285 27708 61287
rect 27764 61285 27788 61287
rect 27844 61285 27868 61287
rect 27924 61285 27951 61287
rect 27442 61271 27951 61285
rect 30015 61303 30029 61359
rect 30085 61303 30099 61359
rect 30015 61279 30031 61303
rect 30083 61279 30099 61303
rect 30015 61223 30029 61279
rect 30085 61223 30099 61279
rect 30015 61199 30031 61223
rect 30083 61199 30099 61223
rect 30015 61143 30029 61199
rect 30085 61143 30099 61199
rect 30015 61129 30031 61143
rect 30083 61129 30099 61143
rect 30015 61119 30099 61129
rect 30015 61063 30029 61119
rect 30085 61063 30099 61119
rect 30015 61053 30099 61063
rect 30015 61039 30031 61053
rect 30083 61039 30099 61053
rect 30015 60983 30029 61039
rect 30085 60983 30099 61039
rect 30015 60959 30031 60983
rect 30083 60959 30099 60983
rect 30015 60903 30029 60959
rect 30085 60903 30099 60959
rect 30015 60879 30031 60903
rect 30083 60879 30099 60903
rect 30015 60823 30029 60879
rect 30085 60823 30099 60879
rect 30015 60809 30031 60823
rect 30083 60809 30099 60823
rect 30015 60799 30099 60809
rect 30015 60743 30029 60799
rect 30085 60743 30099 60799
rect 30015 60733 30099 60743
rect 30015 60719 30031 60733
rect 30083 60719 30099 60733
rect 30015 60663 30029 60719
rect 30085 60663 30099 60719
rect 30015 60639 30031 60663
rect 30083 60639 30099 60663
rect 30015 60583 30029 60639
rect 30085 60583 30099 60639
rect 30015 60559 30031 60583
rect 30083 60559 30099 60583
rect 30015 60503 30029 60559
rect 30085 60503 30099 60559
rect 30015 60489 30031 60503
rect 30083 60489 30099 60503
rect 30015 60477 30099 60489
rect 38211 61384 38221 61440
rect 38277 61384 38287 61440
rect 38211 61378 38223 61384
rect 38275 61378 38287 61384
rect 38211 61366 38287 61378
rect 38211 61360 38223 61366
rect 38275 61360 38287 61366
rect 38211 61304 38221 61360
rect 38277 61304 38287 61360
rect 38211 61302 38287 61304
rect 38211 61280 38223 61302
rect 38275 61280 38287 61302
rect 38211 61224 38221 61280
rect 38277 61224 38287 61280
rect 38211 61200 38223 61224
rect 38275 61200 38287 61224
rect 38211 61144 38221 61200
rect 38277 61144 38287 61200
rect 59738 61229 59802 61239
rect 62523 61229 62587 61239
rect 63795 61229 63859 61239
rect 59738 61223 63859 61229
rect 59262 61167 59326 61181
rect 38211 61122 38223 61144
rect 38275 61122 38287 61144
rect 38211 61120 38287 61122
rect 38211 61064 38221 61120
rect 38277 61064 38287 61120
rect 58567 61147 58631 61161
rect 58567 61091 58571 61147
rect 58627 61091 58631 61147
rect 58567 61077 58631 61091
rect 59262 61153 59268 61167
rect 59320 61153 59326 61167
rect 59738 61171 59744 61223
rect 59796 61171 62529 61223
rect 62581 61171 63801 61223
rect 63853 61171 63859 61223
rect 59738 61165 63859 61171
rect 59738 61155 59802 61165
rect 62523 61155 62587 61165
rect 63795 61155 63859 61165
rect 59262 61097 59266 61153
rect 59322 61097 59326 61153
rect 38211 61058 38223 61064
rect 38275 61058 38287 61064
rect 38211 61046 38287 61058
rect 38211 61040 38223 61046
rect 38275 61040 38287 61046
rect 38211 60984 38221 61040
rect 38277 60984 38287 61040
rect 38211 60982 38287 60984
rect 38211 60960 38223 60982
rect 38275 60960 38287 60982
rect 38211 60904 38221 60960
rect 38277 60904 38287 60960
rect 59262 61073 59268 61097
rect 59320 61073 59326 61097
rect 59262 61017 59266 61073
rect 59322 61017 59326 61073
rect 59262 60993 59268 61017
rect 59320 60993 59326 61017
rect 59262 60937 59266 60993
rect 59322 60937 59326 60993
rect 59262 60923 59268 60937
rect 59320 60923 59326 60937
rect 59262 60910 59326 60923
rect 38211 60880 38223 60904
rect 38275 60880 38287 60904
rect 38211 60824 38221 60880
rect 38277 60824 38287 60880
rect 57187 60838 57251 60848
rect 57977 60838 58041 60848
rect 38211 60802 38223 60824
rect 38275 60802 38287 60824
rect 38211 60800 38287 60802
rect 38211 60744 38221 60800
rect 38277 60744 38287 60800
rect 57184 60832 58041 60838
rect 57184 60780 57193 60832
rect 57245 60780 57983 60832
rect 58035 60780 58041 60832
rect 57184 60774 58041 60780
rect 57187 60764 57251 60774
rect 57977 60764 58041 60774
rect 38211 60738 38223 60744
rect 38275 60738 38287 60744
rect 38211 60726 38287 60738
rect 38211 60720 38223 60726
rect 38275 60720 38287 60726
rect 38211 60664 38221 60720
rect 38277 60664 38287 60720
rect 38211 60662 38287 60664
rect 38211 60640 38223 60662
rect 38275 60640 38287 60662
rect 38211 60584 38221 60640
rect 38277 60584 38287 60640
rect 38211 60560 38223 60584
rect 38275 60560 38287 60584
rect 38211 60504 38221 60560
rect 38277 60504 38287 60560
rect 38211 60482 38223 60504
rect 38275 60482 38287 60504
rect 38211 60480 38287 60482
rect 38211 60424 38221 60480
rect 38277 60424 38287 60480
rect 38211 60418 38223 60424
rect 38275 60418 38287 60424
rect 38211 60406 38287 60418
rect 38211 60400 38223 60406
rect 38275 60400 38287 60406
rect 38211 60344 38221 60400
rect 38277 60344 38287 60400
rect 59263 60669 59327 60700
rect 59263 60613 59267 60669
rect 59323 60613 59327 60669
rect 63439 60615 63503 60629
rect 63439 60613 63443 60615
rect 59263 60603 59327 60613
rect 59263 60589 59269 60603
rect 59321 60589 59327 60603
rect 59263 60533 59267 60589
rect 59323 60533 59327 60589
rect 59263 60509 59269 60533
rect 59321 60509 59327 60533
rect 59263 60453 59267 60509
rect 59323 60453 59327 60509
rect 59263 60429 59269 60453
rect 59321 60429 59327 60453
rect 59263 60373 59267 60429
rect 59323 60373 59327 60429
rect 59263 60359 59269 60373
rect 59321 60359 59327 60373
rect 38211 60342 38287 60344
rect 38211 60320 38223 60342
rect 38275 60320 38287 60342
rect 38211 60264 38221 60320
rect 38277 60264 38287 60320
rect 59090 60337 59154 60351
rect 59090 60281 59094 60337
rect 59150 60281 59154 60337
rect 59090 60267 59154 60281
rect 59263 60349 59327 60359
rect 59263 60293 59267 60349
rect 59323 60293 59327 60349
rect 38211 60240 38223 60264
rect 38275 60240 38287 60264
rect 59263 60262 59327 60293
rect 62032 60561 63443 60613
rect 30017 60164 30098 60192
rect 30017 60142 30031 60164
rect 30083 60142 30098 60164
rect 30017 60086 30029 60142
rect 30085 60086 30098 60142
rect 38211 60184 38221 60240
rect 38277 60184 38287 60240
rect 38211 60162 38223 60184
rect 38275 60162 38287 60184
rect 38211 60136 38287 60162
rect 30017 60062 30031 60086
rect 30083 60062 30098 60086
rect 30017 60006 30029 60062
rect 30085 60006 30098 60062
rect 60032 60109 60437 60120
rect 60032 60053 60046 60109
rect 60102 60107 60126 60109
rect 60182 60107 60206 60109
rect 60262 60107 60286 60109
rect 60342 60107 60366 60109
rect 60102 60055 60112 60107
rect 60356 60055 60366 60107
rect 60102 60053 60126 60055
rect 60182 60053 60206 60055
rect 60262 60053 60286 60055
rect 60342 60053 60366 60055
rect 60422 60053 60437 60109
rect 60032 60042 60437 60053
rect 60676 60112 60905 60126
rect 60676 60056 60682 60112
rect 60738 60110 60762 60112
rect 60818 60110 60842 60112
rect 60752 60058 60762 60110
rect 60818 60058 60828 60110
rect 60738 60056 60762 60058
rect 60818 60056 60842 60058
rect 60898 60056 60905 60112
rect 60676 60042 60905 60056
rect 30017 59984 30031 60006
rect 30083 59984 30098 60006
rect 30017 59982 30098 59984
rect 30017 59926 30029 59982
rect 30085 59926 30098 59982
rect 30017 59920 30031 59926
rect 30083 59920 30098 59926
rect 30017 59908 30098 59920
rect 30017 59902 30031 59908
rect 30083 59902 30098 59908
rect 30017 59846 30029 59902
rect 30085 59846 30098 59902
rect 62032 59885 62084 60561
rect 63439 60559 63443 60561
rect 63499 60613 63503 60615
rect 63499 60561 64898 60613
rect 63499 60559 63503 60561
rect 63439 60545 63503 60559
rect 63439 60271 63503 60285
rect 63439 60269 63443 60271
rect 63084 60217 63443 60269
rect 62149 60111 62445 60136
rect 62205 60109 62229 60111
rect 62285 60109 62309 60111
rect 62365 60109 62389 60111
rect 62227 60057 62229 60109
rect 62291 60057 62303 60109
rect 62365 60057 62367 60109
rect 62205 60055 62229 60057
rect 62285 60055 62309 60057
rect 62365 60055 62389 60057
rect 62149 60030 62445 60055
rect 62668 60112 62895 60129
rect 62668 60056 62673 60112
rect 62729 60110 62753 60112
rect 62809 60110 62833 60112
rect 62743 60058 62753 60110
rect 62809 60058 62819 60110
rect 62729 60056 62753 60058
rect 62809 60056 62833 60058
rect 62889 60056 62895 60112
rect 62668 60039 62895 60056
rect 63084 59991 63136 60217
rect 63439 60215 63443 60217
rect 63499 60269 63503 60271
rect 63499 60217 63834 60269
rect 63499 60215 63503 60217
rect 63439 60201 63503 60215
rect 62841 59939 63136 59991
rect 63782 59991 63834 60217
rect 64030 60104 64251 60121
rect 64030 60048 64032 60104
rect 64088 60102 64112 60104
rect 64168 60102 64192 60104
rect 64102 60050 64112 60102
rect 64168 60050 64178 60102
rect 64088 60048 64112 60050
rect 64168 60048 64192 60050
rect 64248 60048 64251 60104
rect 64030 60032 64251 60048
rect 64477 60111 64775 60126
rect 64477 60055 64478 60111
rect 64534 60109 64558 60111
rect 64614 60109 64638 60111
rect 64694 60109 64718 60111
rect 64556 60057 64558 60109
rect 64620 60057 64632 60109
rect 64694 60057 64696 60109
rect 64534 60055 64558 60057
rect 64614 60055 64638 60057
rect 64694 60055 64718 60057
rect 64774 60055 64775 60111
rect 64477 60040 64775 60055
rect 63782 59939 64083 59991
rect 64846 59963 64898 60561
rect 66015 60110 66442 60125
rect 66015 60054 66040 60110
rect 66096 60108 66120 60110
rect 66176 60108 66200 60110
rect 66256 60108 66280 60110
rect 66336 60108 66360 60110
rect 66096 60056 66106 60108
rect 66350 60056 66360 60108
rect 66096 60054 66120 60056
rect 66176 60054 66200 60056
rect 66256 60054 66280 60056
rect 66336 60054 66360 60056
rect 66416 60054 66442 60110
rect 66015 60040 66442 60054
rect 66669 60107 66896 60123
rect 66669 60051 66674 60107
rect 66730 60105 66754 60107
rect 66810 60105 66834 60107
rect 66744 60053 66754 60105
rect 66810 60053 66820 60105
rect 66730 60051 66754 60053
rect 66810 60051 66834 60053
rect 66890 60051 66896 60107
rect 66669 60035 66896 60051
rect 30017 59844 30098 59846
rect 30017 59822 30031 59844
rect 30083 59822 30098 59844
rect 30017 59766 30029 59822
rect 30085 59766 30098 59822
rect 30017 59742 30031 59766
rect 30083 59742 30098 59766
rect 30017 59686 30029 59742
rect 30085 59686 30098 59742
rect 30017 59664 30031 59686
rect 30083 59664 30098 59686
rect 30017 59662 30098 59664
rect 30017 59606 30029 59662
rect 30085 59606 30098 59662
rect 30017 59600 30031 59606
rect 30083 59600 30098 59606
rect 30017 59588 30098 59600
rect 30017 59582 30031 59588
rect 30083 59582 30098 59588
rect 30017 59526 30029 59582
rect 30085 59526 30098 59582
rect 30017 59524 30098 59526
rect 30017 59502 30031 59524
rect 30083 59502 30098 59524
rect 30017 59446 30029 59502
rect 30085 59446 30098 59502
rect 30017 59422 30031 59446
rect 30083 59422 30098 59446
rect 30017 59366 30029 59422
rect 30085 59366 30098 59422
rect 30017 59344 30031 59366
rect 30083 59344 30098 59366
rect 30017 59342 30098 59344
rect 30017 59286 30029 59342
rect 30085 59286 30098 59342
rect 30017 59280 30031 59286
rect 30083 59280 30098 59286
rect 30017 59268 30098 59280
rect 30017 59262 30031 59268
rect 30083 59262 30098 59268
rect 30017 59206 30029 59262
rect 30085 59206 30098 59262
rect 30017 59204 30098 59206
rect 30017 59182 30031 59204
rect 30083 59182 30098 59204
rect 30017 59126 30029 59182
rect 30085 59126 30098 59182
rect 30017 59102 30031 59126
rect 30083 59102 30098 59126
rect 30017 59046 30029 59102
rect 30085 59046 30098 59102
rect 30017 59024 30031 59046
rect 30083 59024 30098 59046
rect 30017 58997 30098 59024
rect 62524 59036 62588 59052
rect 62524 58984 62530 59036
rect 62582 58984 62588 59036
rect 30015 58704 30094 58723
rect 30015 58648 30026 58704
rect 30082 58648 30094 58704
rect 30015 58634 30028 58648
rect 30080 58634 30094 58648
rect 30015 58624 30094 58634
rect 47725 58694 47789 58708
rect 47725 58638 47729 58694
rect 47785 58638 47789 58694
rect 47725 58624 47789 58638
rect 30015 58568 30026 58624
rect 30082 58568 30094 58624
rect 30015 58558 30094 58568
rect 30015 58544 30028 58558
rect 30080 58544 30094 58558
rect 30015 58488 30026 58544
rect 30082 58488 30094 58544
rect 30015 58464 30028 58488
rect 30080 58464 30094 58488
rect 30015 58408 30026 58464
rect 30082 58408 30094 58464
rect 30015 58384 30028 58408
rect 30080 58384 30094 58408
rect 30015 58328 30026 58384
rect 30082 58328 30094 58384
rect 30015 58314 30028 58328
rect 30080 58314 30094 58328
rect 30015 58304 30094 58314
rect 30015 58248 30026 58304
rect 30082 58248 30094 58304
rect 30015 58238 30094 58248
rect 30015 58224 30028 58238
rect 30080 58224 30094 58238
rect 30015 58168 30026 58224
rect 30082 58168 30094 58224
rect 30015 58144 30028 58168
rect 30080 58144 30094 58168
rect 60032 58205 60084 58726
rect 62524 58441 62588 58984
rect 62524 58389 62530 58441
rect 62582 58389 62588 58441
rect 62524 58373 62588 58389
rect 64336 59034 64400 59050
rect 64336 58982 64342 59034
rect 64394 58982 64400 59034
rect 64336 58441 64400 58982
rect 64336 58389 64342 58441
rect 64394 58389 64400 58441
rect 64336 58373 64400 58389
rect 63026 58213 63090 58227
rect 63026 58205 63030 58213
rect 60032 58157 63030 58205
rect 63086 58205 63090 58213
rect 66032 58205 66084 58812
rect 63086 58157 66084 58205
rect 60032 58153 66084 58157
rect 30015 58088 30026 58144
rect 30082 58088 30094 58144
rect 63026 58143 63090 58153
rect 30015 58064 30028 58088
rect 30080 58064 30094 58088
rect 30015 58008 30026 58064
rect 30082 58008 30094 58064
rect 30015 57994 30028 58008
rect 30080 57994 30094 58008
rect 30015 57984 30094 57994
rect 30015 57928 30026 57984
rect 30082 57928 30094 57984
rect 30015 57918 30094 57928
rect 30015 57904 30028 57918
rect 30080 57904 30094 57918
rect 30015 57848 30026 57904
rect 30082 57848 30094 57904
rect 30015 57824 30028 57848
rect 30080 57824 30094 57848
rect 30015 57768 30026 57824
rect 30082 57768 30094 57824
rect 60839 57872 60891 57882
rect 63832 57872 63896 57882
rect 66839 57872 66891 57882
rect 60891 57868 66839 57872
rect 60891 57820 63836 57868
rect 60839 57810 60891 57820
rect 63832 57812 63836 57820
rect 63892 57820 66839 57868
rect 66891 57820 66892 57872
rect 63892 57812 63896 57820
rect 63832 57798 63896 57812
rect 66839 57810 66891 57820
rect 30015 57744 30028 57768
rect 30080 57744 30094 57768
rect 30015 57688 30026 57744
rect 30082 57688 30094 57744
rect 30015 57674 30028 57688
rect 30080 57674 30094 57688
rect 30015 57664 30094 57674
rect 30015 57608 30026 57664
rect 30082 57608 30094 57664
rect 30015 57598 30094 57608
rect 30015 57584 30028 57598
rect 30080 57584 30094 57598
rect 30015 57528 30026 57584
rect 30082 57528 30094 57584
rect 30015 57510 30094 57528
rect 35576 57569 35640 57583
rect 35576 57513 35580 57569
rect 35636 57513 35640 57569
rect 35576 57499 35640 57513
rect 62524 57577 62588 57596
rect 62524 57525 62530 57577
rect 62582 57525 62588 57577
rect 50146 57197 50210 57211
rect 50146 57141 50150 57197
rect 50206 57141 50210 57197
rect 50146 57127 50210 57141
rect 30010 56904 30089 56931
rect 30010 56882 30023 56904
rect 30075 56882 30089 56904
rect 30010 56826 30021 56882
rect 30077 56826 30089 56882
rect 30010 56802 30023 56826
rect 30075 56802 30089 56826
rect 30010 56746 30021 56802
rect 30077 56746 30089 56802
rect 30010 56724 30023 56746
rect 30075 56724 30089 56746
rect 30010 56722 30089 56724
rect 30010 56666 30021 56722
rect 30077 56666 30089 56722
rect 30010 56660 30023 56666
rect 30075 56660 30089 56666
rect 30010 56648 30089 56660
rect 30010 56642 30023 56648
rect 30075 56642 30089 56648
rect 30010 56586 30021 56642
rect 30077 56586 30089 56642
rect 30010 56584 30089 56586
rect 30010 56562 30023 56584
rect 30075 56562 30089 56584
rect 30010 56506 30021 56562
rect 30077 56506 30089 56562
rect 30010 56482 30023 56506
rect 30075 56482 30089 56506
rect 30010 56426 30021 56482
rect 30077 56426 30089 56482
rect 30010 56404 30023 56426
rect 30075 56404 30089 56426
rect 30010 56377 30089 56404
rect 62411 56367 62475 56377
rect 62524 56367 62588 57525
rect 64522 57585 64586 57601
rect 64522 57533 64528 57585
rect 64580 57533 64586 57585
rect 64522 56384 64586 57533
rect 62411 56363 62588 56367
rect 62411 56307 62415 56363
rect 62471 56307 62588 56363
rect 62411 56303 62588 56307
rect 64458 56370 64586 56384
rect 64458 56314 64462 56370
rect 64518 56314 64586 56370
rect 64458 56310 64586 56314
rect 62411 56293 62475 56303
rect 64458 56300 64522 56310
rect 50105 55829 65151 55862
rect 50105 55827 65063 55829
rect 50105 55775 50111 55827
rect 50163 55775 50175 55827
rect 50227 55775 65063 55827
rect 50105 55773 65063 55775
rect 65119 55773 65151 55829
rect 50105 55734 65151 55773
rect 61448 54450 61512 54464
rect 61448 54394 61452 54450
rect 61508 54394 61512 54450
rect 61448 54380 61512 54394
rect 65422 54455 65486 54469
rect 65422 54399 65426 54455
rect 65482 54399 65486 54455
rect 65422 54385 65486 54399
rect 47747 54337 59547 54360
rect 47697 54327 59547 54337
rect 60420 54327 60484 54337
rect 47697 54323 60484 54327
rect 47697 54321 60424 54323
rect 47697 54269 47703 54321
rect 47755 54269 47767 54321
rect 47819 54269 60424 54321
rect 47697 54267 60424 54269
rect 60480 54267 60484 54323
rect 47697 54263 60484 54267
rect 47697 54253 59547 54263
rect 60420 54253 60484 54263
rect 47747 54232 59547 54253
rect 44401 53770 44465 53784
rect 44401 53714 44405 53770
rect 44461 53714 44465 53770
rect 44401 53700 44465 53714
rect 59007 53774 59071 53784
rect 73815 53774 73879 53784
rect 59007 53770 73879 53774
rect 59007 53714 59011 53770
rect 59067 53714 73819 53770
rect 73875 53714 73879 53770
rect 59007 53710 73879 53714
rect 59007 53700 59071 53710
rect 73815 53700 73879 53710
rect 43625 53347 43689 53361
rect 26895 53187 26901 53303
rect 27017 53187 27024 53303
rect 26895 53171 27024 53187
rect 38571 53303 38700 53320
rect 38571 53187 38577 53303
rect 38693 53187 38700 53303
rect 43625 53291 43629 53347
rect 43685 53291 43689 53347
rect 43625 53277 43689 53291
rect 59007 53351 59071 53361
rect 74506 53351 74570 53361
rect 59007 53347 74570 53351
rect 59007 53291 59011 53347
rect 59067 53291 74510 53347
rect 74566 53291 74570 53347
rect 59007 53287 74570 53291
rect 59007 53277 59071 53287
rect 74506 53277 74570 53287
rect 26064 51829 26070 51945
rect 26186 51829 26193 51945
rect 26064 51813 26193 51829
rect 37711 51945 37840 51962
rect 37711 51829 37717 51945
rect 37833 51829 37840 51945
rect 18904 50612 22238 50643
rect 18904 50610 18943 50612
rect 18999 50610 19023 50612
rect 19079 50610 19103 50612
rect 19159 50610 19183 50612
rect 19239 50610 19263 50612
rect 19319 50610 19343 50612
rect 19399 50610 19423 50612
rect 19479 50610 19503 50612
rect 19559 50610 19583 50612
rect 19639 50610 19663 50612
rect 19719 50610 19743 50612
rect 19799 50610 19823 50612
rect 19879 50610 19903 50612
rect 19959 50610 19983 50612
rect 20039 50610 20063 50612
rect 20119 50610 20143 50612
rect 20199 50610 20223 50612
rect 20279 50610 20303 50612
rect 20359 50610 20383 50612
rect 20439 50610 20463 50612
rect 20519 50610 20543 50612
rect 20599 50610 20623 50612
rect 20679 50610 20703 50612
rect 20759 50610 20783 50612
rect 20839 50610 20863 50612
rect 20919 50610 20943 50612
rect 20999 50610 21023 50612
rect 21079 50610 21103 50612
rect 21159 50610 21183 50612
rect 21239 50610 21263 50612
rect 21319 50610 21343 50612
rect 21399 50610 21423 50612
rect 21479 50610 21503 50612
rect 21559 50610 21583 50612
rect 21639 50610 21663 50612
rect 21719 50610 21743 50612
rect 21799 50610 21823 50612
rect 21879 50610 21903 50612
rect 21959 50610 21983 50612
rect 22039 50610 22063 50612
rect 22119 50610 22143 50612
rect 22199 50610 22238 50612
rect 18904 50558 18913 50610
rect 19093 50558 19103 50610
rect 19159 50558 19169 50610
rect 19413 50558 19423 50610
rect 19479 50558 19489 50610
rect 19733 50558 19743 50610
rect 19799 50558 19809 50610
rect 20053 50558 20063 50610
rect 20119 50558 20129 50610
rect 20373 50558 20383 50610
rect 20439 50558 20449 50610
rect 20693 50558 20703 50610
rect 20759 50558 20769 50610
rect 21013 50558 21023 50610
rect 21079 50558 21089 50610
rect 21333 50558 21343 50610
rect 21399 50558 21409 50610
rect 21653 50558 21663 50610
rect 21719 50558 21729 50610
rect 21973 50558 21983 50610
rect 22039 50558 22049 50610
rect 22229 50558 22238 50610
rect 18904 50556 18943 50558
rect 18999 50556 19023 50558
rect 19079 50556 19103 50558
rect 19159 50556 19183 50558
rect 19239 50556 19263 50558
rect 19319 50556 19343 50558
rect 19399 50556 19423 50558
rect 19479 50556 19503 50558
rect 19559 50556 19583 50558
rect 19639 50556 19663 50558
rect 19719 50556 19743 50558
rect 19799 50556 19823 50558
rect 19879 50556 19903 50558
rect 19959 50556 19983 50558
rect 20039 50556 20063 50558
rect 20119 50556 20143 50558
rect 20199 50556 20223 50558
rect 20279 50556 20303 50558
rect 20359 50556 20383 50558
rect 20439 50556 20463 50558
rect 20519 50556 20543 50558
rect 20599 50556 20623 50558
rect 20679 50556 20703 50558
rect 20759 50556 20783 50558
rect 20839 50556 20863 50558
rect 20919 50556 20943 50558
rect 20999 50556 21023 50558
rect 21079 50556 21103 50558
rect 21159 50556 21183 50558
rect 21239 50556 21263 50558
rect 21319 50556 21343 50558
rect 21399 50556 21423 50558
rect 21479 50556 21503 50558
rect 21559 50556 21583 50558
rect 21639 50556 21663 50558
rect 21719 50556 21743 50558
rect 21799 50556 21823 50558
rect 21879 50556 21903 50558
rect 21959 50556 21983 50558
rect 22039 50556 22063 50558
rect 22119 50556 22143 50558
rect 22199 50556 22238 50558
rect 18904 50526 22238 50556
rect 37711 50037 37840 51829
rect 38571 51631 38700 53187
rect 65054 52864 65118 52878
rect 59045 52830 59173 52840
rect 61795 52830 61859 52840
rect 59045 52826 61859 52830
rect 59045 52824 61799 52826
rect 59045 52772 59051 52824
rect 59103 52772 59115 52824
rect 59167 52772 61799 52824
rect 59045 52770 61799 52772
rect 61855 52770 61859 52826
rect 65054 52808 65058 52864
rect 65114 52808 65118 52864
rect 65054 52794 65118 52808
rect 59045 52766 61859 52770
rect 59045 52756 59173 52766
rect 61795 52756 61859 52766
rect 51008 52624 51136 52655
rect 51008 52572 51014 52624
rect 51066 52572 51078 52624
rect 51130 52572 51136 52624
rect 41382 52111 41481 52130
rect 41382 52081 41405 52111
rect 41457 52081 41481 52111
rect 41382 52025 41403 52081
rect 41459 52025 41481 52081
rect 41382 52001 41405 52025
rect 41457 52001 41481 52025
rect 41382 51945 41403 52001
rect 41459 51945 41481 52001
rect 41382 51931 41405 51945
rect 41457 51931 41481 51945
rect 41382 51921 41481 51931
rect 41382 51865 41403 51921
rect 41459 51865 41481 51921
rect 41382 51855 41481 51865
rect 41382 51841 41405 51855
rect 41457 51841 41481 51855
rect 41382 51785 41403 51841
rect 41459 51785 41481 51841
rect 41382 51761 41405 51785
rect 41457 51761 41481 51785
rect 41382 51705 41403 51761
rect 41459 51705 41481 51761
rect 39459 51660 39587 51676
rect 38571 51591 38848 51631
rect 38571 51539 38774 51591
rect 38826 51539 38848 51591
rect 38571 51502 38848 51539
rect 39459 51544 39465 51660
rect 39581 51544 39587 51660
rect 41382 51675 41405 51705
rect 41457 51675 41481 51705
rect 41382 51657 41481 51675
rect 43111 52088 43163 52098
rect 39459 51528 39587 51544
rect 42188 51593 42240 51603
rect 38768 51120 38832 51130
rect 38768 51114 39837 51120
rect 38768 51062 38774 51114
rect 38826 51062 39837 51114
rect 38768 51056 39837 51062
rect 42188 51105 42240 51541
rect 38768 51046 38832 51056
rect 38213 50782 38277 50792
rect 39838 50782 39902 50792
rect 38213 50776 39902 50782
rect 38213 50724 38219 50776
rect 38271 50724 39844 50776
rect 39896 50724 39902 50776
rect 38213 50718 39902 50724
rect 38213 50708 38277 50718
rect 39838 50708 39902 50718
rect 39459 50431 39587 50447
rect 39459 50315 39465 50431
rect 39581 50315 39587 50431
rect 39459 50299 39587 50315
rect 41369 50292 41458 50313
rect 41369 50236 41385 50292
rect 41441 50236 41458 50292
rect 41369 50222 41387 50236
rect 41439 50222 41458 50236
rect 41369 50212 41458 50222
rect 41369 50156 41385 50212
rect 41441 50156 41458 50212
rect 41369 50146 41458 50156
rect 41369 50132 41387 50146
rect 41439 50132 41458 50146
rect 41369 50076 41385 50132
rect 41441 50076 41458 50132
rect 41369 50056 41458 50076
rect 37711 49993 38278 50037
rect 37711 49941 38218 49993
rect 38270 49941 38278 49993
rect 37711 49908 38278 49941
rect 42188 49989 42240 51053
rect 42188 49927 42240 49937
rect 42690 51281 42742 51291
rect 42690 49681 42742 51229
rect 43111 50488 43163 52036
rect 44705 52083 44778 52108
rect 44705 52027 44713 52083
rect 44769 52027 44778 52083
rect 44705 52017 44778 52027
rect 44705 52003 44715 52017
rect 44767 52003 44778 52017
rect 44705 51947 44713 52003
rect 44769 51947 44778 52003
rect 44705 51923 44715 51947
rect 44767 51923 44778 51947
rect 44705 51867 44713 51923
rect 44769 51867 44778 51923
rect 44705 51843 44715 51867
rect 44767 51843 44778 51867
rect 44705 51787 44713 51843
rect 44769 51787 44778 51843
rect 44705 51773 44715 51787
rect 44767 51773 44778 51787
rect 44705 51763 44778 51773
rect 44705 51707 44713 51763
rect 44769 51707 44778 51763
rect 44705 51682 44778 51707
rect 44700 51442 44797 51459
rect 44700 51386 44720 51442
rect 44776 51386 44797 51442
rect 44700 51372 44722 51386
rect 44774 51372 44797 51386
rect 44700 51362 44797 51372
rect 44700 51306 44720 51362
rect 44776 51306 44797 51362
rect 44700 51296 44797 51306
rect 44700 51282 44722 51296
rect 44774 51282 44797 51296
rect 44700 51226 44720 51282
rect 44776 51226 44797 51282
rect 44700 51210 44797 51226
rect 47078 50604 47206 50620
rect 47078 50552 47084 50604
rect 47136 50552 47148 50604
rect 47200 50552 47206 50604
rect 43111 49696 43163 50436
rect 44698 50481 44793 50518
rect 44698 50425 44717 50481
rect 44773 50425 44793 50481
rect 44698 50415 44793 50425
rect 44698 50401 44719 50415
rect 44771 50401 44793 50415
rect 44698 50345 44717 50401
rect 44773 50345 44793 50401
rect 44698 50321 44719 50345
rect 44771 50321 44793 50345
rect 44698 50265 44717 50321
rect 44773 50265 44793 50321
rect 44698 50241 44719 50265
rect 44771 50241 44793 50265
rect 44698 50185 44717 50241
rect 44773 50185 44793 50241
rect 44698 50171 44719 50185
rect 44771 50171 44793 50185
rect 44698 50161 44793 50171
rect 44698 50105 44717 50161
rect 44773 50105 44793 50161
rect 44698 50069 44793 50105
rect 44710 49843 44773 49855
rect 44710 49787 44713 49843
rect 44769 49787 44773 49843
rect 44710 49773 44715 49787
rect 44767 49773 44773 49787
rect 44710 49763 44773 49773
rect 44710 49707 44713 49763
rect 44769 49707 44773 49763
rect 44710 49697 44773 49707
rect 31543 49549 32246 49601
rect 31645 49498 31725 49514
rect 31645 49442 31657 49498
rect 31713 49442 31725 49498
rect 31645 49420 31659 49442
rect 31711 49420 31725 49442
rect 31645 49418 31725 49420
rect 31645 49362 31657 49418
rect 31713 49362 31725 49418
rect 31645 49356 31659 49362
rect 31711 49356 31725 49362
rect 31645 49344 31725 49356
rect 31645 49338 31659 49344
rect 31711 49338 31725 49344
rect 31645 49282 31657 49338
rect 31713 49282 31725 49338
rect 31645 49280 31725 49282
rect 31645 49258 31659 49280
rect 31711 49258 31725 49280
rect 16501 49183 16737 49203
rect 31645 49202 31657 49258
rect 31713 49202 31725 49258
rect 31645 49187 31725 49202
rect 16501 48967 16511 49183
rect 16727 48967 16737 49183
rect 16501 48947 16737 48967
rect 24103 49128 24231 49144
rect 24103 49012 24109 49128
rect 24225 49012 24231 49128
rect 18912 47604 22242 47637
rect 18912 47602 18949 47604
rect 19005 47602 19029 47604
rect 19085 47602 19109 47604
rect 19165 47602 19189 47604
rect 19245 47602 19269 47604
rect 19325 47602 19349 47604
rect 19405 47602 19429 47604
rect 19485 47602 19509 47604
rect 19565 47602 19589 47604
rect 19645 47602 19669 47604
rect 19725 47602 19749 47604
rect 19805 47602 19829 47604
rect 19885 47602 19909 47604
rect 19965 47602 19989 47604
rect 20045 47602 20069 47604
rect 20125 47602 20149 47604
rect 20205 47602 20229 47604
rect 20285 47602 20309 47604
rect 20365 47602 20389 47604
rect 20445 47602 20469 47604
rect 20525 47602 20549 47604
rect 20605 47602 20629 47604
rect 20685 47602 20709 47604
rect 20765 47602 20789 47604
rect 20845 47602 20869 47604
rect 20925 47602 20949 47604
rect 21005 47602 21029 47604
rect 21085 47602 21109 47604
rect 21165 47602 21189 47604
rect 21245 47602 21269 47604
rect 21325 47602 21349 47604
rect 21405 47602 21429 47604
rect 21485 47602 21509 47604
rect 21565 47602 21589 47604
rect 21645 47602 21669 47604
rect 21725 47602 21749 47604
rect 21805 47602 21829 47604
rect 21885 47602 21909 47604
rect 21965 47602 21989 47604
rect 22045 47602 22069 47604
rect 22125 47602 22149 47604
rect 22205 47602 22242 47604
rect 18912 47550 18919 47602
rect 19099 47550 19109 47602
rect 19165 47550 19175 47602
rect 19419 47550 19429 47602
rect 19485 47550 19495 47602
rect 19739 47550 19749 47602
rect 19805 47550 19815 47602
rect 20059 47550 20069 47602
rect 20125 47550 20135 47602
rect 20379 47550 20389 47602
rect 20445 47550 20455 47602
rect 20699 47550 20709 47602
rect 20765 47550 20775 47602
rect 21019 47550 21029 47602
rect 21085 47550 21095 47602
rect 21339 47550 21349 47602
rect 21405 47550 21415 47602
rect 21659 47550 21669 47602
rect 21725 47550 21735 47602
rect 21979 47550 21989 47602
rect 22045 47550 22055 47602
rect 22235 47550 22242 47602
rect 18912 47548 18949 47550
rect 19005 47548 19029 47550
rect 19085 47548 19109 47550
rect 19165 47548 19189 47550
rect 19245 47548 19269 47550
rect 19325 47548 19349 47550
rect 19405 47548 19429 47550
rect 19485 47548 19509 47550
rect 19565 47548 19589 47550
rect 19645 47548 19669 47550
rect 19725 47548 19749 47550
rect 19805 47548 19829 47550
rect 19885 47548 19909 47550
rect 19965 47548 19989 47550
rect 20045 47548 20069 47550
rect 20125 47548 20149 47550
rect 20205 47548 20229 47550
rect 20285 47548 20309 47550
rect 20365 47548 20389 47550
rect 20445 47548 20469 47550
rect 20525 47548 20549 47550
rect 20605 47548 20629 47550
rect 20685 47548 20709 47550
rect 20765 47548 20789 47550
rect 20845 47548 20869 47550
rect 20925 47548 20949 47550
rect 21005 47548 21029 47550
rect 21085 47548 21109 47550
rect 21165 47548 21189 47550
rect 21245 47548 21269 47550
rect 21325 47548 21349 47550
rect 21405 47548 21429 47550
rect 21485 47548 21509 47550
rect 21565 47548 21589 47550
rect 21645 47548 21669 47550
rect 21725 47548 21749 47550
rect 21805 47548 21829 47550
rect 21885 47548 21909 47550
rect 21965 47548 21989 47550
rect 22045 47548 22069 47550
rect 22125 47548 22149 47550
rect 22205 47548 22242 47550
rect 18912 47515 22242 47548
rect 18926 43076 22233 43097
rect 18926 43020 18951 43076
rect 19007 43074 19031 43076
rect 19087 43074 19111 43076
rect 19167 43074 19191 43076
rect 19247 43074 19271 43076
rect 19327 43074 19351 43076
rect 19407 43074 19431 43076
rect 19487 43074 19511 43076
rect 19567 43074 19591 43076
rect 19647 43074 19671 43076
rect 19727 43074 19751 43076
rect 19807 43074 19831 43076
rect 19887 43074 19911 43076
rect 19967 43074 19991 43076
rect 20047 43074 20071 43076
rect 20127 43074 20151 43076
rect 20207 43074 20231 43076
rect 20287 43074 20311 43076
rect 20367 43074 20391 43076
rect 20447 43074 20471 43076
rect 20527 43074 20551 43076
rect 20607 43074 20631 43076
rect 20687 43074 20711 43076
rect 20767 43074 20791 43076
rect 20847 43074 20871 43076
rect 20927 43074 20951 43076
rect 21007 43074 21031 43076
rect 21087 43074 21111 43076
rect 21167 43074 21191 43076
rect 21247 43074 21271 43076
rect 21327 43074 21351 43076
rect 21407 43074 21431 43076
rect 21487 43074 21511 43076
rect 21567 43074 21591 43076
rect 21647 43074 21671 43076
rect 21727 43074 21751 43076
rect 21807 43074 21831 43076
rect 21887 43074 21911 43076
rect 21967 43074 21991 43076
rect 22047 43074 22071 43076
rect 22127 43074 22151 43076
rect 19007 43022 19017 43074
rect 19261 43022 19271 43074
rect 19327 43022 19337 43074
rect 19581 43022 19591 43074
rect 19647 43022 19657 43074
rect 19901 43022 19911 43074
rect 19967 43022 19977 43074
rect 20221 43022 20231 43074
rect 20287 43022 20297 43074
rect 20541 43022 20551 43074
rect 20607 43022 20617 43074
rect 20861 43022 20871 43074
rect 20927 43022 20937 43074
rect 21181 43022 21191 43074
rect 21247 43022 21257 43074
rect 21501 43022 21511 43074
rect 21567 43022 21577 43074
rect 21821 43022 21831 43074
rect 21887 43022 21897 43074
rect 22141 43022 22151 43074
rect 19007 43020 19031 43022
rect 19087 43020 19111 43022
rect 19167 43020 19191 43022
rect 19247 43020 19271 43022
rect 19327 43020 19351 43022
rect 19407 43020 19431 43022
rect 19487 43020 19511 43022
rect 19567 43020 19591 43022
rect 19647 43020 19671 43022
rect 19727 43020 19751 43022
rect 19807 43020 19831 43022
rect 19887 43020 19911 43022
rect 19967 43020 19991 43022
rect 20047 43020 20071 43022
rect 20127 43020 20151 43022
rect 20207 43020 20231 43022
rect 20287 43020 20311 43022
rect 20367 43020 20391 43022
rect 20447 43020 20471 43022
rect 20527 43020 20551 43022
rect 20607 43020 20631 43022
rect 20687 43020 20711 43022
rect 20767 43020 20791 43022
rect 20847 43020 20871 43022
rect 20927 43020 20951 43022
rect 21007 43020 21031 43022
rect 21087 43020 21111 43022
rect 21167 43020 21191 43022
rect 21247 43020 21271 43022
rect 21327 43020 21351 43022
rect 21407 43020 21431 43022
rect 21487 43020 21511 43022
rect 21567 43020 21591 43022
rect 21647 43020 21671 43022
rect 21727 43020 21751 43022
rect 21807 43020 21831 43022
rect 21887 43020 21911 43022
rect 21967 43020 21991 43022
rect 22047 43020 22071 43022
rect 22127 43020 22151 43022
rect 22207 43020 22233 43076
rect 18926 42999 22233 43020
rect 16498 41642 16734 41662
rect 16498 41426 16508 41642
rect 16724 41426 16734 41642
rect 16498 41406 16734 41426
rect 18920 40081 22242 40107
rect 18920 40079 18953 40081
rect 19009 40079 19033 40081
rect 19089 40079 19113 40081
rect 19169 40079 19193 40081
rect 19249 40079 19273 40081
rect 19329 40079 19353 40081
rect 19409 40079 19433 40081
rect 19489 40079 19513 40081
rect 19569 40079 19593 40081
rect 19649 40079 19673 40081
rect 19729 40079 19753 40081
rect 19809 40079 19833 40081
rect 19889 40079 19913 40081
rect 19969 40079 19993 40081
rect 20049 40079 20073 40081
rect 20129 40079 20153 40081
rect 20209 40079 20233 40081
rect 20289 40079 20313 40081
rect 20369 40079 20393 40081
rect 20449 40079 20473 40081
rect 20529 40079 20553 40081
rect 20609 40079 20633 40081
rect 20689 40079 20713 40081
rect 20769 40079 20793 40081
rect 20849 40079 20873 40081
rect 20929 40079 20953 40081
rect 21009 40079 21033 40081
rect 21089 40079 21113 40081
rect 21169 40079 21193 40081
rect 21249 40079 21273 40081
rect 21329 40079 21353 40081
rect 21409 40079 21433 40081
rect 21489 40079 21513 40081
rect 21569 40079 21593 40081
rect 21649 40079 21673 40081
rect 21729 40079 21753 40081
rect 21809 40079 21833 40081
rect 21889 40079 21913 40081
rect 21969 40079 21993 40081
rect 22049 40079 22073 40081
rect 22129 40079 22153 40081
rect 22209 40079 22242 40081
rect 18920 40027 18923 40079
rect 19103 40027 19113 40079
rect 19169 40027 19179 40079
rect 19423 40027 19433 40079
rect 19489 40027 19499 40079
rect 19743 40027 19753 40079
rect 19809 40027 19819 40079
rect 20063 40027 20073 40079
rect 20129 40027 20139 40079
rect 20383 40027 20393 40079
rect 20449 40027 20459 40079
rect 20703 40027 20713 40079
rect 20769 40027 20779 40079
rect 21023 40027 21033 40079
rect 21089 40027 21099 40079
rect 21343 40027 21353 40079
rect 21409 40027 21419 40079
rect 21663 40027 21673 40079
rect 21729 40027 21739 40079
rect 21983 40027 21993 40079
rect 22049 40027 22059 40079
rect 22239 40027 22242 40079
rect 18920 40025 18953 40027
rect 19009 40025 19033 40027
rect 19089 40025 19113 40027
rect 19169 40025 19193 40027
rect 19249 40025 19273 40027
rect 19329 40025 19353 40027
rect 19409 40025 19433 40027
rect 19489 40025 19513 40027
rect 19569 40025 19593 40027
rect 19649 40025 19673 40027
rect 19729 40025 19753 40027
rect 19809 40025 19833 40027
rect 19889 40025 19913 40027
rect 19969 40025 19993 40027
rect 20049 40025 20073 40027
rect 20129 40025 20153 40027
rect 20209 40025 20233 40027
rect 20289 40025 20313 40027
rect 20369 40025 20393 40027
rect 20449 40025 20473 40027
rect 20529 40025 20553 40027
rect 20609 40025 20633 40027
rect 20689 40025 20713 40027
rect 20769 40025 20793 40027
rect 20849 40025 20873 40027
rect 20929 40025 20953 40027
rect 21009 40025 21033 40027
rect 21089 40025 21113 40027
rect 21169 40025 21193 40027
rect 21249 40025 21273 40027
rect 21329 40025 21353 40027
rect 21409 40025 21433 40027
rect 21489 40025 21513 40027
rect 21569 40025 21593 40027
rect 21649 40025 21673 40027
rect 21729 40025 21753 40027
rect 21809 40025 21833 40027
rect 21889 40025 21913 40027
rect 21969 40025 21993 40027
rect 22049 40025 22073 40027
rect 22129 40025 22153 40027
rect 22209 40025 22242 40027
rect 18920 39999 22242 40025
rect 24103 38118 24231 49012
rect 31642 48959 31729 48977
rect 31642 48903 31657 48959
rect 31713 48903 31729 48959
rect 31642 48889 31659 48903
rect 31711 48889 31729 48903
rect 31642 48879 31729 48889
rect 31642 48823 31657 48879
rect 31713 48823 31729 48879
rect 31642 48813 31729 48823
rect 31642 48799 31659 48813
rect 31711 48799 31729 48813
rect 29916 48741 30418 48793
rect 31642 48743 31657 48799
rect 31713 48743 31729 48799
rect 29916 45022 29968 48741
rect 31642 48726 31729 48743
rect 29155 44970 29968 45022
rect 24103 38002 24109 38118
rect 24225 38002 24231 38118
rect 24103 37986 24231 38002
rect 25964 41598 26092 41614
rect 25964 41482 25970 41598
rect 26086 41482 26092 41598
rect 25964 30353 26092 41482
rect 29155 39473 29207 44970
rect 29916 41251 29968 44970
rect 32194 45830 32246 49549
rect 41367 49442 41462 49479
rect 41367 49386 41386 49442
rect 41442 49386 41462 49442
rect 41367 49376 41462 49386
rect 41367 49362 41388 49376
rect 41440 49362 41462 49376
rect 41367 49306 41386 49362
rect 41442 49306 41462 49362
rect 41367 49282 41388 49306
rect 41440 49282 41462 49306
rect 41367 49226 41386 49282
rect 41442 49226 41462 49282
rect 41367 49202 41388 49226
rect 41440 49202 41462 49226
rect 41367 49146 41386 49202
rect 41442 49146 41462 49202
rect 41367 49132 41388 49146
rect 41440 49132 41462 49146
rect 41367 49122 41462 49132
rect 41367 49066 41386 49122
rect 41442 49066 41462 49122
rect 39459 49018 39587 49034
rect 41367 49030 41462 49066
rect 39459 48902 39465 49018
rect 39581 48902 39587 49018
rect 42690 48904 42742 49629
rect 43105 49682 43169 49696
rect 43105 49626 43109 49682
rect 43165 49626 43169 49682
rect 43105 49612 43169 49626
rect 44710 49683 44715 49697
rect 44767 49683 44773 49697
rect 44710 49627 44713 49683
rect 44769 49627 44773 49683
rect 44710 49616 44773 49627
rect 39459 48886 39587 48902
rect 42684 48890 42748 48904
rect 42684 48834 42688 48890
rect 42744 48834 42748 48890
rect 42684 48820 42748 48834
rect 43111 48888 43163 49612
rect 38768 48480 38832 48489
rect 38768 48473 39823 48480
rect 38768 48421 38774 48473
rect 38826 48421 39823 48473
rect 38768 48416 39823 48421
rect 42186 48463 42238 48473
rect 38768 48405 38832 48416
rect 38213 48140 38277 48150
rect 39831 48140 39895 48150
rect 38213 48134 39895 48140
rect 38213 48082 38219 48134
rect 38271 48082 39837 48134
rect 39889 48082 39895 48134
rect 38213 48076 39895 48082
rect 38213 48066 38277 48076
rect 39831 48066 39895 48076
rect 39459 47789 39587 47805
rect 39459 47673 39465 47789
rect 39581 47673 39587 47789
rect 39459 47657 39587 47673
rect 41369 47651 41436 47669
rect 41369 47595 41374 47651
rect 41430 47595 41436 47651
rect 41369 47581 41376 47595
rect 41428 47581 41436 47595
rect 41369 47571 41436 47581
rect 41369 47515 41374 47571
rect 41430 47515 41436 47571
rect 41369 47505 41436 47515
rect 41369 47491 41376 47505
rect 41428 47491 41436 47505
rect 41369 47435 41374 47491
rect 41430 47435 41436 47491
rect 41369 47417 41436 47435
rect 42186 46793 42238 48411
rect 42186 46735 42238 46741
rect 42690 48081 42742 48820
rect 42690 46481 42742 48029
rect 43111 47288 43163 48836
rect 44701 48729 44766 48744
rect 44701 48715 44707 48729
rect 44759 48715 44766 48729
rect 44701 48659 44705 48715
rect 44761 48659 44766 48715
rect 44701 48635 44707 48659
rect 44759 48635 44766 48659
rect 44701 48579 44705 48635
rect 44761 48579 44766 48635
rect 44701 48555 44707 48579
rect 44759 48555 44766 48579
rect 44701 48499 44705 48555
rect 44761 48499 44766 48555
rect 44701 48485 44707 48499
rect 44759 48485 44766 48499
rect 44701 48470 44766 48485
rect 44696 48251 44778 48271
rect 44696 48195 44709 48251
rect 44765 48195 44778 48251
rect 44696 48181 44711 48195
rect 44763 48181 44778 48195
rect 44696 48171 44778 48181
rect 44696 48115 44709 48171
rect 44765 48115 44778 48171
rect 44696 48105 44778 48115
rect 44696 48091 44711 48105
rect 44763 48091 44778 48105
rect 44696 48035 44709 48091
rect 44765 48035 44778 48091
rect 44696 48015 44778 48035
rect 43111 47225 43163 47236
rect 44705 47277 44775 47309
rect 44705 47221 44712 47277
rect 44768 47221 44775 47277
rect 44705 47211 44775 47221
rect 44705 47197 44714 47211
rect 44766 47197 44775 47211
rect 44705 47141 44712 47197
rect 44768 47141 44775 47197
rect 44705 47117 44714 47141
rect 44766 47117 44775 47141
rect 44705 47061 44712 47117
rect 44768 47061 44775 47117
rect 44705 47037 44714 47061
rect 44766 47037 44775 47061
rect 44705 46981 44712 47037
rect 44768 46981 44775 47037
rect 44705 46967 44714 46981
rect 44766 46967 44775 46981
rect 44705 46957 44775 46967
rect 44705 46901 44712 46957
rect 44768 46901 44775 46957
rect 44705 46869 44775 46901
rect 45493 46792 45621 46808
rect 45493 46740 45499 46792
rect 45551 46740 45563 46792
rect 45615 46740 45621 46792
rect 42690 46419 42742 46429
rect 44703 46641 44771 46656
rect 44703 46585 44709 46641
rect 44765 46585 44771 46641
rect 44703 46571 44711 46585
rect 44763 46571 44771 46585
rect 44703 46561 44771 46571
rect 44703 46505 44709 46561
rect 44765 46505 44771 46561
rect 44703 46495 44771 46505
rect 44703 46481 44711 46495
rect 44763 46481 44771 46495
rect 44703 46425 44709 46481
rect 44765 46425 44771 46481
rect 44703 46411 44771 46425
rect 45493 45873 45621 46740
rect 32194 45778 33007 45830
rect 32194 42060 32246 45778
rect 31537 42008 32246 42060
rect 31642 41918 31707 41954
rect 31642 41904 31648 41918
rect 31700 41904 31707 41918
rect 31642 41848 31646 41904
rect 31702 41848 31707 41904
rect 31642 41824 31648 41848
rect 31700 41824 31707 41848
rect 31642 41768 31646 41824
rect 31702 41768 31707 41824
rect 31642 41744 31648 41768
rect 31700 41744 31707 41768
rect 31642 41688 31646 41744
rect 31702 41688 31707 41744
rect 31642 41674 31648 41688
rect 31700 41674 31707 41688
rect 31642 41639 31707 41674
rect 31644 41416 31716 41436
rect 31644 41360 31652 41416
rect 31708 41360 31716 41416
rect 31644 41346 31654 41360
rect 31706 41346 31716 41360
rect 31644 41336 31716 41346
rect 31644 41280 31652 41336
rect 31708 41280 31716 41336
rect 31644 41270 31716 41280
rect 31644 41256 31654 41270
rect 31706 41256 31716 41270
rect 29916 41199 30342 41251
rect 31644 41200 31652 41256
rect 31708 41200 31716 41256
rect 31644 41181 31716 41200
rect 32955 40281 33007 45778
rect 32903 40267 33007 40281
rect 32903 40211 32928 40267
rect 32984 40211 33007 40267
rect 32903 40197 33007 40211
rect 29155 39459 29259 39473
rect 29155 39403 29178 39459
rect 29234 39403 29259 39459
rect 29155 39389 29259 39403
rect 29155 33893 29207 39389
rect 31522 38536 32178 38584
rect 31519 38535 32178 38536
rect 31522 38532 32178 38535
rect 31577 38445 31650 38478
rect 31577 38431 31587 38445
rect 31639 38431 31650 38445
rect 31577 38375 31585 38431
rect 31641 38375 31650 38431
rect 31577 38351 31587 38375
rect 31639 38351 31650 38375
rect 31577 38295 31585 38351
rect 31641 38295 31650 38351
rect 31577 38271 31587 38295
rect 31639 38271 31650 38295
rect 31577 38215 31585 38271
rect 31641 38215 31650 38271
rect 31577 38201 31587 38215
rect 31639 38201 31650 38215
rect 31577 38169 31650 38201
rect 31576 37937 31648 37957
rect 31576 37881 31584 37937
rect 31640 37881 31648 37937
rect 31576 37867 31586 37881
rect 31638 37867 31648 37881
rect 31576 37857 31648 37867
rect 31576 37801 31584 37857
rect 31640 37801 31648 37857
rect 31576 37791 31648 37801
rect 31576 37777 31586 37791
rect 31638 37777 31648 37791
rect 29848 37745 30279 37777
rect 29848 37736 30282 37745
rect 29848 37725 30279 37736
rect 29848 33893 29900 37725
rect 31576 37721 31584 37777
rect 31640 37721 31648 37777
rect 31576 37702 31648 37721
rect 29155 33841 29900 33893
rect 25964 30237 25970 30353
rect 26086 30237 26092 30353
rect 25964 30221 26092 30237
rect 29848 30009 29900 33841
rect 32126 34699 32178 38532
rect 32955 34699 33007 40197
rect 40313 45745 45621 45873
rect 38871 38091 38935 38105
rect 38871 38035 38875 38091
rect 38931 38035 38935 38091
rect 38871 38021 38935 38035
rect 32126 34647 33007 34699
rect 32126 30815 32178 34647
rect 40313 31625 40441 45745
rect 47078 45098 47206 50552
rect 51008 45687 51136 52572
rect 60493 52617 60557 52627
rect 61422 52617 61486 52627
rect 60493 52613 61492 52617
rect 60493 52611 61426 52613
rect 60493 52559 60499 52611
rect 60551 52559 61426 52611
rect 60493 52557 61426 52559
rect 61482 52557 61492 52613
rect 60493 52553 61492 52557
rect 65432 52614 65496 52624
rect 66493 52614 66557 52624
rect 65432 52610 66567 52614
rect 65432 52554 65436 52610
rect 65492 52608 66567 52610
rect 65492 52556 66499 52608
rect 66551 52556 66567 52608
rect 65492 52554 66567 52556
rect 60493 52543 60557 52553
rect 61422 52543 61486 52553
rect 65432 52550 66567 52554
rect 65432 52540 65496 52550
rect 66493 52540 66557 52550
rect 51815 51554 51879 51564
rect 51815 51550 77029 51554
rect 51815 51494 51819 51550
rect 51875 51494 77029 51550
rect 51815 51490 77029 51494
rect 51815 51480 51879 51490
rect 53176 50877 53240 50887
rect 53176 50873 74671 50877
rect 53176 50817 53180 50873
rect 53236 50817 74671 50873
rect 53176 50813 74671 50817
rect 53176 50803 53240 50813
rect 59046 49842 59174 49852
rect 65054 49842 65118 49852
rect 59046 49836 65118 49842
rect 59046 49784 59052 49836
rect 59104 49784 59116 49836
rect 59168 49784 65060 49836
rect 65112 49784 65118 49836
rect 59046 49778 65118 49784
rect 59046 49768 59174 49778
rect 65054 49768 65118 49778
rect 51008 45635 51014 45687
rect 51066 45635 51078 45687
rect 51130 45635 51136 45687
rect 51008 45619 51136 45635
rect 53593 49430 53721 49455
rect 53593 49378 53599 49430
rect 53651 49378 53663 49430
rect 53715 49378 53721 49430
rect 42910 44970 47206 45098
rect 42910 39388 43038 44970
rect 53593 44825 53721 49378
rect 74607 48824 74671 50813
rect 76965 50027 77029 51490
rect 76965 49971 76969 50027
rect 77025 49971 77029 50027
rect 76965 49957 77029 49971
rect 76967 49616 77031 49630
rect 76967 49560 76971 49616
rect 77027 49560 77031 49616
rect 76967 48824 77031 49560
rect 74607 48760 77031 48824
rect 62809 48600 62877 48626
rect 62809 48544 62815 48600
rect 62871 48544 62877 48600
rect 62809 48534 62877 48544
rect 64162 48610 64226 48624
rect 64162 48554 64166 48610
rect 64222 48554 64226 48610
rect 64162 48540 64226 48554
rect 62809 48520 62817 48534
rect 62869 48520 62877 48534
rect 62809 48464 62815 48520
rect 62871 48464 62877 48520
rect 62809 48440 62817 48464
rect 62869 48440 62877 48464
rect 62809 48384 62815 48440
rect 62871 48384 62877 48440
rect 62809 48360 62817 48384
rect 62869 48360 62877 48384
rect 62809 48304 62815 48360
rect 62871 48304 62877 48360
rect 62809 48290 62817 48304
rect 62869 48290 62877 48304
rect 62809 48280 62877 48290
rect 62809 48224 62815 48280
rect 62871 48224 62877 48280
rect 62809 48198 62877 48224
rect 99950 48169 103284 48206
rect 99950 48167 99989 48169
rect 100045 48167 100069 48169
rect 100125 48167 100149 48169
rect 100205 48167 100229 48169
rect 100285 48167 100309 48169
rect 100365 48167 100389 48169
rect 100445 48167 100469 48169
rect 100525 48167 100549 48169
rect 100605 48167 100629 48169
rect 100685 48167 100709 48169
rect 100765 48167 100789 48169
rect 100845 48167 100869 48169
rect 100925 48167 100949 48169
rect 101005 48167 101029 48169
rect 101085 48167 101109 48169
rect 101165 48167 101189 48169
rect 101245 48167 101269 48169
rect 101325 48167 101349 48169
rect 101405 48167 101429 48169
rect 101485 48167 101509 48169
rect 101565 48167 101589 48169
rect 101645 48167 101669 48169
rect 101725 48167 101749 48169
rect 101805 48167 101829 48169
rect 101885 48167 101909 48169
rect 101965 48167 101989 48169
rect 102045 48167 102069 48169
rect 102125 48167 102149 48169
rect 102205 48167 102229 48169
rect 102285 48167 102309 48169
rect 102365 48167 102389 48169
rect 102445 48167 102469 48169
rect 102525 48167 102549 48169
rect 102605 48167 102629 48169
rect 102685 48167 102709 48169
rect 102765 48167 102789 48169
rect 102845 48167 102869 48169
rect 102925 48167 102949 48169
rect 103005 48167 103029 48169
rect 103085 48167 103109 48169
rect 103165 48167 103189 48169
rect 103245 48167 103284 48169
rect 60493 48119 60557 48131
rect 62737 48119 62801 48129
rect 60493 48117 62801 48119
rect 60493 48065 60499 48117
rect 60551 48113 62801 48117
rect 60551 48065 62743 48113
rect 60493 48061 62743 48065
rect 62795 48061 62801 48113
rect 60493 48055 62801 48061
rect 60493 48049 60557 48055
rect 62737 48045 62801 48055
rect 64111 48123 64175 48133
rect 66493 48123 66557 48133
rect 64111 48117 66561 48123
rect 64111 48065 64117 48117
rect 64169 48065 66499 48117
rect 66551 48065 66561 48117
rect 99950 48115 99959 48167
rect 100139 48115 100149 48167
rect 100205 48115 100215 48167
rect 100459 48115 100469 48167
rect 100525 48115 100535 48167
rect 100779 48115 100789 48167
rect 100845 48115 100855 48167
rect 101099 48115 101109 48167
rect 101165 48115 101175 48167
rect 101419 48115 101429 48167
rect 101485 48115 101495 48167
rect 101739 48115 101749 48167
rect 101805 48115 101815 48167
rect 102059 48115 102069 48167
rect 102125 48115 102135 48167
rect 102379 48115 102389 48167
rect 102445 48115 102455 48167
rect 102699 48115 102709 48167
rect 102765 48115 102775 48167
rect 103019 48115 103029 48167
rect 103085 48115 103095 48167
rect 103275 48115 103284 48167
rect 99950 48113 99989 48115
rect 100045 48113 100069 48115
rect 100125 48113 100149 48115
rect 100205 48113 100229 48115
rect 100285 48113 100309 48115
rect 100365 48113 100389 48115
rect 100445 48113 100469 48115
rect 100525 48113 100549 48115
rect 100605 48113 100629 48115
rect 100685 48113 100709 48115
rect 100765 48113 100789 48115
rect 100845 48113 100869 48115
rect 100925 48113 100949 48115
rect 101005 48113 101029 48115
rect 101085 48113 101109 48115
rect 101165 48113 101189 48115
rect 101245 48113 101269 48115
rect 101325 48113 101349 48115
rect 101405 48113 101429 48115
rect 101485 48113 101509 48115
rect 101565 48113 101589 48115
rect 101645 48113 101669 48115
rect 101725 48113 101749 48115
rect 101805 48113 101829 48115
rect 101885 48113 101909 48115
rect 101965 48113 101989 48115
rect 102045 48113 102069 48115
rect 102125 48113 102149 48115
rect 102205 48113 102229 48115
rect 102285 48113 102309 48115
rect 102365 48113 102389 48115
rect 102445 48113 102469 48115
rect 102525 48113 102549 48115
rect 102605 48113 102629 48115
rect 102685 48113 102709 48115
rect 102765 48113 102789 48115
rect 102845 48113 102869 48115
rect 102925 48113 102949 48115
rect 103005 48113 103029 48115
rect 103085 48113 103109 48115
rect 103165 48113 103189 48115
rect 103245 48113 103284 48115
rect 99950 48077 103284 48113
rect 64111 48059 66561 48065
rect 64111 48049 64175 48059
rect 66493 48049 66557 48059
rect 93160 48036 93224 48050
rect 93160 48034 93164 48036
rect 93033 47982 93164 48034
rect 93160 47980 93164 47982
rect 93220 47980 93224 48036
rect 93160 47966 93224 47980
rect 92246 47884 92310 47898
rect 92246 47828 92250 47884
rect 92306 47828 92310 47884
rect 92246 47814 92310 47828
rect 64185 47670 64249 47804
rect 64185 47614 64189 47670
rect 64245 47614 64249 47670
rect 96440 47733 96514 47746
rect 96440 47677 96449 47733
rect 96505 47677 96514 47733
rect 96440 47663 96451 47677
rect 96503 47663 96514 47677
rect 96440 47653 96514 47663
rect 64185 47600 64249 47614
rect 94913 47631 94986 47643
rect 94913 47601 94923 47631
rect 94975 47601 94986 47631
rect 94913 47545 94921 47601
rect 94977 47545 94986 47601
rect 94913 47515 94923 47545
rect 94975 47515 94986 47545
rect 94913 47504 94986 47515
rect 96440 47597 96449 47653
rect 96505 47597 96514 47653
rect 96440 47587 96514 47597
rect 96440 47573 96451 47587
rect 96503 47573 96514 47587
rect 96440 47517 96449 47573
rect 96505 47517 96514 47573
rect 96440 47505 96514 47517
rect 65881 47351 66037 47388
rect 65881 47295 65891 47351
rect 65947 47349 65971 47351
rect 65953 47297 65965 47349
rect 65947 47295 65971 47297
rect 66027 47295 66037 47351
rect 65881 47258 66037 47295
rect 94913 47214 94999 47226
rect 94913 47200 94930 47214
rect 94982 47200 94999 47214
rect 94913 47144 94928 47200
rect 94984 47144 94999 47200
rect 94913 47120 94930 47144
rect 94982 47120 94999 47144
rect 59644 47081 59708 47095
rect 59644 47025 59648 47081
rect 59704 47025 59708 47081
rect 59644 47011 59708 47025
rect 67296 47081 67360 47095
rect 67296 47025 67300 47081
rect 67356 47025 67360 47081
rect 67296 47011 67360 47025
rect 94913 47064 94928 47120
rect 94984 47064 94999 47120
rect 94913 47040 94930 47064
rect 94982 47040 94999 47064
rect 94913 46984 94928 47040
rect 94984 46984 94999 47040
rect 94913 46970 94930 46984
rect 94982 46970 94999 46984
rect 94913 46958 94999 46970
rect 96429 47220 96515 47232
rect 96429 47206 96446 47220
rect 96498 47206 96515 47220
rect 96429 47150 96444 47206
rect 96500 47150 96515 47206
rect 96429 47126 96446 47150
rect 96498 47126 96515 47150
rect 96429 47070 96444 47126
rect 96500 47070 96515 47126
rect 96429 47046 96446 47070
rect 96498 47046 96515 47070
rect 96429 46990 96444 47046
rect 96500 46990 96515 47046
rect 96429 46976 96446 46990
rect 96498 46976 96515 46990
rect 96429 46964 96515 46976
rect 92194 46812 92374 46822
rect 92854 46749 93115 46762
rect 92854 46747 92876 46749
rect 92932 46747 92956 46749
rect 93012 46747 93036 46749
rect 93092 46747 93115 46749
rect 92854 46695 92862 46747
rect 93106 46695 93115 46747
rect 92854 46693 92876 46695
rect 92932 46693 92956 46695
rect 93012 46693 93036 46695
rect 93092 46693 93115 46695
rect 92854 46680 93115 46693
rect 104650 46746 104886 46766
rect 92194 46622 92374 46632
rect 104650 46530 104660 46746
rect 104876 46530 104886 46746
rect 104650 46510 104886 46530
rect 96440 46407 96514 46420
rect 96440 46351 96449 46407
rect 96505 46351 96514 46407
rect 96440 46337 96451 46351
rect 96503 46337 96514 46351
rect 96440 46327 96514 46337
rect 94920 46295 94990 46312
rect 94920 46265 94929 46295
rect 94981 46265 94990 46295
rect 94920 46209 94927 46265
rect 94983 46209 94990 46265
rect 94920 46179 94929 46209
rect 94981 46179 94990 46209
rect 96440 46271 96449 46327
rect 96505 46271 96514 46327
rect 96440 46261 96514 46271
rect 96440 46247 96451 46261
rect 96503 46247 96514 46261
rect 96440 46191 96449 46247
rect 96505 46191 96514 46247
rect 96440 46179 96514 46191
rect 94920 46163 94990 46179
rect 61491 46059 61543 46069
rect 53593 44773 53599 44825
rect 53651 44773 53663 44825
rect 53715 44773 53721 44825
rect 53593 44757 53721 44773
rect 56123 45643 56187 45657
rect 56123 45587 56127 45643
rect 56183 45587 56187 45643
rect 56123 44733 56187 45587
rect 60004 45634 60056 46036
rect 60873 46007 61491 46059
rect 61491 45997 61543 46007
rect 65322 46059 65374 46069
rect 65374 46007 66192 46059
rect 65322 45997 65374 46007
rect 63406 45657 63458 45686
rect 63401 45643 63465 45657
rect 63401 45634 63405 45643
rect 60004 45587 63405 45634
rect 63461 45634 63465 45643
rect 66999 45634 67051 46118
rect 63461 45587 67051 45634
rect 94908 45834 94993 45855
rect 94908 45812 94924 45834
rect 94976 45812 94993 45834
rect 94908 45756 94922 45812
rect 94978 45756 94993 45812
rect 94908 45732 94924 45756
rect 94976 45732 94993 45756
rect 94908 45676 94922 45732
rect 94978 45676 94993 45732
rect 94908 45654 94924 45676
rect 94976 45654 94993 45676
rect 94908 45633 94993 45654
rect 96435 45854 96521 45866
rect 96435 45840 96452 45854
rect 96504 45840 96521 45854
rect 96435 45784 96450 45840
rect 96506 45784 96521 45840
rect 96435 45760 96452 45784
rect 96504 45760 96521 45784
rect 96435 45704 96450 45760
rect 96506 45704 96521 45760
rect 96435 45680 96452 45704
rect 96504 45680 96521 45704
rect 96435 45624 96450 45680
rect 96506 45624 96521 45680
rect 60004 45582 67051 45587
rect 92246 45603 92310 45617
rect 63401 45573 63465 45582
rect 92246 45547 92250 45603
rect 92306 45547 92310 45603
rect 96435 45610 96452 45624
rect 96504 45610 96521 45624
rect 96435 45598 96521 45610
rect 92246 45533 92310 45547
rect 92571 45397 92635 45411
rect 92571 45395 92575 45397
rect 92569 45343 92575 45395
rect 92571 45341 92575 45343
rect 92631 45395 92635 45397
rect 93033 45395 93085 45566
rect 92631 45343 93085 45395
rect 92631 45341 92635 45343
rect 92571 45327 92635 45341
rect 99948 45173 103282 45210
rect 99948 45171 99987 45173
rect 100043 45171 100067 45173
rect 100123 45171 100147 45173
rect 100203 45171 100227 45173
rect 100283 45171 100307 45173
rect 100363 45171 100387 45173
rect 100443 45171 100467 45173
rect 100523 45171 100547 45173
rect 100603 45171 100627 45173
rect 100683 45171 100707 45173
rect 100763 45171 100787 45173
rect 100843 45171 100867 45173
rect 100923 45171 100947 45173
rect 101003 45171 101027 45173
rect 101083 45171 101107 45173
rect 101163 45171 101187 45173
rect 101243 45171 101267 45173
rect 101323 45171 101347 45173
rect 101403 45171 101427 45173
rect 101483 45171 101507 45173
rect 101563 45171 101587 45173
rect 101643 45171 101667 45173
rect 101723 45171 101747 45173
rect 101803 45171 101827 45173
rect 101883 45171 101907 45173
rect 101963 45171 101987 45173
rect 102043 45171 102067 45173
rect 102123 45171 102147 45173
rect 102203 45171 102227 45173
rect 102283 45171 102307 45173
rect 102363 45171 102387 45173
rect 102443 45171 102467 45173
rect 102523 45171 102547 45173
rect 102603 45171 102627 45173
rect 102683 45171 102707 45173
rect 102763 45171 102787 45173
rect 102843 45171 102867 45173
rect 102923 45171 102947 45173
rect 103003 45171 103027 45173
rect 103083 45171 103107 45173
rect 103163 45171 103187 45173
rect 103243 45171 103282 45173
rect 99948 45119 99957 45171
rect 100137 45119 100147 45171
rect 100203 45119 100213 45171
rect 100457 45119 100467 45171
rect 100523 45119 100533 45171
rect 100777 45119 100787 45171
rect 100843 45119 100853 45171
rect 101097 45119 101107 45171
rect 101163 45119 101173 45171
rect 101417 45119 101427 45171
rect 101483 45119 101493 45171
rect 101737 45119 101747 45171
rect 101803 45119 101813 45171
rect 102057 45119 102067 45171
rect 102123 45119 102133 45171
rect 102377 45119 102387 45171
rect 102443 45119 102453 45171
rect 102697 45119 102707 45171
rect 102763 45119 102773 45171
rect 103017 45119 103027 45171
rect 103083 45119 103093 45171
rect 103273 45119 103282 45171
rect 99948 45117 99987 45119
rect 100043 45117 100067 45119
rect 100123 45117 100147 45119
rect 100203 45117 100227 45119
rect 100283 45117 100307 45119
rect 100363 45117 100387 45119
rect 100443 45117 100467 45119
rect 100523 45117 100547 45119
rect 100603 45117 100627 45119
rect 100683 45117 100707 45119
rect 100763 45117 100787 45119
rect 100843 45117 100867 45119
rect 100923 45117 100947 45119
rect 101003 45117 101027 45119
rect 101083 45117 101107 45119
rect 101163 45117 101187 45119
rect 101243 45117 101267 45119
rect 101323 45117 101347 45119
rect 101403 45117 101427 45119
rect 101483 45117 101507 45119
rect 101563 45117 101587 45119
rect 101643 45117 101667 45119
rect 101723 45117 101747 45119
rect 101803 45117 101827 45119
rect 101883 45117 101907 45119
rect 101963 45117 101987 45119
rect 102043 45117 102067 45119
rect 102123 45117 102147 45119
rect 102203 45117 102227 45119
rect 102283 45117 102307 45119
rect 102363 45117 102387 45119
rect 102443 45117 102467 45119
rect 102523 45117 102547 45119
rect 102603 45117 102627 45119
rect 102683 45117 102707 45119
rect 102763 45117 102787 45119
rect 102843 45117 102867 45119
rect 102923 45117 102947 45119
rect 103003 45117 103027 45119
rect 103083 45117 103107 45119
rect 103163 45117 103187 45119
rect 103243 45117 103282 45119
rect 99948 45081 103282 45117
rect 71782 45045 71846 45059
rect 63406 44989 63458 45019
rect 71782 44989 71786 45045
rect 71842 44989 71846 45045
rect 61491 44967 61543 44977
rect 63404 44975 63468 44989
rect 63404 44967 63408 44975
rect 61481 44915 61491 44967
rect 61543 44919 63408 44967
rect 63464 44967 63468 44975
rect 65322 44967 65374 44977
rect 71782 44975 71846 44989
rect 63464 44919 65322 44967
rect 61543 44915 65322 44919
rect 65374 44915 65384 44967
rect 61491 44905 61543 44915
rect 63404 44905 63468 44915
rect 65322 44905 65374 44915
rect 56123 44677 56127 44733
rect 56183 44677 56187 44733
rect 56123 44663 56187 44677
rect 80764 44238 80828 44248
rect 79861 44232 80828 44238
rect 79861 44180 80770 44232
rect 80822 44180 80828 44232
rect 79861 44174 80828 44180
rect 56650 44131 56714 44141
rect 62488 44131 62552 44141
rect 66488 44131 66552 44141
rect 69467 44131 69595 44143
rect 42910 39332 42946 39388
rect 43002 39332 43038 39388
rect 42910 39286 43038 39332
rect 46124 44127 69606 44131
rect 46124 44125 69473 44127
rect 46124 44073 56656 44125
rect 56708 44073 62494 44125
rect 62546 44073 66494 44125
rect 66546 44073 69473 44125
rect 46124 44061 69473 44073
rect 46124 44009 56656 44061
rect 56708 44009 62494 44061
rect 62546 44009 66494 44061
rect 66546 44011 69473 44061
rect 69589 44011 69606 44127
rect 66546 44009 69606 44011
rect 46124 44003 69606 44009
rect 44030 38159 44094 38173
rect 44030 38103 44034 38159
rect 44090 38103 44094 38159
rect 44030 38089 44094 38103
rect 46124 34241 46252 44003
rect 56650 43993 56714 44003
rect 62488 43993 62552 44003
rect 66488 43993 66552 44003
rect 69467 43995 69595 44003
rect 57145 43531 57209 43545
rect 57145 43475 57149 43531
rect 57205 43475 57209 43531
rect 56338 43230 56402 43244
rect 56338 43174 56342 43230
rect 56398 43174 56402 43230
rect 56338 43071 56402 43174
rect 57145 43073 57209 43475
rect 58778 43432 58842 43442
rect 64488 43432 64552 43442
rect 68389 43432 68517 43444
rect 58778 43428 68546 43432
rect 58778 43426 68395 43428
rect 58778 43374 58784 43426
rect 58836 43374 64494 43426
rect 64546 43374 68395 43426
rect 58778 43362 68395 43374
rect 58778 43310 58784 43362
rect 58836 43310 60495 43362
rect 60547 43310 64494 43362
rect 64546 43312 68395 43362
rect 68511 43312 68546 43428
rect 64546 43310 68546 43312
rect 58778 43304 68546 43310
rect 71781 43345 71845 43359
rect 58778 43294 58842 43304
rect 60489 43294 60553 43304
rect 64488 43294 64552 43304
rect 68389 43296 68517 43304
rect 71781 43289 71785 43345
rect 71841 43289 71845 43345
rect 71781 43275 71845 43289
rect 61951 43190 62288 43205
rect 61951 43180 61971 43190
rect 62267 43180 62288 43190
rect 60155 43124 60219 43138
rect 60155 43068 60159 43124
rect 60215 43068 60219 43124
rect 60155 43054 60219 43068
rect 61951 43064 61965 43180
rect 62273 43064 62288 43180
rect 61951 43054 61971 43064
rect 62267 43054 62288 43064
rect 64179 43124 64243 43138
rect 64179 43068 64183 43124
rect 64239 43068 64243 43124
rect 64179 43054 64243 43068
rect 66075 43124 66139 43138
rect 66075 43068 66079 43124
rect 66135 43068 66139 43124
rect 66075 43054 66139 43068
rect 67326 43076 67390 43090
rect 61951 43039 62288 43054
rect 67326 43020 67330 43076
rect 67386 43020 67390 43076
rect 67326 43006 67390 43020
rect 78065 43084 78129 43094
rect 79861 43084 79925 44174
rect 80764 44164 80828 44174
rect 80783 43400 80847 43414
rect 80783 43344 80787 43400
rect 80843 43344 80847 43400
rect 80783 43330 80847 43344
rect 78065 43080 79925 43084
rect 78065 43024 78069 43080
rect 78125 43024 79925 43080
rect 78065 43020 79925 43024
rect 78065 43010 78129 43020
rect 62801 42928 62865 42942
rect 62801 42872 62805 42928
rect 62861 42872 62865 42928
rect 62801 42858 62865 42872
rect 64800 42928 64864 42942
rect 64800 42872 64804 42928
rect 64860 42872 64864 42928
rect 64800 42858 64864 42872
rect 65374 42736 65438 42750
rect 61993 42669 62057 42683
rect 61993 42613 61997 42669
rect 62053 42613 62057 42669
rect 61993 42599 62057 42613
rect 63991 42669 64055 42683
rect 63991 42613 63995 42669
rect 64051 42613 64055 42669
rect 65374 42680 65378 42736
rect 65434 42680 65438 42736
rect 65374 42666 65438 42680
rect 70668 42706 70732 42720
rect 70668 42650 70672 42706
rect 70728 42650 70732 42706
rect 70668 42636 70732 42650
rect 63991 42599 64055 42613
rect 79861 42450 79925 43020
rect 80752 42450 80816 42460
rect 79861 42444 80816 42450
rect 79861 42392 80758 42444
rect 80810 42392 80816 42444
rect 79861 42386 80816 42392
rect 80752 42376 80816 42386
rect 60801 42330 60865 42344
rect 60801 42274 60805 42330
rect 60861 42274 60865 42330
rect 60801 42260 60865 42274
rect 66800 42330 66864 42344
rect 66800 42274 66804 42330
rect 66860 42274 66864 42330
rect 66800 42260 66864 42274
rect 59992 42049 60056 42063
rect 59992 41993 59996 42049
rect 60052 41993 60056 42049
rect 59992 41979 60056 41993
rect 65993 42049 66057 42063
rect 65993 41993 65997 42049
rect 66053 41993 66057 42049
rect 65993 41979 66057 41993
rect 57327 41790 57391 41804
rect 57327 41734 57331 41790
rect 57387 41734 57391 41790
rect 57327 41720 57391 41734
rect 71783 41560 71847 41574
rect 56273 41543 56337 41557
rect 56273 41487 56277 41543
rect 56333 41487 56337 41543
rect 71783 41504 71787 41560
rect 71843 41504 71847 41560
rect 71783 41490 71847 41504
rect 80783 41570 80847 41584
rect 80783 41514 80787 41570
rect 80843 41514 80847 41570
rect 80783 41500 80847 41514
rect 56273 41473 56337 41487
rect 64487 41381 64551 41391
rect 66490 41381 66554 41391
rect 70979 41381 71043 41391
rect 64487 41375 71056 41381
rect 64487 41323 64493 41375
rect 64545 41323 66496 41375
rect 66548 41323 70985 41375
rect 71037 41323 71056 41375
rect 61389 41307 61453 41321
rect 56649 41243 56713 41253
rect 58778 41243 58842 41253
rect 46615 41237 58842 41243
rect 61389 41251 61393 41307
rect 61449 41251 61453 41307
rect 61389 41237 61453 41251
rect 63321 41307 63385 41321
rect 63321 41251 63325 41307
rect 63381 41251 63385 41307
rect 63321 41237 63385 41251
rect 64487 41311 71056 41323
rect 64487 41259 64493 41311
rect 64545 41259 66496 41311
rect 66548 41259 70985 41311
rect 71037 41259 71056 41311
rect 64487 41253 71056 41259
rect 64487 41243 64551 41253
rect 66490 41243 66554 41253
rect 70979 41243 71043 41253
rect 46615 41185 56655 41237
rect 56707 41185 58784 41237
rect 58836 41185 58842 41237
rect 46615 41175 58842 41185
rect 46615 41119 46682 41175
rect 46738 41173 58842 41175
rect 46738 41121 56655 41173
rect 56707 41121 58784 41173
rect 58836 41121 58842 41173
rect 46738 41119 58842 41121
rect 46615 41114 58842 41119
rect 46678 41105 46742 41114
rect 56649 41105 56713 41114
rect 58778 41105 58842 41114
rect 70697 41105 70761 41115
rect 71784 41105 71848 41115
rect 70697 41101 71848 41105
rect 70697 41045 70701 41101
rect 70757 41099 71848 41101
rect 70757 41047 71790 41099
rect 71842 41047 71848 41099
rect 70757 41045 71848 41047
rect 70697 41041 71848 41045
rect 70697 41031 70761 41041
rect 71784 41031 71848 41041
rect 60487 40888 60551 40898
rect 62487 40888 62551 40898
rect 70371 40888 70435 40898
rect 60487 40882 70445 40888
rect 60487 40830 60493 40882
rect 60545 40830 62493 40882
rect 62545 40830 70377 40882
rect 70429 40830 70445 40882
rect 60487 40818 70445 40830
rect 60487 40766 60493 40818
rect 60545 40766 62493 40818
rect 62545 40766 70377 40818
rect 70429 40766 70445 40818
rect 60487 40760 70445 40766
rect 60487 40750 60551 40760
rect 62487 40750 62551 40760
rect 70371 40750 70435 40760
rect 57345 40454 68233 40478
rect 46679 40310 46743 40320
rect 53168 40310 53232 40320
rect 46679 40306 53232 40310
rect 46679 40250 46683 40306
rect 46739 40304 53232 40306
rect 46739 40252 53174 40304
rect 53226 40252 53232 40304
rect 46739 40250 53232 40252
rect 57345 40274 57355 40454
rect 68223 40274 68233 40454
rect 57345 40250 68233 40274
rect 46679 40246 53232 40250
rect 46679 40236 46743 40246
rect 53168 40236 53232 40246
rect 51308 39726 51372 39740
rect 51308 39670 51312 39726
rect 51368 39670 51372 39726
rect 51308 39656 51372 39670
rect 53180 39157 53232 40236
rect 57122 40184 57281 40221
rect 54086 39472 54150 39486
rect 54086 39416 54090 39472
rect 54146 39416 54150 39472
rect 54086 39402 54150 39416
rect 52068 38685 52704 38737
rect 52068 38433 52120 38685
rect 52192 38453 52262 38478
rect 52192 38431 52201 38453
rect 52253 38431 52262 38453
rect 52192 38375 52199 38431
rect 52255 38375 52262 38431
rect 52192 38351 52201 38375
rect 52253 38351 52262 38375
rect 52192 38295 52199 38351
rect 52255 38295 52262 38351
rect 52192 38273 52201 38295
rect 52253 38273 52262 38295
rect 52192 38248 52262 38273
rect 50550 38157 50614 38173
rect 50550 38105 50556 38157
rect 50608 38105 50614 38157
rect 50550 36908 50614 38105
rect 52177 37996 52261 38030
rect 52177 37982 52193 37996
rect 52245 37982 52261 37996
rect 52177 37926 52191 37982
rect 52247 37926 52261 37982
rect 52177 37902 52193 37926
rect 52245 37902 52261 37926
rect 52177 37846 52191 37902
rect 52247 37846 52261 37902
rect 52177 37822 52193 37846
rect 52245 37822 52261 37846
rect 52177 37766 52191 37822
rect 52247 37766 52261 37822
rect 52177 37752 52193 37766
rect 52245 37752 52261 37766
rect 52177 37718 52261 37752
rect 52088 37619 52363 37671
rect 50550 36856 50556 36908
rect 50608 36856 50614 36908
rect 50550 36840 50614 36856
rect 51243 36908 51307 36924
rect 51243 36856 51249 36908
rect 51301 36856 51307 36908
rect 51243 36235 51307 36856
rect 51243 36183 51249 36235
rect 51301 36183 51307 36235
rect 51243 36167 51307 36183
rect 51249 34965 51301 34975
rect 50683 34912 50991 34964
rect 50683 34723 50735 34912
rect 50932 34845 51157 34865
rect 50932 34789 50936 34845
rect 50992 34843 51016 34845
rect 51072 34843 51096 34845
rect 51006 34791 51016 34843
rect 51072 34791 51082 34843
rect 50992 34789 51016 34791
rect 51072 34789 51096 34791
rect 51152 34789 51157 34845
rect 50932 34770 51157 34789
rect 50683 34671 50990 34723
rect 46124 34185 46128 34241
rect 46184 34185 46252 34241
rect 46124 34161 46252 34185
rect 50938 34236 50990 34671
rect 51249 34434 51301 34913
rect 51387 34844 51693 34870
rect 51387 34788 51392 34844
rect 51448 34842 51472 34844
rect 51528 34842 51552 34844
rect 51608 34842 51632 34844
rect 51470 34790 51472 34842
rect 51534 34790 51546 34842
rect 51608 34790 51610 34842
rect 51448 34788 51472 34790
rect 51528 34788 51552 34790
rect 51608 34788 51632 34790
rect 51688 34788 51693 34844
rect 51387 34763 51693 34788
rect 51249 34423 51302 34434
rect 51301 34371 51302 34423
rect 51249 34361 51302 34371
rect 50938 34222 51002 34236
rect 50938 34166 50942 34222
rect 50998 34166 51002 34222
rect 50938 34152 51002 34166
rect 50938 33739 50990 34152
rect 50711 33687 50990 33739
rect 50711 33475 50763 33687
rect 50927 33602 51165 33624
rect 50927 33546 50938 33602
rect 50994 33600 51018 33602
rect 51074 33600 51098 33602
rect 51008 33548 51018 33600
rect 51074 33548 51084 33600
rect 50994 33546 51018 33548
rect 51074 33546 51098 33548
rect 51154 33546 51165 33602
rect 50927 33525 51165 33546
rect 50711 33423 50984 33475
rect 51249 33474 51301 34361
rect 51746 34236 51798 34957
rect 52311 34265 52363 37619
rect 52652 34265 52704 38685
rect 53180 38161 53232 39105
rect 56416 39158 56468 39168
rect 53950 39002 54033 39030
rect 53950 38988 53965 39002
rect 54017 38988 54033 39002
rect 53950 38932 53963 38988
rect 54019 38932 54033 38988
rect 53950 38908 53965 38932
rect 54017 38908 54033 38932
rect 53950 38852 53963 38908
rect 54019 38852 54033 38908
rect 53950 38828 53965 38852
rect 54017 38828 54033 38852
rect 53950 38772 53963 38828
rect 54019 38772 54033 38828
rect 53950 38758 53965 38772
rect 54017 38758 54033 38772
rect 53950 38731 54033 38758
rect 54071 38662 54135 38676
rect 54071 38606 54075 38662
rect 54131 38606 54135 38662
rect 54071 38592 54135 38606
rect 53180 36657 53232 38109
rect 54496 37155 54560 37169
rect 54496 37099 54500 37155
rect 54556 37099 54560 37155
rect 54496 37085 54560 37099
rect 55286 37139 55369 37165
rect 55286 37083 55299 37139
rect 55355 37083 55369 37139
rect 55286 37073 55369 37083
rect 55286 37059 55301 37073
rect 55353 37059 55369 37073
rect 55286 37003 55299 37059
rect 55355 37003 55369 37059
rect 55286 36979 55301 37003
rect 55353 36979 55369 37003
rect 55286 36923 55299 36979
rect 55355 36923 55369 36979
rect 55286 36899 55301 36923
rect 55353 36899 55369 36923
rect 55286 36843 55299 36899
rect 55355 36843 55369 36899
rect 55286 36829 55301 36843
rect 55353 36829 55369 36843
rect 55286 36819 55369 36829
rect 55286 36763 55299 36819
rect 55355 36763 55369 36819
rect 55286 36738 55369 36763
rect 51733 34222 51798 34236
rect 51733 34220 51737 34222
rect 51731 34168 51737 34220
rect 51733 34166 51737 34168
rect 51793 34166 51798 34222
rect 52305 34251 52369 34265
rect 52305 34195 52309 34251
rect 52365 34195 52369 34251
rect 52305 34181 52369 34195
rect 52646 34251 52710 34265
rect 52646 34195 52650 34251
rect 52706 34195 52710 34251
rect 52646 34181 52710 34195
rect 51733 34152 51798 34166
rect 51386 33602 51695 33627
rect 51386 33600 51392 33602
rect 51448 33600 51472 33602
rect 51528 33600 51552 33602
rect 51608 33600 51632 33602
rect 51688 33600 51695 33602
rect 51448 33548 51450 33600
rect 51630 33548 51632 33600
rect 51694 33548 51695 33600
rect 51386 33546 51392 33548
rect 51448 33546 51472 33548
rect 51528 33546 51552 33548
rect 51608 33546 51632 33548
rect 51688 33546 51695 33548
rect 51386 33521 51695 33546
rect 51746 33428 51798 34152
rect 51249 33412 51301 33422
rect 40313 31569 40349 31625
rect 40405 31569 40441 31625
rect 51241 32190 51305 32206
rect 51241 32138 51247 32190
rect 51299 32138 51305 32190
rect 40313 31523 40441 31569
rect 50529 31607 50593 31623
rect 50529 31555 50535 31607
rect 50587 31555 50593 31607
rect 49880 31253 50343 31275
rect 49880 31037 49883 31253
rect 50339 31037 50343 31253
rect 49880 31015 50343 31037
rect 31466 30763 32178 30815
rect 31573 30682 31648 30701
rect 31573 30668 31584 30682
rect 31636 30668 31648 30682
rect 31573 30612 31582 30668
rect 31638 30612 31648 30668
rect 31573 30588 31584 30612
rect 31636 30588 31648 30612
rect 31573 30532 31582 30588
rect 31638 30532 31648 30588
rect 31573 30508 31584 30532
rect 31636 30508 31648 30532
rect 31573 30452 31582 30508
rect 31638 30452 31648 30508
rect 31573 30438 31584 30452
rect 31636 30438 31648 30452
rect 31573 30420 31648 30438
rect 38843 30321 38907 30335
rect 38843 30265 38847 30321
rect 38903 30265 38907 30321
rect 38843 30251 38907 30265
rect 44019 30331 44083 30345
rect 44019 30275 44023 30331
rect 44079 30275 44083 30331
rect 44019 30261 44083 30275
rect 50529 30329 50593 31555
rect 51241 31611 51305 32138
rect 51241 31559 51247 31611
rect 51299 31559 51305 31611
rect 51241 31543 51305 31559
rect 52311 30825 52363 34181
rect 52058 30773 52363 30825
rect 52177 30713 52258 30727
rect 52177 30657 52189 30713
rect 52245 30657 52258 30713
rect 52177 30635 52191 30657
rect 52243 30635 52258 30657
rect 52177 30633 52258 30635
rect 52177 30577 52189 30633
rect 52245 30577 52258 30633
rect 52177 30571 52191 30577
rect 52243 30571 52258 30577
rect 52177 30559 52258 30571
rect 52177 30553 52191 30559
rect 52243 30553 52258 30559
rect 52177 30497 52189 30553
rect 52245 30497 52258 30553
rect 52177 30495 52258 30497
rect 52177 30473 52191 30495
rect 52243 30473 52258 30495
rect 52177 30417 52189 30473
rect 52245 30417 52258 30473
rect 52177 30404 52258 30417
rect 50529 30277 50535 30329
rect 50587 30277 50593 30329
rect 50529 30261 50593 30277
rect 31572 30195 31647 30206
rect 31572 30181 31583 30195
rect 31635 30181 31647 30195
rect 31572 30125 31581 30181
rect 31637 30125 31647 30181
rect 31572 30101 31583 30125
rect 31635 30101 31647 30125
rect 31572 30045 31581 30101
rect 31637 30045 31647 30101
rect 31572 30021 31583 30045
rect 31635 30021 31647 30045
rect 29848 29958 30312 30009
rect 29929 29957 30312 29958
rect 31572 29965 31581 30021
rect 31637 29965 31647 30021
rect 52187 30168 52253 30195
rect 52187 30146 52194 30168
rect 52246 30146 52253 30168
rect 52187 30090 52192 30146
rect 52248 30090 52253 30146
rect 52187 30066 52194 30090
rect 52246 30066 52253 30090
rect 31572 29951 31583 29965
rect 31635 29951 31647 29965
rect 31572 29941 31647 29951
rect 52065 29848 52117 30016
rect 52187 30010 52192 30066
rect 52248 30010 52253 30066
rect 52187 29988 52194 30010
rect 52246 29988 52253 30010
rect 52187 29962 52253 29988
rect 52652 29848 52704 34181
rect 53180 33459 53232 36605
rect 55596 36427 55660 36441
rect 55596 36371 55600 36427
rect 55656 36371 55660 36427
rect 54209 36346 54273 36360
rect 55596 36357 55660 36371
rect 54209 36290 54213 36346
rect 54269 36290 54273 36346
rect 54209 36276 54273 36290
rect 55168 35553 55232 35567
rect 55168 35497 55172 35553
rect 55228 35497 55232 35553
rect 55168 35483 55232 35497
rect 55335 35544 55401 35561
rect 55335 35488 55340 35544
rect 55396 35488 55401 35544
rect 55335 35478 55401 35488
rect 55335 35464 55342 35478
rect 55394 35464 55401 35478
rect 55335 35408 55340 35464
rect 55396 35408 55401 35464
rect 55335 35384 55342 35408
rect 55394 35384 55401 35408
rect 55335 35328 55340 35384
rect 55396 35328 55401 35384
rect 55335 35304 55342 35328
rect 55394 35304 55401 35328
rect 55335 35248 55340 35304
rect 55396 35248 55401 35304
rect 55335 35234 55342 35248
rect 55394 35234 55401 35248
rect 55335 35224 55401 35234
rect 55335 35168 55340 35224
rect 55396 35168 55401 35224
rect 55335 35152 55401 35168
rect 53180 33397 53232 33407
rect 53679 35056 53731 35066
rect 52065 29796 52704 29848
rect 53679 31857 53731 35004
rect 55596 34801 55660 34815
rect 54882 34747 54946 34761
rect 54882 34691 54886 34747
rect 54942 34691 54946 34747
rect 55596 34745 55600 34801
rect 55656 34745 55660 34801
rect 55596 34731 55660 34745
rect 54882 34677 54946 34691
rect 56416 34424 56468 39106
rect 55168 33955 55232 33969
rect 55168 33899 55172 33955
rect 55228 33899 55232 33955
rect 55168 33885 55232 33899
rect 55335 33941 55399 33962
rect 55335 33885 55339 33941
rect 55395 33885 55399 33941
rect 55335 33875 55399 33885
rect 55335 33861 55341 33875
rect 55393 33861 55399 33875
rect 55335 33805 55339 33861
rect 55395 33805 55399 33861
rect 55335 33781 55341 33805
rect 55393 33781 55399 33805
rect 55335 33725 55339 33781
rect 55395 33725 55399 33781
rect 55335 33701 55341 33725
rect 55393 33701 55399 33725
rect 55335 33645 55339 33701
rect 55395 33645 55399 33701
rect 55335 33631 55341 33645
rect 55393 33631 55399 33645
rect 55335 33621 55399 33631
rect 55335 33565 55339 33621
rect 55395 33565 55399 33621
rect 55335 33544 55399 33565
rect 55945 33457 55997 33473
rect 54882 33147 54946 33161
rect 54882 33091 54886 33147
rect 54942 33091 54946 33147
rect 54882 33077 54946 33091
rect 55596 33143 55660 33157
rect 55596 33087 55600 33143
rect 55656 33087 55660 33143
rect 55596 33073 55660 33087
rect 54496 32353 54560 32367
rect 54496 32297 54500 32353
rect 54556 32297 54560 32353
rect 54496 32283 54560 32297
rect 55336 32340 55404 32362
rect 55336 32284 55342 32340
rect 55398 32284 55404 32340
rect 55336 32274 55404 32284
rect 55336 32260 55344 32274
rect 55396 32260 55404 32274
rect 55336 32204 55342 32260
rect 55398 32204 55404 32260
rect 55336 32180 55344 32204
rect 55396 32180 55404 32204
rect 55336 32124 55342 32180
rect 55398 32124 55404 32180
rect 55336 32100 55344 32124
rect 55396 32100 55404 32124
rect 55336 32044 55342 32100
rect 55398 32044 55404 32100
rect 55336 32030 55344 32044
rect 55396 32030 55404 32044
rect 55336 32020 55404 32030
rect 55336 31964 55342 32020
rect 55398 31964 55404 32020
rect 55336 31942 55404 31964
rect 53679 30332 53731 31805
rect 55945 31857 55997 33405
rect 55596 31604 55660 31618
rect 54209 31545 54273 31559
rect 54209 31489 54213 31545
rect 54269 31489 54273 31545
rect 55596 31548 55600 31604
rect 55656 31548 55660 31604
rect 55596 31534 55660 31548
rect 54209 31475 54273 31489
rect 55596 31260 55660 31290
rect 55596 31246 55602 31260
rect 55654 31246 55660 31260
rect 55596 31190 55600 31246
rect 55656 31190 55660 31246
rect 55596 31166 55602 31190
rect 55654 31166 55660 31190
rect 55596 31110 55600 31166
rect 55656 31110 55660 31166
rect 55596 31086 55602 31110
rect 55654 31086 55660 31110
rect 55596 31030 55600 31086
rect 55656 31030 55660 31086
rect 55596 31016 55602 31030
rect 55654 31016 55660 31030
rect 55596 30986 55660 31016
rect 55596 30469 55660 30483
rect 55596 30413 55600 30469
rect 55656 30413 55660 30469
rect 55596 30399 55660 30413
rect 53679 29745 53731 30280
rect 54044 30060 54108 30074
rect 54044 30004 54048 30060
rect 54104 30004 54108 30060
rect 54044 29990 54108 30004
rect 53679 29079 53731 29693
rect 53901 29580 53984 29609
rect 53901 29566 53916 29580
rect 53968 29566 53984 29580
rect 53901 29510 53914 29566
rect 53970 29510 53984 29566
rect 53901 29486 53916 29510
rect 53968 29486 53984 29510
rect 53901 29430 53914 29486
rect 53970 29430 53984 29486
rect 53901 29406 53916 29430
rect 53968 29406 53984 29430
rect 53901 29350 53914 29406
rect 53970 29350 53984 29406
rect 53901 29336 53916 29350
rect 53968 29336 53984 29350
rect 53901 29308 53984 29336
rect 54066 29251 54130 29265
rect 54066 29195 54070 29251
rect 54126 29195 54130 29251
rect 54066 29181 54130 29195
rect 55945 29151 55997 31805
rect 56416 29745 56468 34372
rect 56416 29683 56468 29693
rect 56815 36659 56867 36669
rect 56815 35057 56867 36607
rect 55945 29089 55997 29099
rect 46328 29069 46392 29079
rect 53667 29069 53731 29079
rect 46328 29065 53731 29069
rect 46328 29009 46332 29065
rect 46388 29063 53731 29065
rect 46388 29011 53673 29063
rect 53725 29011 53731 29063
rect 46388 29009 53731 29011
rect 46328 29005 53731 29009
rect 46328 28995 46392 29005
rect 53667 28995 53731 29005
rect 56815 27811 56867 35005
rect 57122 34688 57133 40184
rect 57269 34688 57281 40184
rect 68333 40195 68493 40216
rect 68333 38459 68345 40195
rect 68481 38459 68493 40195
rect 80780 39806 80844 39820
rect 71759 39729 71865 39765
rect 80780 39750 80784 39806
rect 80840 39750 80844 39806
rect 80780 39736 80844 39750
rect 71759 39673 71784 39729
rect 71840 39673 71865 39729
rect 71759 39638 71865 39673
rect 78022 39514 78086 39528
rect 78022 39458 78026 39514
rect 78082 39458 78086 39514
rect 78022 39444 78086 39458
rect 71784 39246 71848 39260
rect 71784 39190 71788 39246
rect 71844 39190 71848 39246
rect 71784 39176 71848 39190
rect 68333 38438 68493 38459
rect 80780 38015 80844 38029
rect 68351 37968 68478 37986
rect 68351 37020 68356 37968
rect 68472 37020 68478 37968
rect 71779 37983 71843 37997
rect 71779 37927 71783 37983
rect 71839 37927 71843 37983
rect 80780 37959 80784 38015
rect 80840 37959 80844 38015
rect 80780 37945 80844 37959
rect 71779 37913 71843 37927
rect 70730 37550 70794 37560
rect 71784 37550 71848 37560
rect 70730 37546 71848 37550
rect 70730 37490 70734 37546
rect 70790 37544 71848 37546
rect 70790 37492 71790 37544
rect 71842 37492 71848 37544
rect 70790 37490 71848 37492
rect 70730 37486 71848 37490
rect 70730 37476 70794 37486
rect 71784 37476 71848 37486
rect 80779 37028 80843 37038
rect 68351 37002 68478 37020
rect 80188 37022 80843 37028
rect 80188 36970 80785 37022
rect 80837 36970 80843 37022
rect 80188 36964 80843 36970
rect 71796 36198 71860 36212
rect 68337 36132 68492 36161
rect 68337 35356 68346 36132
rect 68482 35356 68492 36132
rect 71796 36142 71800 36198
rect 71856 36142 71860 36198
rect 71796 36128 71860 36142
rect 78079 35928 78143 35938
rect 80188 35928 80252 36964
rect 80779 36954 80843 36964
rect 80785 36208 80849 36222
rect 80785 36152 80789 36208
rect 80845 36152 80849 36208
rect 80785 36138 80849 36152
rect 78062 35924 80847 35928
rect 78062 35868 78083 35924
rect 78139 35868 80847 35924
rect 78062 35864 80847 35868
rect 78079 35854 78143 35864
rect 70793 35698 70857 35708
rect 71786 35698 71850 35708
rect 70793 35694 71850 35698
rect 70793 35638 70797 35694
rect 70853 35692 71850 35694
rect 70853 35640 71792 35692
rect 71844 35640 71850 35692
rect 70853 35638 71850 35640
rect 70793 35634 71850 35638
rect 70793 35624 70857 35634
rect 71786 35624 71850 35634
rect 80783 35535 80847 35864
rect 80783 35483 80789 35535
rect 80841 35483 80847 35535
rect 80783 35467 80847 35483
rect 68337 35328 68492 35356
rect 57122 34652 57281 34688
rect 63577 34536 68312 34569
rect 63577 34400 63596 34536
rect 68292 34400 68312 34536
rect 63577 34368 68312 34400
rect 71785 34401 71849 34415
rect 71785 34345 71789 34401
rect 71845 34345 71849 34401
rect 71785 34331 71849 34345
rect 80785 34398 80849 34412
rect 80785 34342 80789 34398
rect 80845 34342 80849 34398
rect 80785 34328 80849 34342
rect 62317 33440 62370 33450
rect 81638 33440 81702 33456
rect 62317 33439 81644 33440
rect 62369 33388 81644 33439
rect 81696 33388 81702 33440
rect 62369 33387 81702 33388
rect 62317 33377 62370 33387
rect 81638 33372 81702 33387
rect 93160 33172 93224 33186
rect 80302 31867 80355 31877
rect 74865 31866 80355 31867
rect 74865 31814 80302 31866
rect 80354 31814 80355 31866
rect 74865 31739 74918 31814
rect 80302 31804 80355 31814
rect 70014 31686 74918 31739
rect 82589 31673 82653 33138
rect 92936 33118 93164 33172
rect 92583 32549 92647 32563
rect 92583 32493 92587 32549
rect 92643 32493 92647 32549
rect 92583 32479 92647 32493
rect 92936 32422 92990 33118
rect 93160 33116 93164 33118
rect 93220 33116 93224 33172
rect 93160 33102 93224 33116
rect 93725 32487 93789 32501
rect 93076 32435 93729 32487
rect 93725 32431 93729 32435
rect 93785 32431 93789 32487
rect 93725 32417 93789 32431
rect 92118 32301 92182 32315
rect 92118 32245 92122 32301
rect 92178 32245 92182 32301
rect 92118 32231 92182 32245
rect 97194 32139 97275 32153
rect 97194 32117 97208 32139
rect 97260 32117 97275 32139
rect 95669 32055 95739 32070
rect 95669 31999 95676 32055
rect 95732 31999 95739 32055
rect 95669 31993 95678 31999
rect 95730 31993 95739 31999
rect 95669 31981 95739 31993
rect 95669 31975 95678 31981
rect 95730 31975 95739 31981
rect 95669 31919 95676 31975
rect 95732 31919 95739 31975
rect 97194 32061 97206 32117
rect 97262 32061 97275 32117
rect 97194 32037 97208 32061
rect 97260 32037 97275 32061
rect 97194 31981 97206 32037
rect 97262 31981 97275 32037
rect 97194 31959 97208 31981
rect 97260 31959 97275 31981
rect 97194 31945 97275 31959
rect 93395 31897 93626 31913
rect 95669 31904 95739 31919
rect 93395 31841 93402 31897
rect 93458 31895 93482 31897
rect 93538 31895 93562 31897
rect 93472 31843 93482 31895
rect 93538 31843 93548 31895
rect 93458 31841 93482 31843
rect 93538 31841 93562 31843
rect 93618 31841 93626 31897
rect 93395 31826 93626 31841
rect 90840 31673 90904 31683
rect 82589 31667 90904 31673
rect 82589 31615 90846 31667
rect 90898 31615 90904 31667
rect 82589 31609 90904 31615
rect 90840 31599 90904 31609
rect 95662 31581 95743 31595
rect 95662 31559 95676 31581
rect 95728 31559 95743 31581
rect 95662 31503 95674 31559
rect 95730 31503 95743 31559
rect 95662 31479 95676 31503
rect 95728 31479 95743 31503
rect 95662 31423 95674 31479
rect 95730 31423 95743 31479
rect 95662 31401 95676 31423
rect 95728 31401 95743 31423
rect 95662 31387 95743 31401
rect 97181 31594 97262 31608
rect 97181 31572 97195 31594
rect 97247 31572 97262 31594
rect 97181 31516 97193 31572
rect 97249 31516 97262 31572
rect 97181 31492 97195 31516
rect 97247 31492 97262 31516
rect 97181 31436 97193 31492
rect 97249 31436 97262 31492
rect 97181 31414 97195 31436
rect 97247 31414 97262 31436
rect 97181 31400 97262 31414
rect 93456 31356 93625 31369
rect 93456 31300 93472 31356
rect 93528 31354 93552 31356
rect 93534 31302 93546 31354
rect 93528 31300 93552 31302
rect 93608 31300 93625 31356
rect 93456 31287 93625 31300
rect 92122 31241 92186 31255
rect 92122 31185 92126 31241
rect 92182 31185 92186 31241
rect 92122 31171 92186 31185
rect 99696 31237 103017 31264
rect 99696 31235 99728 31237
rect 99784 31235 99808 31237
rect 99864 31235 99888 31237
rect 99944 31235 99968 31237
rect 100024 31235 100048 31237
rect 100104 31235 100128 31237
rect 100184 31235 100208 31237
rect 100264 31235 100288 31237
rect 100344 31235 100368 31237
rect 100424 31235 100448 31237
rect 100504 31235 100528 31237
rect 100584 31235 100608 31237
rect 100664 31235 100688 31237
rect 100744 31235 100768 31237
rect 100824 31235 100848 31237
rect 100904 31235 100928 31237
rect 100984 31235 101008 31237
rect 101064 31235 101088 31237
rect 101144 31235 101168 31237
rect 101224 31235 101248 31237
rect 101304 31235 101328 31237
rect 101384 31235 101408 31237
rect 101464 31235 101488 31237
rect 101544 31235 101568 31237
rect 101624 31235 101648 31237
rect 101704 31235 101728 31237
rect 101784 31235 101808 31237
rect 101864 31235 101888 31237
rect 101944 31235 101968 31237
rect 102024 31235 102048 31237
rect 102104 31235 102128 31237
rect 102184 31235 102208 31237
rect 102264 31235 102288 31237
rect 102344 31235 102368 31237
rect 102424 31235 102448 31237
rect 102504 31235 102528 31237
rect 102584 31235 102608 31237
rect 102664 31235 102688 31237
rect 102744 31235 102768 31237
rect 102824 31235 102848 31237
rect 102904 31235 102928 31237
rect 102984 31235 103017 31237
rect 99696 31183 99698 31235
rect 99878 31183 99888 31235
rect 99944 31183 99954 31235
rect 100198 31183 100208 31235
rect 100264 31183 100274 31235
rect 100518 31183 100528 31235
rect 100584 31183 100594 31235
rect 100838 31183 100848 31235
rect 100904 31183 100914 31235
rect 101158 31183 101168 31235
rect 101224 31183 101234 31235
rect 101478 31183 101488 31235
rect 101544 31183 101554 31235
rect 101798 31183 101808 31235
rect 101864 31183 101874 31235
rect 102118 31183 102128 31235
rect 102184 31183 102194 31235
rect 102438 31183 102448 31235
rect 102504 31183 102514 31235
rect 102758 31183 102768 31235
rect 102824 31183 102834 31235
rect 103014 31183 103017 31235
rect 99696 31181 99728 31183
rect 99784 31181 99808 31183
rect 99864 31181 99888 31183
rect 99944 31181 99968 31183
rect 100024 31181 100048 31183
rect 100104 31181 100128 31183
rect 100184 31181 100208 31183
rect 100264 31181 100288 31183
rect 100344 31181 100368 31183
rect 100424 31181 100448 31183
rect 100504 31181 100528 31183
rect 100584 31181 100608 31183
rect 100664 31181 100688 31183
rect 100744 31181 100768 31183
rect 100824 31181 100848 31183
rect 100904 31181 100928 31183
rect 100984 31181 101008 31183
rect 101064 31181 101088 31183
rect 101144 31181 101168 31183
rect 101224 31181 101248 31183
rect 101304 31181 101328 31183
rect 101384 31181 101408 31183
rect 101464 31181 101488 31183
rect 101544 31181 101568 31183
rect 101624 31181 101648 31183
rect 101704 31181 101728 31183
rect 101784 31181 101808 31183
rect 101864 31181 101888 31183
rect 101944 31181 101968 31183
rect 102024 31181 102048 31183
rect 102104 31181 102128 31183
rect 102184 31181 102208 31183
rect 102264 31181 102288 31183
rect 102344 31181 102368 31183
rect 102424 31181 102448 31183
rect 102504 31181 102528 31183
rect 102584 31181 102608 31183
rect 102664 31181 102688 31183
rect 102744 31181 102768 31183
rect 102824 31181 102848 31183
rect 102904 31181 102928 31183
rect 102984 31181 103017 31183
rect 99696 31155 103017 31181
rect 92121 30972 92185 30986
rect 92121 30916 92125 30972
rect 92181 30916 92185 30972
rect 92121 30902 92185 30916
rect 93446 30808 93531 30827
rect 93446 30752 93460 30808
rect 93516 30752 93531 30808
rect 93446 30733 93531 30752
rect 97186 30803 97267 30817
rect 97186 30781 97200 30803
rect 97252 30781 97267 30803
rect 95665 30724 95743 30739
rect 95665 30694 95678 30724
rect 95730 30694 95743 30724
rect 95665 30638 95676 30694
rect 95732 30638 95743 30694
rect 95665 30608 95678 30638
rect 95730 30608 95743 30638
rect 97186 30725 97198 30781
rect 97254 30725 97267 30781
rect 97186 30701 97200 30725
rect 97252 30701 97267 30725
rect 97186 30645 97198 30701
rect 97254 30645 97267 30701
rect 97186 30623 97200 30645
rect 97252 30623 97267 30645
rect 97186 30609 97267 30623
rect 95665 30594 95743 30608
rect 81638 30334 81702 30344
rect 90828 30334 90892 30344
rect 81638 30328 90892 30334
rect 81638 30276 81644 30328
rect 81696 30276 90834 30328
rect 90886 30276 90892 30328
rect 81638 30270 90892 30276
rect 81638 30260 81702 30270
rect 90828 30260 90892 30270
rect 94065 30267 94161 30297
rect 94065 30211 94085 30267
rect 94141 30211 94161 30267
rect 94065 30181 94161 30211
rect 95657 30250 95738 30264
rect 95657 30228 95671 30250
rect 95723 30228 95738 30250
rect 95657 30172 95669 30228
rect 95725 30172 95738 30228
rect 95657 30148 95671 30172
rect 95723 30148 95738 30172
rect 95657 30092 95669 30148
rect 95725 30092 95738 30148
rect 95657 30070 95671 30092
rect 95723 30070 95738 30092
rect 95657 30056 95738 30070
rect 97186 30247 97267 30261
rect 97186 30225 97200 30247
rect 97252 30225 97267 30247
rect 97186 30169 97198 30225
rect 97254 30169 97267 30225
rect 97186 30145 97200 30169
rect 97252 30145 97267 30169
rect 97186 30089 97198 30145
rect 97254 30089 97267 30145
rect 97186 30067 97200 30089
rect 97252 30067 97267 30089
rect 97186 30053 97267 30067
rect 92121 29903 92185 29917
rect 92121 29847 92125 29903
rect 92181 29847 92185 29903
rect 92121 29833 92185 29847
rect 104567 29812 104803 29832
rect 93064 29725 93243 29739
rect 93064 29669 93085 29725
rect 93141 29723 93165 29725
rect 93147 29671 93159 29723
rect 93141 29669 93165 29671
rect 93221 29669 93243 29725
rect 93064 29656 93243 29669
rect 104567 29596 104577 29812
rect 104793 29596 104803 29812
rect 92118 29580 92182 29594
rect 92118 29524 92122 29580
rect 92178 29524 92182 29580
rect 104567 29576 104803 29596
rect 92118 29510 92182 29524
rect 97203 29423 97284 29437
rect 97203 29401 97217 29423
rect 97269 29401 97284 29423
rect 95668 29334 95742 29354
rect 95668 29304 95679 29334
rect 95731 29304 95742 29334
rect 95668 29248 95677 29304
rect 95733 29248 95742 29304
rect 95668 29218 95679 29248
rect 95731 29218 95742 29248
rect 97203 29345 97215 29401
rect 97271 29345 97284 29401
rect 97203 29321 97217 29345
rect 97269 29321 97284 29345
rect 97203 29265 97215 29321
rect 97271 29265 97284 29321
rect 97203 29243 97217 29265
rect 97269 29243 97284 29265
rect 97203 29229 97284 29243
rect 95668 29199 95742 29218
rect 93608 29177 93828 29194
rect 93608 29121 93610 29177
rect 93666 29175 93690 29177
rect 93746 29175 93770 29177
rect 93680 29123 93690 29175
rect 93746 29123 93756 29175
rect 93666 29121 93690 29123
rect 93746 29121 93770 29123
rect 93826 29121 93828 29177
rect 93608 29104 93828 29121
rect 80302 28938 80355 28948
rect 90836 28938 90889 28948
rect 80302 28937 90889 28938
rect 80354 28885 90836 28937
rect 90888 28885 90889 28937
rect 80302 28875 80355 28885
rect 90836 28875 90889 28885
rect 95656 28897 95737 28911
rect 95656 28875 95670 28897
rect 95722 28875 95737 28897
rect 95656 28819 95668 28875
rect 95724 28819 95737 28875
rect 95656 28795 95670 28819
rect 95722 28795 95737 28819
rect 95656 28739 95668 28795
rect 95724 28739 95737 28795
rect 95656 28717 95670 28739
rect 95722 28717 95737 28739
rect 95656 28703 95737 28717
rect 97186 28875 97267 28889
rect 97186 28853 97200 28875
rect 97252 28853 97267 28875
rect 97186 28797 97198 28853
rect 97254 28797 97267 28853
rect 97186 28773 97200 28797
rect 97252 28773 97267 28797
rect 97186 28717 97198 28773
rect 97254 28717 97267 28773
rect 97186 28695 97200 28717
rect 97252 28695 97267 28717
rect 97186 28681 97267 28695
rect 93458 28634 93603 28645
rect 93458 28578 93462 28634
rect 93518 28632 93542 28634
rect 93524 28580 93536 28632
rect 93518 28578 93542 28580
rect 93598 28578 93603 28634
rect 93458 28567 93603 28578
rect 92129 28510 92193 28524
rect 92129 28454 92133 28510
rect 92189 28454 92193 28510
rect 92129 28440 92193 28454
rect 99693 28238 103053 28265
rect 92118 28205 92182 28219
rect 92118 28149 92122 28205
rect 92178 28149 92182 28205
rect 99693 28182 99705 28238
rect 99761 28236 99785 28238
rect 99841 28236 99865 28238
rect 99921 28236 99945 28238
rect 100001 28236 100025 28238
rect 100081 28236 100105 28238
rect 100161 28236 100185 28238
rect 100241 28236 100265 28238
rect 100321 28236 100345 28238
rect 100401 28236 100425 28238
rect 100481 28236 100505 28238
rect 100561 28236 100585 28238
rect 100641 28236 100665 28238
rect 100721 28236 100745 28238
rect 100801 28236 100825 28238
rect 100881 28236 100905 28238
rect 100961 28236 100985 28238
rect 101041 28236 101065 28238
rect 101121 28236 101145 28238
rect 101201 28236 101225 28238
rect 101281 28236 101305 28238
rect 101361 28236 101385 28238
rect 101441 28236 101465 28238
rect 101521 28236 101545 28238
rect 101601 28236 101625 28238
rect 101681 28236 101705 28238
rect 101761 28236 101785 28238
rect 101841 28236 101865 28238
rect 101921 28236 101945 28238
rect 102001 28236 102025 28238
rect 102081 28236 102105 28238
rect 102161 28236 102185 28238
rect 102241 28236 102265 28238
rect 102321 28236 102345 28238
rect 102401 28236 102425 28238
rect 102481 28236 102505 28238
rect 102561 28236 102585 28238
rect 102641 28236 102665 28238
rect 102721 28236 102745 28238
rect 102801 28236 102825 28238
rect 102881 28236 102905 28238
rect 102961 28236 102985 28238
rect 99767 28184 99779 28236
rect 99841 28184 99843 28236
rect 100023 28184 100025 28236
rect 100087 28184 100099 28236
rect 100161 28184 100163 28236
rect 100343 28184 100345 28236
rect 100407 28184 100419 28236
rect 100481 28184 100483 28236
rect 100663 28184 100665 28236
rect 100727 28184 100739 28236
rect 100801 28184 100803 28236
rect 100983 28184 100985 28236
rect 101047 28184 101059 28236
rect 101121 28184 101123 28236
rect 101303 28184 101305 28236
rect 101367 28184 101379 28236
rect 101441 28184 101443 28236
rect 101623 28184 101625 28236
rect 101687 28184 101699 28236
rect 101761 28184 101763 28236
rect 101943 28184 101945 28236
rect 102007 28184 102019 28236
rect 102081 28184 102083 28236
rect 102263 28184 102265 28236
rect 102327 28184 102339 28236
rect 102401 28184 102403 28236
rect 102583 28184 102585 28236
rect 102647 28184 102659 28236
rect 102721 28184 102723 28236
rect 102903 28184 102905 28236
rect 102967 28184 102979 28236
rect 99761 28182 99785 28184
rect 99841 28182 99865 28184
rect 99921 28182 99945 28184
rect 100001 28182 100025 28184
rect 100081 28182 100105 28184
rect 100161 28182 100185 28184
rect 100241 28182 100265 28184
rect 100321 28182 100345 28184
rect 100401 28182 100425 28184
rect 100481 28182 100505 28184
rect 100561 28182 100585 28184
rect 100641 28182 100665 28184
rect 100721 28182 100745 28184
rect 100801 28182 100825 28184
rect 100881 28182 100905 28184
rect 100961 28182 100985 28184
rect 101041 28182 101065 28184
rect 101121 28182 101145 28184
rect 101201 28182 101225 28184
rect 101281 28182 101305 28184
rect 101361 28182 101385 28184
rect 101441 28182 101465 28184
rect 101521 28182 101545 28184
rect 101601 28182 101625 28184
rect 101681 28182 101705 28184
rect 101761 28182 101785 28184
rect 101841 28182 101865 28184
rect 101921 28182 101945 28184
rect 102001 28182 102025 28184
rect 102081 28182 102105 28184
rect 102161 28182 102185 28184
rect 102241 28182 102265 28184
rect 102321 28182 102345 28184
rect 102401 28182 102425 28184
rect 102481 28182 102505 28184
rect 102561 28182 102585 28184
rect 102641 28182 102665 28184
rect 102721 28182 102745 28184
rect 102801 28182 102825 28184
rect 102881 28182 102905 28184
rect 102961 28182 102985 28184
rect 103041 28182 103053 28238
rect 99693 28156 103053 28182
rect 92118 28135 92182 28149
rect 94066 28091 94162 28121
rect 94066 28035 94086 28091
rect 94142 28035 94162 28091
rect 94066 28005 94162 28035
rect 97193 28044 97274 28058
rect 97193 28022 97207 28044
rect 97259 28022 97274 28044
rect 97193 27966 97205 28022
rect 97261 27966 97274 28022
rect 95666 27947 95745 27966
rect 95666 27891 95677 27947
rect 95733 27891 95745 27947
rect 95666 27885 95679 27891
rect 95731 27885 95745 27891
rect 95666 27873 95745 27885
rect 95666 27867 95679 27873
rect 95731 27867 95745 27873
rect 95666 27811 95677 27867
rect 95733 27811 95745 27867
rect 97193 27942 97207 27966
rect 97259 27942 97274 27966
rect 97193 27886 97205 27942
rect 97261 27886 97274 27942
rect 97193 27864 97207 27886
rect 97259 27864 97274 27886
rect 97193 27850 97274 27864
rect 95666 27793 95745 27811
rect 56815 27749 56867 27759
rect 93453 27545 93580 27563
rect 93453 27543 93488 27545
rect 93544 27543 93580 27545
rect 93453 27491 93458 27543
rect 93574 27491 93580 27543
rect 93453 27489 93488 27491
rect 93544 27489 93580 27491
rect 93453 27471 93580 27489
rect 95659 27497 95740 27511
rect 95659 27475 95673 27497
rect 95725 27475 95740 27497
rect 95659 27419 95671 27475
rect 95727 27419 95740 27475
rect 95659 27395 95673 27419
rect 95725 27395 95740 27419
rect 95659 27339 95671 27395
rect 95727 27339 95740 27395
rect 95659 27317 95673 27339
rect 95725 27317 95740 27339
rect 95659 27303 95740 27317
rect 97183 27491 97264 27505
rect 97183 27469 97197 27491
rect 97249 27469 97264 27491
rect 97183 27413 97195 27469
rect 97251 27413 97264 27469
rect 97183 27389 97197 27413
rect 97249 27389 97264 27413
rect 97183 27333 97195 27389
rect 97251 27333 97264 27389
rect 97183 27311 97197 27333
rect 97249 27311 97264 27333
rect 97183 27297 97264 27311
rect 92125 27140 92189 27154
rect 92125 27084 92129 27140
rect 92185 27084 92189 27140
rect 92125 27070 92189 27084
rect 60764 26710 62498 26763
rect 62445 26429 62498 26710
rect 80526 26429 80579 26439
rect 62445 26428 80579 26429
rect 62445 26376 80526 26428
rect 80578 26376 80579 26428
rect 80526 26366 80579 26376
rect 93160 26232 93224 26246
rect 92936 26178 93164 26232
rect 92583 25609 92647 25623
rect 92583 25553 92587 25609
rect 92643 25553 92647 25609
rect 92583 25539 92647 25553
rect 92936 25482 92990 26178
rect 93160 26176 93164 26178
rect 93220 26176 93224 26232
rect 93160 26162 93224 26176
rect 93725 25547 93789 25561
rect 93076 25495 93729 25547
rect 93725 25491 93729 25495
rect 93785 25491 93789 25547
rect 93725 25477 93789 25491
rect 92118 25361 92182 25375
rect 92118 25305 92122 25361
rect 92178 25305 92182 25361
rect 92118 25291 92182 25305
rect 97194 25199 97275 25213
rect 97194 25177 97208 25199
rect 97260 25177 97275 25199
rect 79683 25119 79736 25129
rect 75902 25118 79736 25119
rect 75902 25066 79683 25118
rect 79735 25066 79736 25118
rect 79683 25056 79736 25066
rect 95669 25115 95739 25130
rect 95669 25059 95676 25115
rect 95732 25059 95739 25115
rect 95669 25053 95678 25059
rect 95730 25053 95739 25059
rect 95669 25041 95739 25053
rect 95669 25035 95678 25041
rect 95730 25035 95739 25041
rect 95669 24979 95676 25035
rect 95732 24979 95739 25035
rect 97194 25121 97206 25177
rect 97262 25121 97275 25177
rect 97194 25097 97208 25121
rect 97260 25097 97275 25121
rect 97194 25041 97206 25097
rect 97262 25041 97275 25097
rect 97194 25019 97208 25041
rect 97260 25019 97275 25041
rect 97194 25005 97275 25019
rect 93395 24957 93626 24973
rect 95669 24964 95739 24979
rect 93395 24901 93402 24957
rect 93458 24955 93482 24957
rect 93538 24955 93562 24957
rect 93472 24903 93482 24955
rect 93538 24903 93548 24955
rect 93458 24901 93482 24903
rect 93538 24901 93562 24903
rect 93618 24901 93626 24957
rect 93395 24886 93626 24901
rect 83095 24738 83170 24748
rect 90824 24743 90899 24748
rect 90824 24738 90904 24743
rect 83095 24726 90904 24738
rect 83095 24674 83106 24726
rect 83158 24674 90835 24726
rect 90887 24674 90904 24726
rect 83095 24663 90904 24674
rect 83095 24653 83170 24663
rect 90824 24659 90904 24663
rect 90824 24653 90899 24659
rect 95662 24641 95743 24655
rect 95662 24619 95676 24641
rect 95728 24619 95743 24641
rect 95662 24563 95674 24619
rect 95730 24563 95743 24619
rect 95662 24539 95676 24563
rect 95728 24539 95743 24563
rect 95662 24483 95674 24539
rect 95730 24483 95743 24539
rect 95662 24461 95676 24483
rect 95728 24461 95743 24483
rect 95662 24447 95743 24461
rect 97181 24654 97262 24668
rect 97181 24632 97195 24654
rect 97247 24632 97262 24654
rect 97181 24576 97193 24632
rect 97249 24576 97262 24632
rect 97181 24552 97195 24576
rect 97247 24552 97262 24576
rect 97181 24496 97193 24552
rect 97249 24496 97262 24552
rect 97181 24474 97195 24496
rect 97247 24474 97262 24496
rect 97181 24460 97262 24474
rect 93456 24416 93625 24429
rect 93456 24360 93472 24416
rect 93528 24414 93552 24416
rect 93534 24362 93546 24414
rect 93528 24360 93552 24362
rect 93608 24360 93625 24416
rect 93456 24347 93625 24360
rect 92122 24301 92186 24315
rect 57416 24239 78201 24264
rect 57416 24103 57420 24239
rect 78196 24103 78201 24239
rect 92122 24245 92126 24301
rect 92182 24245 92186 24301
rect 92122 24231 92186 24245
rect 99693 24304 103024 24341
rect 99693 24302 99730 24304
rect 99786 24302 99810 24304
rect 99866 24302 99890 24304
rect 99946 24302 99970 24304
rect 100026 24302 100050 24304
rect 100106 24302 100130 24304
rect 100186 24302 100210 24304
rect 100266 24302 100290 24304
rect 100346 24302 100370 24304
rect 100426 24302 100450 24304
rect 100506 24302 100530 24304
rect 100586 24302 100610 24304
rect 100666 24302 100690 24304
rect 100746 24302 100770 24304
rect 100826 24302 100850 24304
rect 100906 24302 100930 24304
rect 100986 24302 101010 24304
rect 101066 24302 101090 24304
rect 101146 24302 101170 24304
rect 101226 24302 101250 24304
rect 101306 24302 101330 24304
rect 101386 24302 101410 24304
rect 101466 24302 101490 24304
rect 101546 24302 101570 24304
rect 101626 24302 101650 24304
rect 101706 24302 101730 24304
rect 101786 24302 101810 24304
rect 101866 24302 101890 24304
rect 101946 24302 101970 24304
rect 102026 24302 102050 24304
rect 102106 24302 102130 24304
rect 102186 24302 102210 24304
rect 102266 24302 102290 24304
rect 102346 24302 102370 24304
rect 102426 24302 102450 24304
rect 102506 24302 102530 24304
rect 102586 24302 102610 24304
rect 102666 24302 102690 24304
rect 102746 24302 102770 24304
rect 102826 24302 102850 24304
rect 102906 24302 102930 24304
rect 102986 24302 103024 24304
rect 99693 24250 99700 24302
rect 99880 24250 99890 24302
rect 99946 24250 99956 24302
rect 100200 24250 100210 24302
rect 100266 24250 100276 24302
rect 100520 24250 100530 24302
rect 100586 24250 100596 24302
rect 100840 24250 100850 24302
rect 100906 24250 100916 24302
rect 101160 24250 101170 24302
rect 101226 24250 101236 24302
rect 101480 24250 101490 24302
rect 101546 24250 101556 24302
rect 101800 24250 101810 24302
rect 101866 24250 101876 24302
rect 102120 24250 102130 24302
rect 102186 24250 102196 24302
rect 102440 24250 102450 24302
rect 102506 24250 102516 24302
rect 102760 24250 102770 24302
rect 102826 24250 102836 24302
rect 103016 24250 103024 24302
rect 99693 24248 99730 24250
rect 99786 24248 99810 24250
rect 99866 24248 99890 24250
rect 99946 24248 99970 24250
rect 100026 24248 100050 24250
rect 100106 24248 100130 24250
rect 100186 24248 100210 24250
rect 100266 24248 100290 24250
rect 100346 24248 100370 24250
rect 100426 24248 100450 24250
rect 100506 24248 100530 24250
rect 100586 24248 100610 24250
rect 100666 24248 100690 24250
rect 100746 24248 100770 24250
rect 100826 24248 100850 24250
rect 100906 24248 100930 24250
rect 100986 24248 101010 24250
rect 101066 24248 101090 24250
rect 101146 24248 101170 24250
rect 101226 24248 101250 24250
rect 101306 24248 101330 24250
rect 101386 24248 101410 24250
rect 101466 24248 101490 24250
rect 101546 24248 101570 24250
rect 101626 24248 101650 24250
rect 101706 24248 101730 24250
rect 101786 24248 101810 24250
rect 101866 24248 101890 24250
rect 101946 24248 101970 24250
rect 102026 24248 102050 24250
rect 102106 24248 102130 24250
rect 102186 24248 102210 24250
rect 102266 24248 102290 24250
rect 102346 24248 102370 24250
rect 102426 24248 102450 24250
rect 102506 24248 102530 24250
rect 102586 24248 102610 24250
rect 102666 24248 102690 24250
rect 102746 24248 102770 24250
rect 102826 24248 102850 24250
rect 102906 24248 102930 24250
rect 102986 24248 103024 24250
rect 99693 24211 103024 24248
rect 57416 24079 78201 24103
rect 92121 24032 92185 24046
rect 92121 23976 92125 24032
rect 92181 23976 92185 24032
rect 92121 23962 92185 23976
rect 93446 23868 93531 23887
rect 93446 23812 93460 23868
rect 93516 23812 93531 23868
rect 93446 23793 93531 23812
rect 97186 23863 97267 23877
rect 97186 23841 97200 23863
rect 97252 23841 97267 23863
rect 95665 23784 95743 23799
rect 95665 23754 95678 23784
rect 95730 23754 95743 23784
rect 95665 23698 95676 23754
rect 95732 23698 95743 23754
rect 95665 23668 95678 23698
rect 95730 23668 95743 23698
rect 97186 23785 97198 23841
rect 97254 23785 97267 23841
rect 97186 23761 97200 23785
rect 97252 23761 97267 23785
rect 97186 23705 97198 23761
rect 97254 23705 97267 23761
rect 97186 23683 97200 23705
rect 97252 23683 97267 23705
rect 97186 23669 97267 23683
rect 95665 23654 95743 23668
rect 90828 23394 90892 23404
rect 80511 23387 90892 23394
rect 80511 23381 90835 23387
rect 80511 23329 80526 23381
rect 80578 23335 90835 23381
rect 90887 23335 90892 23387
rect 80578 23329 90892 23335
rect 80526 23319 80579 23329
rect 90828 23320 90892 23329
rect 94065 23327 94161 23357
rect 90835 23319 90888 23320
rect 94065 23271 94085 23327
rect 94141 23271 94161 23327
rect 94065 23241 94161 23271
rect 95657 23310 95738 23324
rect 95657 23288 95671 23310
rect 95723 23288 95738 23310
rect 95657 23232 95669 23288
rect 95725 23232 95738 23288
rect 95657 23208 95671 23232
rect 95723 23208 95738 23232
rect 95657 23152 95669 23208
rect 95725 23152 95738 23208
rect 95657 23130 95671 23152
rect 95723 23130 95738 23152
rect 95657 23116 95738 23130
rect 97186 23307 97267 23321
rect 97186 23285 97200 23307
rect 97252 23285 97267 23307
rect 97186 23229 97198 23285
rect 97254 23229 97267 23285
rect 97186 23205 97200 23229
rect 97252 23205 97267 23229
rect 97186 23149 97198 23205
rect 97254 23149 97267 23205
rect 97186 23127 97200 23149
rect 97252 23127 97267 23149
rect 97186 23113 97267 23127
rect 92121 22963 92185 22977
rect 92121 22907 92125 22963
rect 92181 22907 92185 22963
rect 92121 22893 92185 22907
rect 104583 22872 104819 22892
rect 93064 22785 93243 22799
rect 93064 22729 93085 22785
rect 93141 22783 93165 22785
rect 93147 22731 93159 22783
rect 93141 22729 93165 22731
rect 93221 22729 93243 22785
rect 93064 22716 93243 22729
rect 104583 22656 104593 22872
rect 104809 22656 104819 22872
rect 92118 22640 92182 22654
rect 92118 22584 92122 22640
rect 92178 22584 92182 22640
rect 104583 22636 104819 22656
rect 92118 22570 92182 22584
rect 97203 22483 97284 22497
rect 97203 22461 97217 22483
rect 97269 22461 97284 22483
rect 95668 22394 95742 22414
rect 95668 22364 95679 22394
rect 95731 22364 95742 22394
rect 95668 22308 95677 22364
rect 95733 22308 95742 22364
rect 95668 22278 95679 22308
rect 95731 22278 95742 22308
rect 97203 22405 97215 22461
rect 97271 22405 97284 22461
rect 97203 22381 97217 22405
rect 97269 22381 97284 22405
rect 97203 22325 97215 22381
rect 97271 22325 97284 22381
rect 97203 22303 97217 22325
rect 97269 22303 97284 22325
rect 97203 22289 97284 22303
rect 95668 22259 95742 22278
rect 93608 22237 93828 22254
rect 93608 22181 93610 22237
rect 93666 22235 93690 22237
rect 93746 22235 93770 22237
rect 93680 22183 93690 22235
rect 93746 22183 93756 22235
rect 93666 22181 93690 22183
rect 93746 22181 93770 22183
rect 93826 22181 93828 22237
rect 93608 22164 93828 22181
rect 79683 22005 79737 22015
rect 90840 22005 90900 22015
rect 79681 22004 90900 22005
rect 79681 21952 79684 22004
rect 79736 22001 90900 22004
rect 79736 21952 90844 22001
rect 79681 21949 90844 21952
rect 90896 21949 90900 22001
rect 79681 21945 90900 21949
rect 79683 21942 79737 21945
rect 90840 21935 90900 21945
rect 95656 21957 95737 21971
rect 95656 21935 95670 21957
rect 95722 21935 95737 21957
rect 95656 21879 95668 21935
rect 95724 21879 95737 21935
rect 95656 21855 95670 21879
rect 95722 21855 95737 21879
rect 95656 21799 95668 21855
rect 95724 21799 95737 21855
rect 95656 21777 95670 21799
rect 95722 21777 95737 21799
rect 95656 21763 95737 21777
rect 97186 21935 97267 21949
rect 97186 21913 97200 21935
rect 97252 21913 97267 21935
rect 97186 21857 97198 21913
rect 97254 21857 97267 21913
rect 97186 21833 97200 21857
rect 97252 21833 97267 21857
rect 97186 21777 97198 21833
rect 97254 21777 97267 21833
rect 97186 21755 97200 21777
rect 97252 21755 97267 21777
rect 97186 21741 97267 21755
rect 93458 21694 93603 21705
rect 93458 21638 93462 21694
rect 93518 21692 93542 21694
rect 93524 21640 93536 21692
rect 93518 21638 93542 21640
rect 93598 21638 93603 21694
rect 93458 21627 93603 21638
rect 92129 21570 92193 21584
rect 92129 21514 92133 21570
rect 92189 21514 92193 21570
rect 92129 21500 92193 21514
rect 99681 21298 103027 21324
rect 92118 21265 92182 21279
rect 92118 21209 92122 21265
rect 92178 21209 92182 21265
rect 99681 21242 99686 21298
rect 99742 21296 99766 21298
rect 99822 21296 99846 21298
rect 99902 21296 99926 21298
rect 99982 21296 100006 21298
rect 100062 21296 100086 21298
rect 100142 21296 100166 21298
rect 100222 21296 100246 21298
rect 100302 21296 100326 21298
rect 100382 21296 100406 21298
rect 100462 21296 100486 21298
rect 100542 21296 100566 21298
rect 100622 21296 100646 21298
rect 100702 21296 100726 21298
rect 100782 21296 100806 21298
rect 100862 21296 100886 21298
rect 100942 21296 100966 21298
rect 101022 21296 101046 21298
rect 101102 21296 101126 21298
rect 101182 21296 101206 21298
rect 101262 21296 101286 21298
rect 101342 21296 101366 21298
rect 101422 21296 101446 21298
rect 101502 21296 101526 21298
rect 101582 21296 101606 21298
rect 101662 21296 101686 21298
rect 101742 21296 101766 21298
rect 101822 21296 101846 21298
rect 101902 21296 101926 21298
rect 101982 21296 102006 21298
rect 102062 21296 102086 21298
rect 102142 21296 102166 21298
rect 102222 21296 102246 21298
rect 102302 21296 102326 21298
rect 102382 21296 102406 21298
rect 102462 21296 102486 21298
rect 102542 21296 102566 21298
rect 102622 21296 102646 21298
rect 102702 21296 102726 21298
rect 102782 21296 102806 21298
rect 102862 21296 102886 21298
rect 102942 21296 102966 21298
rect 99748 21244 99760 21296
rect 99822 21244 99824 21296
rect 100004 21244 100006 21296
rect 100068 21244 100080 21296
rect 100142 21244 100144 21296
rect 100324 21244 100326 21296
rect 100388 21244 100400 21296
rect 100462 21244 100464 21296
rect 100644 21244 100646 21296
rect 100708 21244 100720 21296
rect 100782 21244 100784 21296
rect 100964 21244 100966 21296
rect 101028 21244 101040 21296
rect 101102 21244 101104 21296
rect 101284 21244 101286 21296
rect 101348 21244 101360 21296
rect 101422 21244 101424 21296
rect 101604 21244 101606 21296
rect 101668 21244 101680 21296
rect 101742 21244 101744 21296
rect 101924 21244 101926 21296
rect 101988 21244 102000 21296
rect 102062 21244 102064 21296
rect 102244 21244 102246 21296
rect 102308 21244 102320 21296
rect 102382 21244 102384 21296
rect 102564 21244 102566 21296
rect 102628 21244 102640 21296
rect 102702 21244 102704 21296
rect 102884 21244 102886 21296
rect 102948 21244 102960 21296
rect 99742 21242 99766 21244
rect 99822 21242 99846 21244
rect 99902 21242 99926 21244
rect 99982 21242 100006 21244
rect 100062 21242 100086 21244
rect 100142 21242 100166 21244
rect 100222 21242 100246 21244
rect 100302 21242 100326 21244
rect 100382 21242 100406 21244
rect 100462 21242 100486 21244
rect 100542 21242 100566 21244
rect 100622 21242 100646 21244
rect 100702 21242 100726 21244
rect 100782 21242 100806 21244
rect 100862 21242 100886 21244
rect 100942 21242 100966 21244
rect 101022 21242 101046 21244
rect 101102 21242 101126 21244
rect 101182 21242 101206 21244
rect 101262 21242 101286 21244
rect 101342 21242 101366 21244
rect 101422 21242 101446 21244
rect 101502 21242 101526 21244
rect 101582 21242 101606 21244
rect 101662 21242 101686 21244
rect 101742 21242 101766 21244
rect 101822 21242 101846 21244
rect 101902 21242 101926 21244
rect 101982 21242 102006 21244
rect 102062 21242 102086 21244
rect 102142 21242 102166 21244
rect 102222 21242 102246 21244
rect 102302 21242 102326 21244
rect 102382 21242 102406 21244
rect 102462 21242 102486 21244
rect 102542 21242 102566 21244
rect 102622 21242 102646 21244
rect 102702 21242 102726 21244
rect 102782 21242 102806 21244
rect 102862 21242 102886 21244
rect 102942 21242 102966 21244
rect 103022 21242 103027 21298
rect 99681 21216 103027 21242
rect 92118 21195 92182 21209
rect 94066 21151 94162 21181
rect 94066 21095 94086 21151
rect 94142 21095 94162 21151
rect 94066 21065 94162 21095
rect 97193 21104 97274 21118
rect 97193 21082 97207 21104
rect 97259 21082 97274 21104
rect 97193 21026 97205 21082
rect 97261 21026 97274 21082
rect 95666 21007 95745 21026
rect 95666 20951 95677 21007
rect 95733 20951 95745 21007
rect 95666 20945 95679 20951
rect 95731 20945 95745 20951
rect 95666 20933 95745 20945
rect 95666 20927 95679 20933
rect 95731 20927 95745 20933
rect 95666 20871 95677 20927
rect 95733 20871 95745 20927
rect 97193 21002 97207 21026
rect 97259 21002 97274 21026
rect 97193 20946 97205 21002
rect 97261 20946 97274 21002
rect 97193 20924 97207 20946
rect 97259 20924 97274 20946
rect 97193 20910 97274 20924
rect 95666 20853 95745 20871
rect 93453 20605 93580 20623
rect 93453 20603 93488 20605
rect 93544 20603 93580 20605
rect 93453 20551 93458 20603
rect 93574 20551 93580 20603
rect 93453 20549 93488 20551
rect 93544 20549 93580 20551
rect 93453 20531 93580 20549
rect 95659 20557 95740 20571
rect 95659 20535 95673 20557
rect 95725 20535 95740 20557
rect 95659 20479 95671 20535
rect 95727 20479 95740 20535
rect 95659 20455 95673 20479
rect 95725 20455 95740 20479
rect 95659 20399 95671 20455
rect 95727 20399 95740 20455
rect 95659 20377 95673 20399
rect 95725 20377 95740 20399
rect 95659 20363 95740 20377
rect 97183 20551 97264 20565
rect 97183 20529 97197 20551
rect 97249 20529 97264 20551
rect 97183 20473 97195 20529
rect 97251 20473 97264 20529
rect 97183 20449 97197 20473
rect 97249 20449 97264 20473
rect 97183 20393 97195 20449
rect 97251 20393 97264 20449
rect 97183 20371 97197 20393
rect 97249 20371 97264 20393
rect 97183 20357 97264 20371
rect 92125 20200 92189 20214
rect 92125 20144 92129 20200
rect 92185 20144 92189 20200
rect 92125 20130 92189 20144
rect 53499 17174 53591 17210
rect 53499 17118 53517 17174
rect 53573 17118 53591 17174
rect 53499 17108 53591 17118
rect 53499 17094 53519 17108
rect 53571 17094 53591 17108
rect 53499 17038 53517 17094
rect 53573 17038 53591 17094
rect 53499 17014 53519 17038
rect 53571 17014 53591 17038
rect 53499 16958 53517 17014
rect 53573 16958 53591 17014
rect 53499 16934 53519 16958
rect 53571 16934 53591 16958
rect 53499 16878 53517 16934
rect 53573 16878 53591 16934
rect 53499 16864 53519 16878
rect 53571 16864 53591 16878
rect 53499 16854 53591 16864
rect 53499 16798 53517 16854
rect 53573 16798 53591 16854
rect 53499 16788 53591 16798
rect 53499 16774 53519 16788
rect 53571 16774 53591 16788
rect 53499 16718 53517 16774
rect 53573 16718 53591 16774
rect 53499 16694 53519 16718
rect 53571 16694 53591 16718
rect 53499 16638 53517 16694
rect 53573 16638 53591 16694
rect 53499 16614 53519 16638
rect 53571 16614 53591 16638
rect 53499 16558 53517 16614
rect 53573 16558 53591 16614
rect 53499 16544 53519 16558
rect 53571 16544 53591 16558
rect 53499 16534 53591 16544
rect 53499 16478 53517 16534
rect 53573 16478 53591 16534
rect 53499 16468 53591 16478
rect 53499 16454 53519 16468
rect 53571 16454 53591 16468
rect 53499 16398 53517 16454
rect 53573 16398 53591 16454
rect 53499 16374 53519 16398
rect 53571 16374 53591 16398
rect 53499 16318 53517 16374
rect 53573 16318 53591 16374
rect 53499 16294 53519 16318
rect 53571 16294 53591 16318
rect 53499 16238 53517 16294
rect 53573 16238 53591 16294
rect 53499 16224 53519 16238
rect 53571 16224 53591 16238
rect 53499 16214 53591 16224
rect 53499 16158 53517 16214
rect 53573 16158 53591 16214
rect 53499 16148 53591 16158
rect 53499 16134 53519 16148
rect 53571 16134 53591 16148
rect 53499 16078 53517 16134
rect 53573 16078 53591 16134
rect 53499 16054 53519 16078
rect 53571 16054 53591 16078
rect 53499 15998 53517 16054
rect 53573 15998 53591 16054
rect 53499 15974 53519 15998
rect 53571 15974 53591 15998
rect 53499 15918 53517 15974
rect 53573 15918 53591 15974
rect 53499 15904 53519 15918
rect 53571 15904 53591 15918
rect 53499 15894 53591 15904
rect 53499 15838 53517 15894
rect 53573 15838 53591 15894
rect 53499 15828 53591 15838
rect 53499 15814 53519 15828
rect 53571 15814 53591 15828
rect 53499 15758 53517 15814
rect 53573 15758 53591 15814
rect 53499 15734 53519 15758
rect 53571 15734 53591 15758
rect 53499 15678 53517 15734
rect 53573 15678 53591 15734
rect 53499 15654 53519 15678
rect 53571 15654 53591 15678
rect 53499 15598 53517 15654
rect 53573 15598 53591 15654
rect 53499 15584 53519 15598
rect 53571 15584 53591 15598
rect 53499 15574 53591 15584
rect 53499 15518 53517 15574
rect 53573 15518 53591 15574
rect 53499 15508 53591 15518
rect 53499 15494 53519 15508
rect 53571 15494 53591 15508
rect 53499 15438 53517 15494
rect 53573 15438 53591 15494
rect 53499 15414 53519 15438
rect 53571 15414 53591 15438
rect 53499 15358 53517 15414
rect 53573 15358 53591 15414
rect 53499 15334 53519 15358
rect 53571 15334 53591 15358
rect 53499 15278 53517 15334
rect 53573 15278 53591 15334
rect 53499 15264 53519 15278
rect 53571 15264 53591 15278
rect 53499 15254 53591 15264
rect 53499 15198 53517 15254
rect 53573 15198 53591 15254
rect 53499 15188 53591 15198
rect 53499 15174 53519 15188
rect 53571 15174 53591 15188
rect 53499 15118 53517 15174
rect 53573 15118 53591 15174
rect 53499 15094 53519 15118
rect 53571 15094 53591 15118
rect 53499 15038 53517 15094
rect 53573 15038 53591 15094
rect 53499 15014 53519 15038
rect 53571 15014 53591 15038
rect 53499 14958 53517 15014
rect 53573 14958 53591 15014
rect 53499 14944 53519 14958
rect 53571 14944 53591 14958
rect 53499 14934 53591 14944
rect 53499 14878 53517 14934
rect 53573 14878 53591 14934
rect 53499 14868 53591 14878
rect 53499 14854 53519 14868
rect 53571 14854 53591 14868
rect 53499 14798 53517 14854
rect 53573 14798 53591 14854
rect 53499 14774 53519 14798
rect 53571 14774 53591 14798
rect 53499 14718 53517 14774
rect 53573 14718 53591 14774
rect 53499 14694 53519 14718
rect 53571 14694 53591 14718
rect 53499 14638 53517 14694
rect 53573 14638 53591 14694
rect 53499 14624 53519 14638
rect 53571 14624 53591 14638
rect 53499 14614 53591 14624
rect 53499 14558 53517 14614
rect 53573 14558 53591 14614
rect 53499 14548 53591 14558
rect 53499 14534 53519 14548
rect 53571 14534 53591 14548
rect 53499 14478 53517 14534
rect 53573 14478 53591 14534
rect 53499 14454 53519 14478
rect 53571 14454 53591 14478
rect 53499 14398 53517 14454
rect 53573 14398 53591 14454
rect 53499 14374 53519 14398
rect 53571 14374 53591 14398
rect 53499 14318 53517 14374
rect 53573 14318 53591 14374
rect 53499 14304 53519 14318
rect 53571 14304 53591 14318
rect 53499 14294 53591 14304
rect 53499 14238 53517 14294
rect 53573 14238 53591 14294
rect 53499 14228 53591 14238
rect 53499 14214 53519 14228
rect 53571 14214 53591 14228
rect 53499 14158 53517 14214
rect 53573 14158 53591 14214
rect 53499 14134 53519 14158
rect 53571 14134 53591 14158
rect 53499 14078 53517 14134
rect 53573 14078 53591 14134
rect 53499 14054 53519 14078
rect 53571 14054 53591 14078
rect 53499 13998 53517 14054
rect 53573 13998 53591 14054
rect 53499 13984 53519 13998
rect 53571 13984 53591 13998
rect 53499 13974 53591 13984
rect 53499 13918 53517 13974
rect 53573 13918 53591 13974
rect 53499 13882 53591 13918
rect 56494 17167 56608 17207
rect 56494 17111 56523 17167
rect 56579 17111 56608 17167
rect 56494 17101 56608 17111
rect 56494 17087 56525 17101
rect 56577 17087 56608 17101
rect 56494 17031 56523 17087
rect 56579 17031 56608 17087
rect 56494 17007 56525 17031
rect 56577 17007 56608 17031
rect 56494 16951 56523 17007
rect 56579 16951 56608 17007
rect 56494 16927 56525 16951
rect 56577 16927 56608 16951
rect 56494 16871 56523 16927
rect 56579 16871 56608 16927
rect 56494 16857 56525 16871
rect 56577 16857 56608 16871
rect 56494 16847 56608 16857
rect 56494 16791 56523 16847
rect 56579 16791 56608 16847
rect 56494 16781 56608 16791
rect 56494 16767 56525 16781
rect 56577 16767 56608 16781
rect 56494 16711 56523 16767
rect 56579 16711 56608 16767
rect 56494 16687 56525 16711
rect 56577 16687 56608 16711
rect 56494 16631 56523 16687
rect 56579 16631 56608 16687
rect 56494 16607 56525 16631
rect 56577 16607 56608 16631
rect 56494 16551 56523 16607
rect 56579 16551 56608 16607
rect 56494 16537 56525 16551
rect 56577 16537 56608 16551
rect 56494 16527 56608 16537
rect 56494 16471 56523 16527
rect 56579 16471 56608 16527
rect 56494 16461 56608 16471
rect 56494 16447 56525 16461
rect 56577 16447 56608 16461
rect 56494 16391 56523 16447
rect 56579 16391 56608 16447
rect 56494 16367 56525 16391
rect 56577 16367 56608 16391
rect 56494 16311 56523 16367
rect 56579 16311 56608 16367
rect 56494 16287 56525 16311
rect 56577 16287 56608 16311
rect 56494 16231 56523 16287
rect 56579 16231 56608 16287
rect 56494 16217 56525 16231
rect 56577 16217 56608 16231
rect 56494 16207 56608 16217
rect 56494 16151 56523 16207
rect 56579 16151 56608 16207
rect 56494 16141 56608 16151
rect 56494 16127 56525 16141
rect 56577 16127 56608 16141
rect 56494 16071 56523 16127
rect 56579 16071 56608 16127
rect 56494 16047 56525 16071
rect 56577 16047 56608 16071
rect 56494 15991 56523 16047
rect 56579 15991 56608 16047
rect 56494 15967 56525 15991
rect 56577 15967 56608 15991
rect 56494 15911 56523 15967
rect 56579 15911 56608 15967
rect 56494 15897 56525 15911
rect 56577 15897 56608 15911
rect 56494 15887 56608 15897
rect 56494 15831 56523 15887
rect 56579 15831 56608 15887
rect 56494 15821 56608 15831
rect 56494 15807 56525 15821
rect 56577 15807 56608 15821
rect 56494 15751 56523 15807
rect 56579 15751 56608 15807
rect 56494 15727 56525 15751
rect 56577 15727 56608 15751
rect 56494 15671 56523 15727
rect 56579 15671 56608 15727
rect 56494 15647 56525 15671
rect 56577 15647 56608 15671
rect 56494 15591 56523 15647
rect 56579 15591 56608 15647
rect 56494 15577 56525 15591
rect 56577 15577 56608 15591
rect 56494 15567 56608 15577
rect 56494 15511 56523 15567
rect 56579 15511 56608 15567
rect 56494 15501 56608 15511
rect 56494 15487 56525 15501
rect 56577 15487 56608 15501
rect 56494 15431 56523 15487
rect 56579 15431 56608 15487
rect 56494 15407 56525 15431
rect 56577 15407 56608 15431
rect 56494 15351 56523 15407
rect 56579 15351 56608 15407
rect 56494 15327 56525 15351
rect 56577 15327 56608 15351
rect 56494 15271 56523 15327
rect 56579 15271 56608 15327
rect 56494 15257 56525 15271
rect 56577 15257 56608 15271
rect 56494 15247 56608 15257
rect 56494 15191 56523 15247
rect 56579 15191 56608 15247
rect 56494 15181 56608 15191
rect 56494 15167 56525 15181
rect 56577 15167 56608 15181
rect 56494 15111 56523 15167
rect 56579 15111 56608 15167
rect 56494 15087 56525 15111
rect 56577 15087 56608 15111
rect 56494 15031 56523 15087
rect 56579 15031 56608 15087
rect 56494 15007 56525 15031
rect 56577 15007 56608 15031
rect 56494 14951 56523 15007
rect 56579 14951 56608 15007
rect 56494 14937 56525 14951
rect 56577 14937 56608 14951
rect 56494 14927 56608 14937
rect 56494 14871 56523 14927
rect 56579 14871 56608 14927
rect 56494 14861 56608 14871
rect 56494 14847 56525 14861
rect 56577 14847 56608 14861
rect 56494 14791 56523 14847
rect 56579 14791 56608 14847
rect 56494 14767 56525 14791
rect 56577 14767 56608 14791
rect 56494 14711 56523 14767
rect 56579 14711 56608 14767
rect 56494 14687 56525 14711
rect 56577 14687 56608 14711
rect 56494 14631 56523 14687
rect 56579 14631 56608 14687
rect 56494 14617 56525 14631
rect 56577 14617 56608 14631
rect 56494 14607 56608 14617
rect 56494 14551 56523 14607
rect 56579 14551 56608 14607
rect 56494 14541 56608 14551
rect 56494 14527 56525 14541
rect 56577 14527 56608 14541
rect 56494 14471 56523 14527
rect 56579 14471 56608 14527
rect 56494 14447 56525 14471
rect 56577 14447 56608 14471
rect 56494 14391 56523 14447
rect 56579 14391 56608 14447
rect 56494 14367 56525 14391
rect 56577 14367 56608 14391
rect 56494 14311 56523 14367
rect 56579 14311 56608 14367
rect 56494 14297 56525 14311
rect 56577 14297 56608 14311
rect 56494 14287 56608 14297
rect 56494 14231 56523 14287
rect 56579 14231 56608 14287
rect 56494 14221 56608 14231
rect 56494 14207 56525 14221
rect 56577 14207 56608 14221
rect 56494 14151 56523 14207
rect 56579 14151 56608 14207
rect 56494 14127 56525 14151
rect 56577 14127 56608 14151
rect 56494 14071 56523 14127
rect 56579 14071 56608 14127
rect 56494 14047 56525 14071
rect 56577 14047 56608 14071
rect 56494 13991 56523 14047
rect 56579 13991 56608 14047
rect 56494 13977 56525 13991
rect 56577 13977 56608 13991
rect 56494 13967 56608 13977
rect 56494 13911 56523 13967
rect 56579 13911 56608 13967
rect 56494 13872 56608 13911
rect 54915 11930 55151 11950
rect 54915 11714 54925 11930
rect 55141 11714 55151 11930
rect 54915 11694 55151 11714
<< via2 >>
rect 41694 102134 41910 102152
rect 41694 101954 41712 102134
rect 41712 101954 41892 102134
rect 41892 101954 41910 102134
rect 41694 101936 41910 101954
rect 69710 102105 69926 102123
rect 69710 101925 69728 102105
rect 69728 101925 69908 102105
rect 69908 101925 69926 102105
rect 69710 101907 69926 101925
rect 81760 102106 81976 102124
rect 81760 101926 81778 102106
rect 81778 101926 81958 102106
rect 81958 101926 81976 102106
rect 81760 101908 81976 101926
rect 40267 100688 40269 100710
rect 40269 100688 40321 100710
rect 40321 100688 40323 100710
rect 40267 100676 40323 100688
rect 40267 100654 40269 100676
rect 40269 100654 40321 100676
rect 40321 100654 40323 100676
rect 40267 100624 40269 100630
rect 40269 100624 40321 100630
rect 40321 100624 40323 100630
rect 40267 100612 40323 100624
rect 40267 100574 40269 100612
rect 40269 100574 40321 100612
rect 40321 100574 40323 100612
rect 40267 100548 40323 100550
rect 40267 100496 40269 100548
rect 40269 100496 40321 100548
rect 40321 100496 40323 100548
rect 40267 100494 40323 100496
rect 40267 100432 40269 100470
rect 40269 100432 40321 100470
rect 40321 100432 40323 100470
rect 40267 100420 40323 100432
rect 40267 100414 40269 100420
rect 40269 100414 40321 100420
rect 40321 100414 40323 100420
rect 40267 100368 40269 100390
rect 40269 100368 40321 100390
rect 40321 100368 40323 100390
rect 40267 100356 40323 100368
rect 40267 100334 40269 100356
rect 40269 100334 40321 100356
rect 40321 100334 40323 100356
rect 40267 100304 40269 100310
rect 40269 100304 40321 100310
rect 40321 100304 40323 100310
rect 40267 100292 40323 100304
rect 40267 100254 40269 100292
rect 40269 100254 40321 100292
rect 40321 100254 40323 100292
rect 40267 100228 40323 100230
rect 40267 100176 40269 100228
rect 40269 100176 40321 100228
rect 40321 100176 40323 100228
rect 40267 100174 40323 100176
rect 40267 100112 40269 100150
rect 40269 100112 40321 100150
rect 40321 100112 40323 100150
rect 40267 100100 40323 100112
rect 40267 100094 40269 100100
rect 40269 100094 40321 100100
rect 40321 100094 40323 100100
rect 40267 100048 40269 100070
rect 40269 100048 40321 100070
rect 40321 100048 40323 100070
rect 40267 100036 40323 100048
rect 40267 100014 40269 100036
rect 40269 100014 40321 100036
rect 40321 100014 40323 100036
rect 40267 99984 40269 99990
rect 40269 99984 40321 99990
rect 40321 99984 40323 99990
rect 40267 99972 40323 99984
rect 40267 99934 40269 99972
rect 40269 99934 40321 99972
rect 40321 99934 40323 99972
rect 40267 99908 40323 99910
rect 40267 99856 40269 99908
rect 40269 99856 40321 99908
rect 40321 99856 40323 99908
rect 40267 99854 40323 99856
rect 40267 99792 40269 99830
rect 40269 99792 40321 99830
rect 40321 99792 40323 99830
rect 40267 99780 40323 99792
rect 40267 99774 40269 99780
rect 40269 99774 40321 99780
rect 40321 99774 40323 99780
rect 40267 99728 40269 99750
rect 40269 99728 40321 99750
rect 40321 99728 40323 99750
rect 40267 99716 40323 99728
rect 40267 99694 40269 99716
rect 40269 99694 40321 99716
rect 40321 99694 40323 99716
rect 40267 99664 40269 99670
rect 40269 99664 40321 99670
rect 40321 99664 40323 99670
rect 40267 99652 40323 99664
rect 40267 99614 40269 99652
rect 40269 99614 40321 99652
rect 40321 99614 40323 99652
rect 40267 99588 40323 99590
rect 40267 99536 40269 99588
rect 40269 99536 40321 99588
rect 40321 99536 40323 99588
rect 40267 99534 40323 99536
rect 40267 99472 40269 99510
rect 40269 99472 40321 99510
rect 40321 99472 40323 99510
rect 40267 99460 40323 99472
rect 40267 99454 40269 99460
rect 40269 99454 40321 99460
rect 40321 99454 40323 99460
rect 40267 99408 40269 99430
rect 40269 99408 40321 99430
rect 40321 99408 40323 99430
rect 40267 99396 40323 99408
rect 40267 99374 40269 99396
rect 40269 99374 40321 99396
rect 40321 99374 40323 99396
rect 40267 99344 40269 99350
rect 40269 99344 40321 99350
rect 40321 99344 40323 99350
rect 40267 99332 40323 99344
rect 40267 99294 40269 99332
rect 40269 99294 40321 99332
rect 40321 99294 40323 99332
rect 40267 99268 40323 99270
rect 40267 99216 40269 99268
rect 40269 99216 40321 99268
rect 40321 99216 40323 99268
rect 40267 99214 40323 99216
rect 40267 99152 40269 99190
rect 40269 99152 40321 99190
rect 40321 99152 40323 99190
rect 40267 99140 40323 99152
rect 40267 99134 40269 99140
rect 40269 99134 40321 99140
rect 40321 99134 40323 99140
rect 40267 99088 40269 99110
rect 40269 99088 40321 99110
rect 40321 99088 40323 99110
rect 40267 99076 40323 99088
rect 40267 99054 40269 99076
rect 40269 99054 40321 99076
rect 40321 99054 40323 99076
rect 40267 99024 40269 99030
rect 40269 99024 40321 99030
rect 40321 99024 40323 99030
rect 40267 99012 40323 99024
rect 40267 98974 40269 99012
rect 40269 98974 40321 99012
rect 40321 98974 40323 99012
rect 40267 98948 40323 98950
rect 40267 98896 40269 98948
rect 40269 98896 40321 98948
rect 40321 98896 40323 98948
rect 40267 98894 40323 98896
rect 40267 98832 40269 98870
rect 40269 98832 40321 98870
rect 40321 98832 40323 98870
rect 40267 98820 40323 98832
rect 40267 98814 40269 98820
rect 40269 98814 40321 98820
rect 40321 98814 40323 98820
rect 40267 98768 40269 98790
rect 40269 98768 40321 98790
rect 40321 98768 40323 98790
rect 40267 98756 40323 98768
rect 40267 98734 40269 98756
rect 40269 98734 40321 98756
rect 40321 98734 40323 98756
rect 40267 98704 40269 98710
rect 40269 98704 40321 98710
rect 40321 98704 40323 98710
rect 40267 98692 40323 98704
rect 40267 98654 40269 98692
rect 40269 98654 40321 98692
rect 40321 98654 40323 98692
rect 40267 98628 40323 98630
rect 40267 98576 40269 98628
rect 40269 98576 40321 98628
rect 40321 98576 40323 98628
rect 40267 98574 40323 98576
rect 40267 98512 40269 98550
rect 40269 98512 40321 98550
rect 40321 98512 40323 98550
rect 40267 98500 40323 98512
rect 40267 98494 40269 98500
rect 40269 98494 40321 98500
rect 40321 98494 40323 98500
rect 40267 98448 40269 98470
rect 40269 98448 40321 98470
rect 40321 98448 40323 98470
rect 40267 98436 40323 98448
rect 40267 98414 40269 98436
rect 40269 98414 40321 98436
rect 40321 98414 40323 98436
rect 40267 98384 40269 98390
rect 40269 98384 40321 98390
rect 40321 98384 40323 98390
rect 40267 98372 40323 98384
rect 40267 98334 40269 98372
rect 40269 98334 40321 98372
rect 40321 98334 40323 98372
rect 40267 98308 40323 98310
rect 40267 98256 40269 98308
rect 40269 98256 40321 98308
rect 40321 98256 40323 98308
rect 40267 98254 40323 98256
rect 40267 98192 40269 98230
rect 40269 98192 40321 98230
rect 40321 98192 40323 98230
rect 40267 98180 40323 98192
rect 40267 98174 40269 98180
rect 40269 98174 40321 98180
rect 40321 98174 40323 98180
rect 40267 98128 40269 98150
rect 40269 98128 40321 98150
rect 40321 98128 40323 98150
rect 40267 98116 40323 98128
rect 40267 98094 40269 98116
rect 40269 98094 40321 98116
rect 40321 98094 40323 98116
rect 40267 98064 40269 98070
rect 40269 98064 40321 98070
rect 40321 98064 40323 98070
rect 40267 98052 40323 98064
rect 40267 98014 40269 98052
rect 40269 98014 40321 98052
rect 40321 98014 40323 98052
rect 40267 97988 40323 97990
rect 40267 97936 40269 97988
rect 40269 97936 40321 97988
rect 40321 97936 40323 97988
rect 40267 97934 40323 97936
rect 40267 97872 40269 97910
rect 40269 97872 40321 97910
rect 40321 97872 40323 97910
rect 40267 97860 40323 97872
rect 40267 97854 40269 97860
rect 40269 97854 40321 97860
rect 40321 97854 40323 97860
rect 40267 97808 40269 97830
rect 40269 97808 40321 97830
rect 40321 97808 40323 97830
rect 40267 97796 40323 97808
rect 40267 97774 40269 97796
rect 40269 97774 40321 97796
rect 40321 97774 40323 97796
rect 40267 97744 40269 97750
rect 40269 97744 40321 97750
rect 40321 97744 40323 97750
rect 40267 97732 40323 97744
rect 40267 97694 40269 97732
rect 40269 97694 40321 97732
rect 40321 97694 40323 97732
rect 40267 97668 40323 97670
rect 40267 97616 40269 97668
rect 40269 97616 40321 97668
rect 40321 97616 40323 97668
rect 40267 97614 40323 97616
rect 40267 97552 40269 97590
rect 40269 97552 40321 97590
rect 40321 97552 40323 97590
rect 40267 97540 40323 97552
rect 40267 97534 40269 97540
rect 40269 97534 40321 97540
rect 40321 97534 40323 97540
rect 40267 97488 40269 97510
rect 40269 97488 40321 97510
rect 40321 97488 40323 97510
rect 40267 97476 40323 97488
rect 40267 97454 40269 97476
rect 40269 97454 40321 97476
rect 40321 97454 40323 97476
rect 43268 100694 43270 100716
rect 43270 100694 43322 100716
rect 43322 100694 43324 100716
rect 43268 100682 43324 100694
rect 43268 100660 43270 100682
rect 43270 100660 43322 100682
rect 43322 100660 43324 100682
rect 43268 100630 43270 100636
rect 43270 100630 43322 100636
rect 43322 100630 43324 100636
rect 43268 100618 43324 100630
rect 43268 100580 43270 100618
rect 43270 100580 43322 100618
rect 43322 100580 43324 100618
rect 43268 100554 43324 100556
rect 43268 100502 43270 100554
rect 43270 100502 43322 100554
rect 43322 100502 43324 100554
rect 43268 100500 43324 100502
rect 43268 100438 43270 100476
rect 43270 100438 43322 100476
rect 43322 100438 43324 100476
rect 43268 100426 43324 100438
rect 43268 100420 43270 100426
rect 43270 100420 43322 100426
rect 43322 100420 43324 100426
rect 43268 100374 43270 100396
rect 43270 100374 43322 100396
rect 43322 100374 43324 100396
rect 43268 100362 43324 100374
rect 43268 100340 43270 100362
rect 43270 100340 43322 100362
rect 43322 100340 43324 100362
rect 43268 100310 43270 100316
rect 43270 100310 43322 100316
rect 43322 100310 43324 100316
rect 43268 100298 43324 100310
rect 43268 100260 43270 100298
rect 43270 100260 43322 100298
rect 43322 100260 43324 100298
rect 43268 100234 43324 100236
rect 43268 100182 43270 100234
rect 43270 100182 43322 100234
rect 43322 100182 43324 100234
rect 43268 100180 43324 100182
rect 43268 100118 43270 100156
rect 43270 100118 43322 100156
rect 43322 100118 43324 100156
rect 43268 100106 43324 100118
rect 43268 100100 43270 100106
rect 43270 100100 43322 100106
rect 43322 100100 43324 100106
rect 43268 100054 43270 100076
rect 43270 100054 43322 100076
rect 43322 100054 43324 100076
rect 43268 100042 43324 100054
rect 43268 100020 43270 100042
rect 43270 100020 43322 100042
rect 43322 100020 43324 100042
rect 43268 99990 43270 99996
rect 43270 99990 43322 99996
rect 43322 99990 43324 99996
rect 43268 99978 43324 99990
rect 43268 99940 43270 99978
rect 43270 99940 43322 99978
rect 43322 99940 43324 99978
rect 43268 99914 43324 99916
rect 43268 99862 43270 99914
rect 43270 99862 43322 99914
rect 43322 99862 43324 99914
rect 43268 99860 43324 99862
rect 43268 99798 43270 99836
rect 43270 99798 43322 99836
rect 43322 99798 43324 99836
rect 43268 99786 43324 99798
rect 43268 99780 43270 99786
rect 43270 99780 43322 99786
rect 43322 99780 43324 99786
rect 43268 99734 43270 99756
rect 43270 99734 43322 99756
rect 43322 99734 43324 99756
rect 43268 99722 43324 99734
rect 43268 99700 43270 99722
rect 43270 99700 43322 99722
rect 43322 99700 43324 99722
rect 43268 99670 43270 99676
rect 43270 99670 43322 99676
rect 43322 99670 43324 99676
rect 43268 99658 43324 99670
rect 43268 99620 43270 99658
rect 43270 99620 43322 99658
rect 43322 99620 43324 99658
rect 43268 99594 43324 99596
rect 43268 99542 43270 99594
rect 43270 99542 43322 99594
rect 43322 99542 43324 99594
rect 43268 99540 43324 99542
rect 43268 99478 43270 99516
rect 43270 99478 43322 99516
rect 43322 99478 43324 99516
rect 43268 99466 43324 99478
rect 43268 99460 43270 99466
rect 43270 99460 43322 99466
rect 43322 99460 43324 99466
rect 43268 99414 43270 99436
rect 43270 99414 43322 99436
rect 43322 99414 43324 99436
rect 43268 99402 43324 99414
rect 43268 99380 43270 99402
rect 43270 99380 43322 99402
rect 43322 99380 43324 99402
rect 43268 99350 43270 99356
rect 43270 99350 43322 99356
rect 43322 99350 43324 99356
rect 43268 99338 43324 99350
rect 43268 99300 43270 99338
rect 43270 99300 43322 99338
rect 43322 99300 43324 99338
rect 43268 99274 43324 99276
rect 43268 99222 43270 99274
rect 43270 99222 43322 99274
rect 43322 99222 43324 99274
rect 43268 99220 43324 99222
rect 43268 99158 43270 99196
rect 43270 99158 43322 99196
rect 43322 99158 43324 99196
rect 43268 99146 43324 99158
rect 43268 99140 43270 99146
rect 43270 99140 43322 99146
rect 43322 99140 43324 99146
rect 43268 99094 43270 99116
rect 43270 99094 43322 99116
rect 43322 99094 43324 99116
rect 43268 99082 43324 99094
rect 43268 99060 43270 99082
rect 43270 99060 43322 99082
rect 43322 99060 43324 99082
rect 43268 99030 43270 99036
rect 43270 99030 43322 99036
rect 43322 99030 43324 99036
rect 43268 99018 43324 99030
rect 43268 98980 43270 99018
rect 43270 98980 43322 99018
rect 43322 98980 43324 99018
rect 43268 98954 43324 98956
rect 43268 98902 43270 98954
rect 43270 98902 43322 98954
rect 43322 98902 43324 98954
rect 43268 98900 43324 98902
rect 43268 98838 43270 98876
rect 43270 98838 43322 98876
rect 43322 98838 43324 98876
rect 43268 98826 43324 98838
rect 43268 98820 43270 98826
rect 43270 98820 43322 98826
rect 43322 98820 43324 98826
rect 43268 98774 43270 98796
rect 43270 98774 43322 98796
rect 43322 98774 43324 98796
rect 43268 98762 43324 98774
rect 43268 98740 43270 98762
rect 43270 98740 43322 98762
rect 43322 98740 43324 98762
rect 43268 98710 43270 98716
rect 43270 98710 43322 98716
rect 43322 98710 43324 98716
rect 43268 98698 43324 98710
rect 43268 98660 43270 98698
rect 43270 98660 43322 98698
rect 43322 98660 43324 98698
rect 43268 98634 43324 98636
rect 43268 98582 43270 98634
rect 43270 98582 43322 98634
rect 43322 98582 43324 98634
rect 43268 98580 43324 98582
rect 43268 98518 43270 98556
rect 43270 98518 43322 98556
rect 43322 98518 43324 98556
rect 43268 98506 43324 98518
rect 43268 98500 43270 98506
rect 43270 98500 43322 98506
rect 43322 98500 43324 98506
rect 43268 98454 43270 98476
rect 43270 98454 43322 98476
rect 43322 98454 43324 98476
rect 43268 98442 43324 98454
rect 43268 98420 43270 98442
rect 43270 98420 43322 98442
rect 43322 98420 43324 98442
rect 43268 98390 43270 98396
rect 43270 98390 43322 98396
rect 43322 98390 43324 98396
rect 43268 98378 43324 98390
rect 43268 98340 43270 98378
rect 43270 98340 43322 98378
rect 43322 98340 43324 98378
rect 43268 98314 43324 98316
rect 43268 98262 43270 98314
rect 43270 98262 43322 98314
rect 43322 98262 43324 98314
rect 43268 98260 43324 98262
rect 43268 98198 43270 98236
rect 43270 98198 43322 98236
rect 43322 98198 43324 98236
rect 43268 98186 43324 98198
rect 43268 98180 43270 98186
rect 43270 98180 43322 98186
rect 43322 98180 43324 98186
rect 43268 98134 43270 98156
rect 43270 98134 43322 98156
rect 43322 98134 43324 98156
rect 43268 98122 43324 98134
rect 43268 98100 43270 98122
rect 43270 98100 43322 98122
rect 43322 98100 43324 98122
rect 43268 98070 43270 98076
rect 43270 98070 43322 98076
rect 43322 98070 43324 98076
rect 43268 98058 43324 98070
rect 43268 98020 43270 98058
rect 43270 98020 43322 98058
rect 43322 98020 43324 98058
rect 43268 97994 43324 97996
rect 43268 97942 43270 97994
rect 43270 97942 43322 97994
rect 43322 97942 43324 97994
rect 43268 97940 43324 97942
rect 43268 97878 43270 97916
rect 43270 97878 43322 97916
rect 43322 97878 43324 97916
rect 43268 97866 43324 97878
rect 43268 97860 43270 97866
rect 43270 97860 43322 97866
rect 43322 97860 43324 97866
rect 43268 97814 43270 97836
rect 43270 97814 43322 97836
rect 43322 97814 43324 97836
rect 43268 97802 43324 97814
rect 43268 97780 43270 97802
rect 43270 97780 43322 97802
rect 43322 97780 43324 97802
rect 43268 97750 43270 97756
rect 43270 97750 43322 97756
rect 43322 97750 43324 97756
rect 43268 97738 43324 97750
rect 43268 97700 43270 97738
rect 43270 97700 43322 97738
rect 43322 97700 43324 97738
rect 43268 97674 43324 97676
rect 43268 97622 43270 97674
rect 43270 97622 43322 97674
rect 43322 97622 43324 97674
rect 43268 97620 43324 97622
rect 43268 97558 43270 97596
rect 43270 97558 43322 97596
rect 43322 97558 43324 97596
rect 43268 97546 43324 97558
rect 43268 97540 43270 97546
rect 43270 97540 43322 97546
rect 43322 97540 43324 97546
rect 43268 97494 43270 97516
rect 43270 97494 43322 97516
rect 43322 97494 43324 97516
rect 43268 97482 43324 97494
rect 43268 97460 43270 97482
rect 43270 97460 43322 97482
rect 43322 97460 43324 97482
rect 68273 100742 68329 100752
rect 68273 100696 68329 100742
rect 68273 100616 68329 100672
rect 68273 100536 68329 100592
rect 68273 100456 68329 100512
rect 68273 100376 68329 100432
rect 68273 100296 68329 100352
rect 68273 100216 68329 100272
rect 68273 100136 68329 100192
rect 68273 100056 68329 100112
rect 68273 99976 68329 100032
rect 68273 99896 68329 99952
rect 68273 99816 68329 99872
rect 68273 99736 68329 99792
rect 68273 99656 68329 99712
rect 68273 99576 68329 99632
rect 68273 99496 68329 99552
rect 68273 99416 68329 99472
rect 68273 99336 68329 99392
rect 68273 99256 68329 99312
rect 68273 99176 68329 99232
rect 68273 99096 68329 99152
rect 68273 99016 68329 99072
rect 68273 98936 68329 98992
rect 68273 98856 68329 98912
rect 68273 98776 68329 98832
rect 68273 98696 68329 98752
rect 68273 98616 68329 98672
rect 68273 98536 68329 98592
rect 68273 98456 68329 98512
rect 68273 98376 68329 98432
rect 68273 98296 68329 98352
rect 68273 98216 68329 98272
rect 68273 98136 68329 98192
rect 68273 98056 68329 98112
rect 68273 97976 68329 98032
rect 68273 97896 68329 97952
rect 68273 97816 68329 97872
rect 68273 97736 68329 97792
rect 68273 97656 68329 97712
rect 68273 97576 68329 97632
rect 68273 97496 68329 97552
rect 68273 97426 68329 97472
rect 68273 97416 68329 97426
rect 71274 100755 71330 100765
rect 71274 100709 71330 100755
rect 71274 100629 71330 100685
rect 71274 100549 71330 100605
rect 71274 100469 71330 100525
rect 71274 100389 71330 100445
rect 71274 100309 71330 100365
rect 71274 100229 71330 100285
rect 71274 100149 71330 100205
rect 71274 100069 71330 100125
rect 71274 99989 71330 100045
rect 71274 99909 71330 99965
rect 71274 99829 71330 99885
rect 71274 99749 71330 99805
rect 71274 99669 71330 99725
rect 71274 99589 71330 99645
rect 71274 99509 71330 99565
rect 71274 99429 71330 99485
rect 71274 99349 71330 99405
rect 71274 99269 71330 99325
rect 71274 99189 71330 99245
rect 71274 99109 71330 99165
rect 71274 99029 71330 99085
rect 71274 98949 71330 99005
rect 71274 98869 71330 98925
rect 71274 98789 71330 98845
rect 71274 98709 71330 98765
rect 71274 98629 71330 98685
rect 71274 98549 71330 98605
rect 71274 98469 71330 98525
rect 71274 98389 71330 98445
rect 71274 98309 71330 98365
rect 71274 98229 71330 98285
rect 71274 98149 71330 98205
rect 71274 98069 71330 98125
rect 71274 97989 71330 98045
rect 71274 97909 71330 97965
rect 71274 97829 71330 97885
rect 71274 97749 71330 97805
rect 71274 97669 71330 97725
rect 71274 97589 71330 97645
rect 71274 97509 71330 97565
rect 71274 97439 71330 97485
rect 71274 97429 71330 97439
rect 40434 95818 40490 95820
rect 40434 95766 40436 95818
rect 40436 95766 40488 95818
rect 40488 95766 40490 95818
rect 40434 95764 40490 95766
rect 41612 95814 41668 95816
rect 41612 95762 41614 95814
rect 41614 95762 41666 95814
rect 41666 95762 41668 95814
rect 41612 95760 41668 95762
rect 41829 95821 41885 95823
rect 41829 95769 41831 95821
rect 41831 95769 41883 95821
rect 41883 95769 41885 95821
rect 41829 95767 41885 95769
rect 42963 95818 43019 95820
rect 42963 95766 42965 95818
rect 42965 95766 43017 95818
rect 43017 95766 43019 95818
rect 42963 95764 43019 95766
rect 40544 94314 40600 94316
rect 40544 94262 40546 94314
rect 40546 94262 40598 94314
rect 40598 94262 40600 94314
rect 40544 94260 40600 94262
rect 41658 94300 41714 94302
rect 41658 94248 41660 94300
rect 41660 94248 41712 94300
rect 41712 94248 41714 94300
rect 41658 94246 41714 94248
rect 41871 94301 41927 94303
rect 41871 94249 41873 94301
rect 41873 94249 41925 94301
rect 41925 94249 41927 94301
rect 41871 94247 41927 94249
rect 43035 94301 43091 94303
rect 43035 94249 43037 94301
rect 43037 94249 43089 94301
rect 43089 94249 43091 94301
rect 43035 94247 43091 94249
rect 40390 92665 40446 92721
rect 41676 92464 41678 92510
rect 41678 92464 41730 92510
rect 41730 92464 41732 92510
rect 41676 92454 41732 92464
rect 41676 92400 41678 92430
rect 41678 92400 41730 92430
rect 41730 92400 41732 92430
rect 41676 92388 41732 92400
rect 41676 92374 41678 92388
rect 41678 92374 41730 92388
rect 41730 92374 41732 92388
rect 41676 92336 41678 92350
rect 41678 92336 41730 92350
rect 41730 92336 41732 92350
rect 41676 92324 41732 92336
rect 41676 92294 41678 92324
rect 41678 92294 41730 92324
rect 41730 92294 41732 92324
rect 41139 92263 41195 92273
rect 41139 92217 41141 92263
rect 41141 92217 41193 92263
rect 41193 92217 41195 92263
rect 41139 92147 41141 92193
rect 41141 92147 41193 92193
rect 41193 92147 41195 92193
rect 41139 92137 41195 92147
rect 41676 92260 41732 92270
rect 41676 92214 41678 92260
rect 41678 92214 41730 92260
rect 41730 92214 41732 92260
rect 42223 92266 42279 92276
rect 42223 92220 42225 92266
rect 42225 92220 42277 92266
rect 42277 92220 42279 92266
rect 42223 92150 42225 92196
rect 42225 92150 42277 92196
rect 42277 92150 42279 92196
rect 42223 92140 42279 92150
rect 42899 92035 42955 92091
rect 40521 91629 40577 91631
rect 40521 91577 40523 91629
rect 40523 91577 40575 91629
rect 40575 91577 40577 91629
rect 40521 91575 40577 91577
rect 41676 91623 41732 91625
rect 41676 91571 41678 91623
rect 41678 91571 41730 91623
rect 41730 91571 41732 91623
rect 41676 91569 41732 91571
rect 42794 91634 42850 91636
rect 42794 91582 42796 91634
rect 42796 91582 42848 91634
rect 42848 91582 42850 91634
rect 42794 91580 42850 91582
rect 74529 88708 74531 88746
rect 74531 88708 74583 88746
rect 74583 88708 74585 88746
rect 74529 88696 74585 88708
rect 74529 88690 74531 88696
rect 74531 88690 74583 88696
rect 74583 88690 74585 88696
rect 74529 88644 74531 88666
rect 74531 88644 74583 88666
rect 74583 88644 74585 88666
rect 74529 88632 74585 88644
rect 74529 88610 74531 88632
rect 74531 88610 74583 88632
rect 74583 88610 74585 88632
rect 74529 88580 74531 88586
rect 74531 88580 74583 88586
rect 74583 88580 74585 88586
rect 74529 88568 74585 88580
rect 74529 88530 74531 88568
rect 74531 88530 74583 88568
rect 74583 88530 74585 88568
rect 74529 88504 74585 88506
rect 74529 88452 74531 88504
rect 74531 88452 74583 88504
rect 74583 88452 74585 88504
rect 74529 88450 74585 88452
rect 74529 88388 74531 88426
rect 74531 88388 74583 88426
rect 74583 88388 74585 88426
rect 74529 88376 74585 88388
rect 74529 88370 74531 88376
rect 74531 88370 74583 88376
rect 74583 88370 74585 88376
rect 74529 88324 74531 88346
rect 74531 88324 74583 88346
rect 74583 88324 74585 88346
rect 74529 88312 74585 88324
rect 74529 88290 74531 88312
rect 74531 88290 74583 88312
rect 74583 88290 74585 88312
rect 74529 88260 74531 88266
rect 74531 88260 74583 88266
rect 74583 88260 74585 88266
rect 74529 88248 74585 88260
rect 74529 88210 74531 88248
rect 74531 88210 74583 88248
rect 74583 88210 74585 88248
rect 81057 88708 81059 88746
rect 81059 88708 81111 88746
rect 81111 88708 81113 88746
rect 81057 88696 81113 88708
rect 81057 88690 81059 88696
rect 81059 88690 81111 88696
rect 81111 88690 81113 88696
rect 81057 88644 81059 88666
rect 81059 88644 81111 88666
rect 81111 88644 81113 88666
rect 81057 88632 81113 88644
rect 81057 88610 81059 88632
rect 81059 88610 81111 88632
rect 81111 88610 81113 88632
rect 81057 88580 81059 88586
rect 81059 88580 81111 88586
rect 81111 88580 81113 88586
rect 81057 88568 81113 88580
rect 81057 88530 81059 88568
rect 81059 88530 81111 88568
rect 81111 88530 81113 88568
rect 81057 88504 81113 88506
rect 81057 88452 81059 88504
rect 81059 88452 81111 88504
rect 81111 88452 81113 88504
rect 81057 88450 81113 88452
rect 81057 88388 81059 88426
rect 81059 88388 81111 88426
rect 81111 88388 81113 88426
rect 81057 88376 81113 88388
rect 81057 88370 81059 88376
rect 81059 88370 81111 88376
rect 81111 88370 81113 88376
rect 81057 88324 81059 88346
rect 81059 88324 81111 88346
rect 81111 88324 81113 88346
rect 81057 88312 81113 88324
rect 81057 88290 81059 88312
rect 81059 88290 81111 88312
rect 81111 88290 81113 88312
rect 81057 88260 81059 88266
rect 81059 88260 81111 88266
rect 81111 88260 81113 88266
rect 81057 88248 81113 88260
rect 81057 88210 81059 88248
rect 81059 88210 81111 88248
rect 81111 88210 81113 88248
rect 88673 88708 88675 88746
rect 88675 88708 88727 88746
rect 88727 88708 88729 88746
rect 88673 88696 88729 88708
rect 88673 88690 88675 88696
rect 88675 88690 88727 88696
rect 88727 88690 88729 88696
rect 88673 88644 88675 88666
rect 88675 88644 88727 88666
rect 88727 88644 88729 88666
rect 88673 88632 88729 88644
rect 88673 88610 88675 88632
rect 88675 88610 88727 88632
rect 88727 88610 88729 88632
rect 88673 88580 88675 88586
rect 88675 88580 88727 88586
rect 88727 88580 88729 88586
rect 88673 88568 88729 88580
rect 88673 88530 88675 88568
rect 88675 88530 88727 88568
rect 88727 88530 88729 88568
rect 88673 88504 88729 88506
rect 88673 88452 88675 88504
rect 88675 88452 88727 88504
rect 88727 88452 88729 88504
rect 88673 88450 88729 88452
rect 88673 88388 88675 88426
rect 88675 88388 88727 88426
rect 88727 88388 88729 88426
rect 88673 88376 88729 88388
rect 88673 88370 88675 88376
rect 88675 88370 88727 88376
rect 88727 88370 88729 88376
rect 88673 88324 88675 88346
rect 88675 88324 88727 88346
rect 88727 88324 88729 88346
rect 88673 88312 88729 88324
rect 88673 88290 88675 88312
rect 88675 88290 88727 88312
rect 88727 88290 88729 88312
rect 88673 88260 88675 88266
rect 88675 88260 88727 88266
rect 88727 88260 88729 88266
rect 88673 88248 88729 88260
rect 88673 88210 88675 88248
rect 88675 88210 88727 88248
rect 88727 88210 88729 88248
rect 47243 87418 47299 87420
rect 47323 87418 47379 87420
rect 47403 87418 47459 87420
rect 47483 87418 47539 87420
rect 47563 87418 47619 87420
rect 47243 87366 47265 87418
rect 47265 87366 47277 87418
rect 47277 87366 47299 87418
rect 47323 87366 47329 87418
rect 47329 87366 47341 87418
rect 47341 87366 47379 87418
rect 47403 87366 47405 87418
rect 47405 87366 47457 87418
rect 47457 87366 47459 87418
rect 47483 87366 47521 87418
rect 47521 87366 47533 87418
rect 47533 87366 47539 87418
rect 47563 87366 47585 87418
rect 47585 87366 47597 87418
rect 47597 87366 47619 87418
rect 47243 87364 47299 87366
rect 47323 87364 47379 87366
rect 47403 87364 47459 87366
rect 47483 87364 47539 87366
rect 47563 87364 47619 87366
rect 49054 87420 49110 87422
rect 49134 87420 49190 87422
rect 49214 87420 49270 87422
rect 49294 87420 49350 87422
rect 49374 87420 49430 87422
rect 49054 87368 49076 87420
rect 49076 87368 49088 87420
rect 49088 87368 49110 87420
rect 49134 87368 49140 87420
rect 49140 87368 49152 87420
rect 49152 87368 49190 87420
rect 49214 87368 49216 87420
rect 49216 87368 49268 87420
rect 49268 87368 49270 87420
rect 49294 87368 49332 87420
rect 49332 87368 49344 87420
rect 49344 87368 49350 87420
rect 49374 87368 49396 87420
rect 49396 87368 49408 87420
rect 49408 87368 49430 87420
rect 49054 87366 49110 87368
rect 49134 87366 49190 87368
rect 49214 87366 49270 87368
rect 49294 87366 49350 87368
rect 49374 87366 49430 87368
rect 50849 87416 50905 87418
rect 50929 87416 50985 87418
rect 51009 87416 51065 87418
rect 51089 87416 51145 87418
rect 51169 87416 51225 87418
rect 50849 87364 50871 87416
rect 50871 87364 50883 87416
rect 50883 87364 50905 87416
rect 50929 87364 50935 87416
rect 50935 87364 50947 87416
rect 50947 87364 50985 87416
rect 51009 87364 51011 87416
rect 51011 87364 51063 87416
rect 51063 87364 51065 87416
rect 51089 87364 51127 87416
rect 51127 87364 51139 87416
rect 51139 87364 51145 87416
rect 51169 87364 51191 87416
rect 51191 87364 51203 87416
rect 51203 87364 51225 87416
rect 50849 87362 50905 87364
rect 50929 87362 50985 87364
rect 51009 87362 51065 87364
rect 51089 87362 51145 87364
rect 51169 87362 51225 87364
rect 52648 87414 52704 87416
rect 52728 87414 52784 87416
rect 52808 87414 52864 87416
rect 52888 87414 52944 87416
rect 52968 87414 53024 87416
rect 52648 87362 52670 87414
rect 52670 87362 52682 87414
rect 52682 87362 52704 87414
rect 52728 87362 52734 87414
rect 52734 87362 52746 87414
rect 52746 87362 52784 87414
rect 52808 87362 52810 87414
rect 52810 87362 52862 87414
rect 52862 87362 52864 87414
rect 52888 87362 52926 87414
rect 52926 87362 52938 87414
rect 52938 87362 52944 87414
rect 52968 87362 52990 87414
rect 52990 87362 53002 87414
rect 53002 87362 53024 87414
rect 52648 87360 52704 87362
rect 52728 87360 52784 87362
rect 52808 87360 52864 87362
rect 52888 87360 52944 87362
rect 52968 87360 53024 87362
rect 54439 87418 54495 87420
rect 54519 87418 54575 87420
rect 54599 87418 54655 87420
rect 54679 87418 54735 87420
rect 54759 87418 54815 87420
rect 54439 87366 54461 87418
rect 54461 87366 54473 87418
rect 54473 87366 54495 87418
rect 54519 87366 54525 87418
rect 54525 87366 54537 87418
rect 54537 87366 54575 87418
rect 54599 87366 54601 87418
rect 54601 87366 54653 87418
rect 54653 87366 54655 87418
rect 54679 87366 54717 87418
rect 54717 87366 54729 87418
rect 54729 87366 54735 87418
rect 54759 87366 54781 87418
rect 54781 87366 54793 87418
rect 54793 87366 54815 87418
rect 54439 87364 54495 87366
rect 54519 87364 54575 87366
rect 54599 87364 54655 87366
rect 54679 87364 54735 87366
rect 54759 87364 54815 87366
rect 56241 87414 56297 87416
rect 56321 87414 56377 87416
rect 56401 87414 56457 87416
rect 56481 87414 56537 87416
rect 56561 87414 56617 87416
rect 56241 87362 56263 87414
rect 56263 87362 56275 87414
rect 56275 87362 56297 87414
rect 56321 87362 56327 87414
rect 56327 87362 56339 87414
rect 56339 87362 56377 87414
rect 56401 87362 56403 87414
rect 56403 87362 56455 87414
rect 56455 87362 56457 87414
rect 56481 87362 56519 87414
rect 56519 87362 56531 87414
rect 56531 87362 56537 87414
rect 56561 87362 56583 87414
rect 56583 87362 56595 87414
rect 56595 87362 56617 87414
rect 56241 87360 56297 87362
rect 56321 87360 56377 87362
rect 56401 87360 56457 87362
rect 56481 87360 56537 87362
rect 56561 87360 56617 87362
rect 50167 87198 50383 87216
rect 50167 87018 50185 87198
rect 50185 87018 50365 87198
rect 50365 87018 50383 87198
rect 50167 87000 50383 87018
rect 57888 87224 58344 87242
rect 57888 87044 58344 87224
rect 57888 87026 58344 87044
rect 75074 86705 75076 86743
rect 75076 86705 75128 86743
rect 75128 86705 75130 86743
rect 75074 86693 75130 86705
rect 75074 86687 75076 86693
rect 75076 86687 75128 86693
rect 75128 86687 75130 86693
rect 75074 86641 75076 86663
rect 75076 86641 75128 86663
rect 75128 86641 75130 86663
rect 75074 86629 75130 86641
rect 75074 86607 75076 86629
rect 75076 86607 75128 86629
rect 75128 86607 75130 86629
rect 75074 86577 75076 86583
rect 75076 86577 75128 86583
rect 75128 86577 75130 86583
rect 75074 86565 75130 86577
rect 75074 86527 75076 86565
rect 75076 86527 75128 86565
rect 75128 86527 75130 86565
rect 75074 86501 75130 86503
rect 75074 86449 75076 86501
rect 75076 86449 75128 86501
rect 75128 86449 75130 86501
rect 75074 86447 75130 86449
rect 75074 86385 75076 86423
rect 75076 86385 75128 86423
rect 75128 86385 75130 86423
rect 75074 86373 75130 86385
rect 75074 86367 75076 86373
rect 75076 86367 75128 86373
rect 75128 86367 75130 86373
rect 75074 86321 75076 86343
rect 75076 86321 75128 86343
rect 75128 86321 75130 86343
rect 75074 86309 75130 86321
rect 75074 86287 75076 86309
rect 75076 86287 75128 86309
rect 75128 86287 75130 86309
rect 75074 86257 75076 86263
rect 75076 86257 75128 86263
rect 75128 86257 75130 86263
rect 75074 86245 75130 86257
rect 75074 86207 75076 86245
rect 75076 86207 75128 86245
rect 75128 86207 75130 86245
rect 76162 86705 76164 86743
rect 76164 86705 76216 86743
rect 76216 86705 76218 86743
rect 76162 86693 76218 86705
rect 76162 86687 76164 86693
rect 76164 86687 76216 86693
rect 76216 86687 76218 86693
rect 76162 86641 76164 86663
rect 76164 86641 76216 86663
rect 76216 86641 76218 86663
rect 76162 86629 76218 86641
rect 76162 86607 76164 86629
rect 76164 86607 76216 86629
rect 76216 86607 76218 86629
rect 76162 86577 76164 86583
rect 76164 86577 76216 86583
rect 76216 86577 76218 86583
rect 76162 86565 76218 86577
rect 76162 86527 76164 86565
rect 76164 86527 76216 86565
rect 76216 86527 76218 86565
rect 76162 86501 76218 86503
rect 76162 86449 76164 86501
rect 76164 86449 76216 86501
rect 76216 86449 76218 86501
rect 76162 86447 76218 86449
rect 76162 86385 76164 86423
rect 76164 86385 76216 86423
rect 76216 86385 76218 86423
rect 76162 86373 76218 86385
rect 76162 86367 76164 86373
rect 76164 86367 76216 86373
rect 76216 86367 76218 86373
rect 76162 86321 76164 86343
rect 76164 86321 76216 86343
rect 76216 86321 76218 86343
rect 76162 86309 76218 86321
rect 76162 86287 76164 86309
rect 76164 86287 76216 86309
rect 76216 86287 76218 86309
rect 76162 86257 76164 86263
rect 76164 86257 76216 86263
rect 76216 86257 76218 86263
rect 76162 86245 76218 86257
rect 76162 86207 76164 86245
rect 76164 86207 76216 86245
rect 76216 86207 76218 86245
rect 78338 86705 78340 86743
rect 78340 86705 78392 86743
rect 78392 86705 78394 86743
rect 78338 86693 78394 86705
rect 78338 86687 78340 86693
rect 78340 86687 78392 86693
rect 78392 86687 78394 86693
rect 78338 86641 78340 86663
rect 78340 86641 78392 86663
rect 78392 86641 78394 86663
rect 78338 86629 78394 86641
rect 78338 86607 78340 86629
rect 78340 86607 78392 86629
rect 78392 86607 78394 86629
rect 78338 86577 78340 86583
rect 78340 86577 78392 86583
rect 78392 86577 78394 86583
rect 78338 86565 78394 86577
rect 78338 86527 78340 86565
rect 78340 86527 78392 86565
rect 78392 86527 78394 86565
rect 78338 86501 78394 86503
rect 78338 86449 78340 86501
rect 78340 86449 78392 86501
rect 78392 86449 78394 86501
rect 78338 86447 78394 86449
rect 78338 86385 78340 86423
rect 78340 86385 78392 86423
rect 78392 86385 78394 86423
rect 78338 86373 78394 86385
rect 78338 86367 78340 86373
rect 78340 86367 78392 86373
rect 78392 86367 78394 86373
rect 78338 86321 78340 86343
rect 78340 86321 78392 86343
rect 78392 86321 78394 86343
rect 78338 86309 78394 86321
rect 78338 86287 78340 86309
rect 78340 86287 78392 86309
rect 78392 86287 78394 86309
rect 78338 86257 78340 86263
rect 78340 86257 78392 86263
rect 78392 86257 78394 86263
rect 78338 86245 78394 86257
rect 78338 86207 78340 86245
rect 78340 86207 78392 86245
rect 78392 86207 78394 86245
rect 79426 86705 79428 86743
rect 79428 86705 79480 86743
rect 79480 86705 79482 86743
rect 79426 86693 79482 86705
rect 79426 86687 79428 86693
rect 79428 86687 79480 86693
rect 79480 86687 79482 86693
rect 79426 86641 79428 86663
rect 79428 86641 79480 86663
rect 79480 86641 79482 86663
rect 79426 86629 79482 86641
rect 79426 86607 79428 86629
rect 79428 86607 79480 86629
rect 79480 86607 79482 86629
rect 79426 86577 79428 86583
rect 79428 86577 79480 86583
rect 79480 86577 79482 86583
rect 79426 86565 79482 86577
rect 79426 86527 79428 86565
rect 79428 86527 79480 86565
rect 79480 86527 79482 86565
rect 79426 86501 79482 86503
rect 79426 86449 79428 86501
rect 79428 86449 79480 86501
rect 79480 86449 79482 86501
rect 79426 86447 79482 86449
rect 79426 86385 79428 86423
rect 79428 86385 79480 86423
rect 79480 86385 79482 86423
rect 79426 86373 79482 86385
rect 79426 86367 79428 86373
rect 79428 86367 79480 86373
rect 79480 86367 79482 86373
rect 79426 86321 79428 86343
rect 79428 86321 79480 86343
rect 79480 86321 79482 86343
rect 79426 86309 79482 86321
rect 79426 86287 79428 86309
rect 79428 86287 79480 86309
rect 79480 86287 79482 86309
rect 79426 86257 79428 86263
rect 79428 86257 79480 86263
rect 79480 86257 79482 86263
rect 79426 86245 79482 86257
rect 79426 86207 79428 86245
rect 79428 86207 79480 86245
rect 79480 86207 79482 86245
rect 80514 86705 80516 86743
rect 80516 86705 80568 86743
rect 80568 86705 80570 86743
rect 80514 86693 80570 86705
rect 80514 86687 80516 86693
rect 80516 86687 80568 86693
rect 80568 86687 80570 86693
rect 80514 86641 80516 86663
rect 80516 86641 80568 86663
rect 80568 86641 80570 86663
rect 80514 86629 80570 86641
rect 80514 86607 80516 86629
rect 80516 86607 80568 86629
rect 80568 86607 80570 86629
rect 80514 86577 80516 86583
rect 80516 86577 80568 86583
rect 80568 86577 80570 86583
rect 80514 86565 80570 86577
rect 80514 86527 80516 86565
rect 80516 86527 80568 86565
rect 80568 86527 80570 86565
rect 80514 86501 80570 86503
rect 80514 86449 80516 86501
rect 80516 86449 80568 86501
rect 80568 86449 80570 86501
rect 80514 86447 80570 86449
rect 80514 86385 80516 86423
rect 80516 86385 80568 86423
rect 80568 86385 80570 86423
rect 80514 86373 80570 86385
rect 80514 86367 80516 86373
rect 80516 86367 80568 86373
rect 80568 86367 80570 86373
rect 80514 86321 80516 86343
rect 80516 86321 80568 86343
rect 80568 86321 80570 86343
rect 80514 86309 80570 86321
rect 80514 86287 80516 86309
rect 80516 86287 80568 86309
rect 80568 86287 80570 86309
rect 80514 86257 80516 86263
rect 80516 86257 80568 86263
rect 80568 86257 80570 86263
rect 80514 86245 80570 86257
rect 80514 86207 80516 86245
rect 80516 86207 80568 86245
rect 80568 86207 80570 86245
rect 81602 86705 81604 86743
rect 81604 86705 81656 86743
rect 81656 86705 81658 86743
rect 81602 86693 81658 86705
rect 81602 86687 81604 86693
rect 81604 86687 81656 86693
rect 81656 86687 81658 86693
rect 81602 86641 81604 86663
rect 81604 86641 81656 86663
rect 81656 86641 81658 86663
rect 81602 86629 81658 86641
rect 81602 86607 81604 86629
rect 81604 86607 81656 86629
rect 81656 86607 81658 86629
rect 81602 86577 81604 86583
rect 81604 86577 81656 86583
rect 81656 86577 81658 86583
rect 81602 86565 81658 86577
rect 81602 86527 81604 86565
rect 81604 86527 81656 86565
rect 81656 86527 81658 86565
rect 81602 86501 81658 86503
rect 81602 86449 81604 86501
rect 81604 86449 81656 86501
rect 81656 86449 81658 86501
rect 81602 86447 81658 86449
rect 81602 86385 81604 86423
rect 81604 86385 81656 86423
rect 81656 86385 81658 86423
rect 81602 86373 81658 86385
rect 81602 86367 81604 86373
rect 81604 86367 81656 86373
rect 81656 86367 81658 86373
rect 81602 86321 81604 86343
rect 81604 86321 81656 86343
rect 81656 86321 81658 86343
rect 81602 86309 81658 86321
rect 81602 86287 81604 86309
rect 81604 86287 81656 86309
rect 81656 86287 81658 86309
rect 81602 86257 81604 86263
rect 81604 86257 81656 86263
rect 81656 86257 81658 86263
rect 81602 86245 81658 86257
rect 81602 86207 81604 86245
rect 81604 86207 81656 86245
rect 81656 86207 81658 86245
rect 82690 86705 82692 86743
rect 82692 86705 82744 86743
rect 82744 86705 82746 86743
rect 82690 86693 82746 86705
rect 82690 86687 82692 86693
rect 82692 86687 82744 86693
rect 82744 86687 82746 86693
rect 82690 86641 82692 86663
rect 82692 86641 82744 86663
rect 82744 86641 82746 86663
rect 82690 86629 82746 86641
rect 82690 86607 82692 86629
rect 82692 86607 82744 86629
rect 82744 86607 82746 86629
rect 82690 86577 82692 86583
rect 82692 86577 82744 86583
rect 82744 86577 82746 86583
rect 82690 86565 82746 86577
rect 82690 86527 82692 86565
rect 82692 86527 82744 86565
rect 82744 86527 82746 86565
rect 82690 86501 82746 86503
rect 82690 86449 82692 86501
rect 82692 86449 82744 86501
rect 82744 86449 82746 86501
rect 82690 86447 82746 86449
rect 82690 86385 82692 86423
rect 82692 86385 82744 86423
rect 82744 86385 82746 86423
rect 82690 86373 82746 86385
rect 82690 86367 82692 86373
rect 82692 86367 82744 86373
rect 82744 86367 82746 86373
rect 82690 86321 82692 86343
rect 82692 86321 82744 86343
rect 82744 86321 82746 86343
rect 82690 86309 82746 86321
rect 82690 86287 82692 86309
rect 82692 86287 82744 86309
rect 82744 86287 82746 86309
rect 82690 86257 82692 86263
rect 82692 86257 82744 86263
rect 82744 86257 82746 86263
rect 82690 86245 82746 86257
rect 82690 86207 82692 86245
rect 82692 86207 82744 86245
rect 82744 86207 82746 86245
rect 83778 86705 83780 86743
rect 83780 86705 83832 86743
rect 83832 86705 83834 86743
rect 83778 86693 83834 86705
rect 83778 86687 83780 86693
rect 83780 86687 83832 86693
rect 83832 86687 83834 86693
rect 83778 86641 83780 86663
rect 83780 86641 83832 86663
rect 83832 86641 83834 86663
rect 83778 86629 83834 86641
rect 83778 86607 83780 86629
rect 83780 86607 83832 86629
rect 83832 86607 83834 86629
rect 83778 86577 83780 86583
rect 83780 86577 83832 86583
rect 83832 86577 83834 86583
rect 83778 86565 83834 86577
rect 83778 86527 83780 86565
rect 83780 86527 83832 86565
rect 83832 86527 83834 86565
rect 83778 86501 83834 86503
rect 83778 86449 83780 86501
rect 83780 86449 83832 86501
rect 83832 86449 83834 86501
rect 83778 86447 83834 86449
rect 83778 86385 83780 86423
rect 83780 86385 83832 86423
rect 83832 86385 83834 86423
rect 83778 86373 83834 86385
rect 83778 86367 83780 86373
rect 83780 86367 83832 86373
rect 83832 86367 83834 86373
rect 83778 86321 83780 86343
rect 83780 86321 83832 86343
rect 83832 86321 83834 86343
rect 83778 86309 83834 86321
rect 83778 86287 83780 86309
rect 83780 86287 83832 86309
rect 83832 86287 83834 86309
rect 83778 86257 83780 86263
rect 83780 86257 83832 86263
rect 83832 86257 83834 86263
rect 83778 86245 83834 86257
rect 83778 86207 83780 86245
rect 83780 86207 83832 86245
rect 83832 86207 83834 86245
rect 85954 86705 85956 86743
rect 85956 86705 86008 86743
rect 86008 86705 86010 86743
rect 85954 86693 86010 86705
rect 85954 86687 85956 86693
rect 85956 86687 86008 86693
rect 86008 86687 86010 86693
rect 85954 86641 85956 86663
rect 85956 86641 86008 86663
rect 86008 86641 86010 86663
rect 85954 86629 86010 86641
rect 85954 86607 85956 86629
rect 85956 86607 86008 86629
rect 86008 86607 86010 86629
rect 85954 86577 85956 86583
rect 85956 86577 86008 86583
rect 86008 86577 86010 86583
rect 85954 86565 86010 86577
rect 85954 86527 85956 86565
rect 85956 86527 86008 86565
rect 86008 86527 86010 86565
rect 85954 86501 86010 86503
rect 85954 86449 85956 86501
rect 85956 86449 86008 86501
rect 86008 86449 86010 86501
rect 85954 86447 86010 86449
rect 85954 86385 85956 86423
rect 85956 86385 86008 86423
rect 86008 86385 86010 86423
rect 85954 86373 86010 86385
rect 85954 86367 85956 86373
rect 85956 86367 86008 86373
rect 86008 86367 86010 86373
rect 85954 86321 85956 86343
rect 85956 86321 86008 86343
rect 86008 86321 86010 86343
rect 85954 86309 86010 86321
rect 85954 86287 85956 86309
rect 85956 86287 86008 86309
rect 86008 86287 86010 86309
rect 85954 86257 85956 86263
rect 85956 86257 86008 86263
rect 86008 86257 86010 86263
rect 85954 86245 86010 86257
rect 85954 86207 85956 86245
rect 85956 86207 86008 86245
rect 86008 86207 86010 86245
rect 87042 86705 87044 86743
rect 87044 86705 87096 86743
rect 87096 86705 87098 86743
rect 87042 86693 87098 86705
rect 87042 86687 87044 86693
rect 87044 86687 87096 86693
rect 87096 86687 87098 86693
rect 87042 86641 87044 86663
rect 87044 86641 87096 86663
rect 87096 86641 87098 86663
rect 87042 86629 87098 86641
rect 87042 86607 87044 86629
rect 87044 86607 87096 86629
rect 87096 86607 87098 86629
rect 87042 86577 87044 86583
rect 87044 86577 87096 86583
rect 87096 86577 87098 86583
rect 87042 86565 87098 86577
rect 87042 86527 87044 86565
rect 87044 86527 87096 86565
rect 87096 86527 87098 86565
rect 87042 86501 87098 86503
rect 87042 86449 87044 86501
rect 87044 86449 87096 86501
rect 87096 86449 87098 86501
rect 87042 86447 87098 86449
rect 87042 86385 87044 86423
rect 87044 86385 87096 86423
rect 87096 86385 87098 86423
rect 87042 86373 87098 86385
rect 87042 86367 87044 86373
rect 87044 86367 87096 86373
rect 87096 86367 87098 86373
rect 87042 86321 87044 86343
rect 87044 86321 87096 86343
rect 87096 86321 87098 86343
rect 87042 86309 87098 86321
rect 87042 86287 87044 86309
rect 87044 86287 87096 86309
rect 87096 86287 87098 86309
rect 87042 86257 87044 86263
rect 87044 86257 87096 86263
rect 87096 86257 87098 86263
rect 87042 86245 87098 86257
rect 87042 86207 87044 86245
rect 87044 86207 87096 86245
rect 87096 86207 87098 86245
rect 88130 86705 88132 86743
rect 88132 86705 88184 86743
rect 88184 86705 88186 86743
rect 88130 86693 88186 86705
rect 88130 86687 88132 86693
rect 88132 86687 88184 86693
rect 88184 86687 88186 86693
rect 88130 86641 88132 86663
rect 88132 86641 88184 86663
rect 88184 86641 88186 86663
rect 88130 86629 88186 86641
rect 88130 86607 88132 86629
rect 88132 86607 88184 86629
rect 88184 86607 88186 86629
rect 88130 86577 88132 86583
rect 88132 86577 88184 86583
rect 88184 86577 88186 86583
rect 88130 86565 88186 86577
rect 88130 86527 88132 86565
rect 88132 86527 88184 86565
rect 88184 86527 88186 86565
rect 88130 86501 88186 86503
rect 88130 86449 88132 86501
rect 88132 86449 88184 86501
rect 88184 86449 88186 86501
rect 88130 86447 88186 86449
rect 88130 86385 88132 86423
rect 88132 86385 88184 86423
rect 88184 86385 88186 86423
rect 88130 86373 88186 86385
rect 88130 86367 88132 86373
rect 88132 86367 88184 86373
rect 88184 86367 88186 86373
rect 88130 86321 88132 86343
rect 88132 86321 88184 86343
rect 88184 86321 88186 86343
rect 88130 86309 88186 86321
rect 88130 86287 88132 86309
rect 88132 86287 88184 86309
rect 88184 86287 88186 86309
rect 88130 86257 88132 86263
rect 88132 86257 88184 86263
rect 88184 86257 88186 86263
rect 88130 86245 88186 86257
rect 88130 86207 88132 86245
rect 88132 86207 88184 86245
rect 88184 86207 88186 86245
rect 48541 78611 48597 78613
rect 48541 78559 48543 78611
rect 48543 78559 48595 78611
rect 48595 78559 48597 78611
rect 48541 78557 48597 78559
rect 50232 78612 50288 78614
rect 50232 78560 50234 78612
rect 50234 78560 50286 78612
rect 50286 78560 50288 78612
rect 50232 78558 50288 78560
rect 51937 78611 51993 78613
rect 51937 78559 51939 78611
rect 51939 78559 51991 78611
rect 51991 78559 51993 78611
rect 51937 78557 51993 78559
rect 53733 78611 53789 78613
rect 53733 78559 53735 78611
rect 53735 78559 53787 78611
rect 53787 78559 53789 78611
rect 53733 78557 53789 78559
rect 55562 78611 55618 78613
rect 55562 78559 55564 78611
rect 55564 78559 55616 78611
rect 55616 78559 55618 78611
rect 55562 78557 55618 78559
rect 47403 78419 47459 78421
rect 47483 78419 47539 78421
rect 47563 78419 47619 78421
rect 47403 78367 47421 78419
rect 47421 78367 47459 78419
rect 47483 78367 47485 78419
rect 47485 78367 47537 78419
rect 47537 78367 47539 78419
rect 47563 78367 47601 78419
rect 47601 78367 47619 78419
rect 47403 78365 47459 78367
rect 47483 78365 47539 78367
rect 47563 78365 47619 78367
rect 49198 78418 49254 78420
rect 49278 78418 49334 78420
rect 49358 78418 49414 78420
rect 49198 78366 49216 78418
rect 49216 78366 49254 78418
rect 49278 78366 49280 78418
rect 49280 78366 49332 78418
rect 49332 78366 49334 78418
rect 49358 78366 49396 78418
rect 49396 78366 49414 78418
rect 49198 78364 49254 78366
rect 49278 78364 49334 78366
rect 49358 78364 49414 78366
rect 50998 78420 51054 78422
rect 51078 78420 51134 78422
rect 51158 78420 51214 78422
rect 50998 78368 51016 78420
rect 51016 78368 51054 78420
rect 51078 78368 51080 78420
rect 51080 78368 51132 78420
rect 51132 78368 51134 78420
rect 51158 78368 51196 78420
rect 51196 78368 51214 78420
rect 50998 78366 51054 78368
rect 51078 78366 51134 78368
rect 51158 78366 51214 78368
rect 52796 78419 52852 78421
rect 52876 78419 52932 78421
rect 52956 78419 53012 78421
rect 52796 78367 52814 78419
rect 52814 78367 52852 78419
rect 52876 78367 52878 78419
rect 52878 78367 52930 78419
rect 52930 78367 52932 78419
rect 52956 78367 52994 78419
rect 52994 78367 53012 78419
rect 52796 78365 52852 78367
rect 52876 78365 52932 78367
rect 52956 78365 53012 78367
rect 54594 78420 54650 78422
rect 54674 78420 54730 78422
rect 54754 78420 54810 78422
rect 54594 78368 54612 78420
rect 54612 78368 54650 78420
rect 54674 78368 54676 78420
rect 54676 78368 54728 78420
rect 54728 78368 54730 78420
rect 54754 78368 54792 78420
rect 54792 78368 54810 78420
rect 54594 78366 54650 78368
rect 54674 78366 54730 78368
rect 54754 78366 54810 78368
rect 56397 78419 56453 78421
rect 56477 78419 56533 78421
rect 56557 78419 56613 78421
rect 56397 78367 56415 78419
rect 56415 78367 56453 78419
rect 56477 78367 56479 78419
rect 56479 78367 56531 78419
rect 56531 78367 56533 78419
rect 56557 78367 56595 78419
rect 56595 78367 56613 78419
rect 56397 78365 56453 78367
rect 56477 78365 56533 78367
rect 56557 78365 56613 78367
rect 57274 78420 57330 78422
rect 57274 78368 57276 78420
rect 57276 78368 57328 78420
rect 57328 78368 57330 78420
rect 57274 78366 57330 78368
rect 48254 75243 48310 75261
rect 48254 75205 48256 75243
rect 48256 75205 48308 75243
rect 48308 75205 48310 75243
rect 49376 75209 49432 75265
rect 48254 75179 48310 75181
rect 48254 75127 48256 75179
rect 48256 75127 48308 75179
rect 48308 75127 48310 75179
rect 48254 75125 48310 75127
rect 48254 75063 48256 75101
rect 48256 75063 48308 75101
rect 48308 75063 48310 75101
rect 48254 75045 48310 75063
rect 30048 73736 30104 73738
rect 30128 73736 30184 73738
rect 30208 73736 30264 73738
rect 30288 73736 30344 73738
rect 30048 73684 30094 73736
rect 30094 73684 30104 73736
rect 30128 73684 30158 73736
rect 30158 73684 30170 73736
rect 30170 73684 30184 73736
rect 30208 73684 30222 73736
rect 30222 73684 30234 73736
rect 30234 73684 30264 73736
rect 30288 73684 30298 73736
rect 30298 73684 30344 73736
rect 30048 73682 30104 73684
rect 30128 73682 30184 73684
rect 30208 73682 30264 73684
rect 30288 73682 30344 73684
rect 30703 73429 30759 73431
rect 30783 73429 30839 73431
rect 30863 73429 30919 73431
rect 30703 73377 30741 73429
rect 30741 73377 30753 73429
rect 30753 73377 30759 73429
rect 30783 73377 30805 73429
rect 30805 73377 30817 73429
rect 30817 73377 30839 73429
rect 30863 73377 30869 73429
rect 30869 73377 30881 73429
rect 30881 73377 30919 73429
rect 30703 73375 30759 73377
rect 30783 73375 30839 73377
rect 30863 73375 30919 73377
rect 31038 73440 31094 73442
rect 31038 73388 31040 73440
rect 31040 73388 31092 73440
rect 31092 73388 31094 73440
rect 31038 73386 31094 73388
rect 31134 73194 31190 73196
rect 31214 73194 31270 73196
rect 31294 73194 31350 73196
rect 31374 73194 31430 73196
rect 31134 73142 31180 73194
rect 31180 73142 31190 73194
rect 31214 73142 31244 73194
rect 31244 73142 31256 73194
rect 31256 73142 31270 73194
rect 31294 73142 31308 73194
rect 31308 73142 31320 73194
rect 31320 73142 31350 73194
rect 31374 73142 31384 73194
rect 31384 73142 31430 73194
rect 31134 73140 31190 73142
rect 31214 73140 31270 73142
rect 31294 73140 31350 73142
rect 31374 73140 31430 73142
rect 30027 67266 30029 67296
rect 30029 67266 30081 67296
rect 30081 67266 30083 67296
rect 30027 67254 30083 67266
rect 30027 67240 30029 67254
rect 30029 67240 30081 67254
rect 30081 67240 30083 67254
rect 30027 67202 30029 67216
rect 30029 67202 30081 67216
rect 30081 67202 30083 67216
rect 30027 67190 30083 67202
rect 30027 67160 30029 67190
rect 30029 67160 30081 67190
rect 30081 67160 30083 67190
rect 30027 67126 30083 67136
rect 30027 67080 30029 67126
rect 30029 67080 30081 67126
rect 30081 67080 30083 67126
rect 30027 67010 30029 67056
rect 30029 67010 30081 67056
rect 30081 67010 30083 67056
rect 30027 67000 30083 67010
rect 43629 67077 43685 67079
rect 43629 67025 43631 67077
rect 43631 67025 43683 67077
rect 43683 67025 43685 67077
rect 43629 67023 43685 67025
rect 30027 66946 30029 66976
rect 30029 66946 30081 66976
rect 30081 66946 30083 66976
rect 30027 66934 30083 66946
rect 30027 66920 30029 66934
rect 30029 66920 30081 66934
rect 30081 66920 30083 66934
rect 30027 66882 30029 66896
rect 30029 66882 30081 66896
rect 30081 66882 30083 66896
rect 30027 66870 30083 66882
rect 30027 66840 30029 66870
rect 30029 66840 30081 66870
rect 30081 66840 30083 66870
rect 44405 66414 44461 66416
rect 44405 66362 44407 66414
rect 44407 66362 44459 66414
rect 44459 66362 44461 66414
rect 44405 66360 44461 66362
rect 30027 66125 30029 66155
rect 30029 66125 30081 66155
rect 30081 66125 30083 66155
rect 30027 66113 30083 66125
rect 30027 66099 30029 66113
rect 30029 66099 30081 66113
rect 30081 66099 30083 66113
rect 35623 66125 35679 66181
rect 30027 66061 30029 66075
rect 30029 66061 30081 66075
rect 30081 66061 30083 66075
rect 30027 66049 30083 66061
rect 30027 66019 30029 66049
rect 30029 66019 30081 66049
rect 30081 66019 30083 66049
rect 30027 65985 30083 65995
rect 30027 65939 30029 65985
rect 30029 65939 30081 65985
rect 30081 65939 30083 65985
rect 30027 65869 30029 65915
rect 30029 65869 30081 65915
rect 30081 65869 30083 65915
rect 30027 65859 30083 65869
rect 30027 65805 30029 65835
rect 30029 65805 30081 65835
rect 30081 65805 30083 65835
rect 30027 65793 30083 65805
rect 30027 65779 30029 65793
rect 30029 65779 30081 65793
rect 30081 65779 30083 65793
rect 30027 65741 30029 65755
rect 30029 65741 30081 65755
rect 30081 65741 30083 65755
rect 30027 65729 30083 65741
rect 30027 65699 30029 65729
rect 30029 65699 30081 65729
rect 30081 65699 30083 65729
rect 30027 65665 30083 65675
rect 30027 65619 30029 65665
rect 30029 65619 30081 65665
rect 30081 65619 30083 65665
rect 30027 65549 30029 65595
rect 30029 65549 30081 65595
rect 30081 65549 30083 65595
rect 30027 65539 30083 65549
rect 30027 65485 30029 65515
rect 30029 65485 30081 65515
rect 30081 65485 30083 65515
rect 30027 65473 30083 65485
rect 30027 65459 30029 65473
rect 30029 65459 30081 65473
rect 30081 65459 30083 65473
rect 30027 65421 30029 65435
rect 30029 65421 30081 65435
rect 30081 65421 30083 65435
rect 30027 65409 30083 65421
rect 30027 65379 30029 65409
rect 30029 65379 30081 65409
rect 30081 65379 30083 65409
rect 30027 65345 30083 65355
rect 30027 65299 30029 65345
rect 30029 65299 30081 65345
rect 30081 65299 30083 65345
rect 30027 65229 30029 65275
rect 30029 65229 30081 65275
rect 30081 65229 30083 65275
rect 30027 65219 30083 65229
rect 30027 65165 30029 65195
rect 30029 65165 30081 65195
rect 30081 65165 30083 65195
rect 30027 65153 30083 65165
rect 30027 65139 30029 65153
rect 30029 65139 30081 65153
rect 30081 65139 30083 65153
rect 30027 65101 30029 65115
rect 30029 65101 30081 65115
rect 30081 65101 30083 65115
rect 30027 65089 30083 65101
rect 30027 65059 30029 65089
rect 30029 65059 30081 65089
rect 30081 65059 30083 65089
rect 30032 64599 30034 64629
rect 30034 64599 30086 64629
rect 30086 64599 30088 64629
rect 30032 64587 30088 64599
rect 30032 64573 30034 64587
rect 30034 64573 30086 64587
rect 30086 64573 30088 64587
rect 30032 64535 30034 64549
rect 30034 64535 30086 64549
rect 30086 64535 30088 64549
rect 30032 64523 30088 64535
rect 30032 64493 30034 64523
rect 30034 64493 30086 64523
rect 30086 64493 30088 64523
rect 30032 64459 30088 64469
rect 30032 64413 30034 64459
rect 30034 64413 30086 64459
rect 30086 64413 30088 64459
rect 30032 64343 30034 64389
rect 30034 64343 30086 64389
rect 30086 64343 30088 64389
rect 30032 64333 30088 64343
rect 30032 64279 30034 64309
rect 30034 64279 30086 64309
rect 30086 64279 30088 64309
rect 30032 64267 30088 64279
rect 30032 64253 30034 64267
rect 30034 64253 30086 64267
rect 30086 64253 30088 64267
rect 30032 64215 30034 64229
rect 30034 64215 30086 64229
rect 30086 64215 30088 64229
rect 30032 64203 30088 64215
rect 30032 64173 30034 64203
rect 30034 64173 30086 64203
rect 30086 64173 30088 64203
rect 30032 64139 30088 64149
rect 30032 64093 30034 64139
rect 30034 64093 30086 64139
rect 30086 64093 30088 64139
rect 30032 64023 30034 64069
rect 30034 64023 30086 64069
rect 30086 64023 30088 64069
rect 30032 64013 30088 64023
rect 30032 63959 30034 63989
rect 30034 63959 30086 63989
rect 30086 63959 30088 63989
rect 30032 63947 30088 63959
rect 30032 63933 30034 63947
rect 30034 63933 30086 63947
rect 30086 63933 30088 63947
rect 30032 63895 30034 63909
rect 30034 63895 30086 63909
rect 30086 63895 30088 63909
rect 30032 63883 30088 63895
rect 30032 63853 30034 63883
rect 30034 63853 30086 63883
rect 30086 63853 30088 63883
rect 30032 63819 30088 63829
rect 30032 63773 30034 63819
rect 30034 63773 30086 63819
rect 30086 63773 30088 63819
rect 57459 77168 57469 84824
rect 57469 77168 57585 84824
rect 57585 77168 57595 84824
rect 67310 84834 67606 84836
rect 48239 74792 48295 74794
rect 48239 74740 48241 74792
rect 48241 74740 48293 74792
rect 48293 74740 48295 74792
rect 48239 74738 48295 74740
rect 48239 74676 48241 74714
rect 48241 74676 48293 74714
rect 48293 74676 48295 74714
rect 48239 74664 48295 74676
rect 48239 74658 48241 74664
rect 48241 74658 48293 74664
rect 48293 74658 48295 74664
rect 48239 74612 48241 74634
rect 48241 74612 48293 74634
rect 48293 74612 48295 74634
rect 48239 74600 48295 74612
rect 48239 74578 48241 74600
rect 48241 74578 48293 74600
rect 48293 74578 48295 74600
rect 48239 74548 48241 74554
rect 48241 74548 48293 74554
rect 48293 74548 48295 74554
rect 48239 74536 48295 74548
rect 48239 74498 48241 74536
rect 48241 74498 48293 74536
rect 48293 74498 48295 74536
rect 48239 74472 48295 74474
rect 48239 74420 48241 74472
rect 48241 74420 48293 74472
rect 48293 74420 48295 74472
rect 48239 74418 48295 74420
rect 48618 74403 48674 74459
rect 51438 74928 53174 75064
rect 53757 75065 54533 75075
rect 53757 74949 54533 75065
rect 53757 74939 54533 74949
rect 55456 75055 56312 75065
rect 55456 74939 56312 75055
rect 55456 74929 56312 74939
rect 57047 74783 57183 74793
rect 51186 74736 51322 74738
rect 51186 71804 51322 74736
rect 51186 71802 51322 71804
rect 57047 71787 57183 74783
rect 57047 71777 57183 71787
rect 67310 71662 67606 84834
rect 74529 84708 74531 84746
rect 74531 84708 74583 84746
rect 74583 84708 74585 84746
rect 74529 84696 74585 84708
rect 74529 84690 74531 84696
rect 74531 84690 74583 84696
rect 74583 84690 74585 84696
rect 74529 84644 74531 84666
rect 74531 84644 74583 84666
rect 74583 84644 74585 84666
rect 74529 84632 74585 84644
rect 74529 84610 74531 84632
rect 74531 84610 74583 84632
rect 74583 84610 74585 84632
rect 74529 84580 74531 84586
rect 74531 84580 74583 84586
rect 74583 84580 74585 84586
rect 74529 84568 74585 84580
rect 74529 84530 74531 84568
rect 74531 84530 74583 84568
rect 74583 84530 74585 84568
rect 74529 84504 74585 84506
rect 74529 84452 74531 84504
rect 74531 84452 74583 84504
rect 74583 84452 74585 84504
rect 74529 84450 74585 84452
rect 74529 84388 74531 84426
rect 74531 84388 74583 84426
rect 74583 84388 74585 84426
rect 74529 84376 74585 84388
rect 74529 84370 74531 84376
rect 74531 84370 74583 84376
rect 74583 84370 74585 84376
rect 74529 84324 74531 84346
rect 74531 84324 74583 84346
rect 74583 84324 74585 84346
rect 74529 84312 74585 84324
rect 74529 84290 74531 84312
rect 74531 84290 74583 84312
rect 74583 84290 74585 84312
rect 74529 84260 74531 84266
rect 74531 84260 74583 84266
rect 74583 84260 74585 84266
rect 74529 84248 74585 84260
rect 74529 84210 74531 84248
rect 74531 84210 74583 84248
rect 74583 84210 74585 84248
rect 75617 84708 75619 84746
rect 75619 84708 75671 84746
rect 75671 84708 75673 84746
rect 75617 84696 75673 84708
rect 75617 84690 75619 84696
rect 75619 84690 75671 84696
rect 75671 84690 75673 84696
rect 75617 84644 75619 84666
rect 75619 84644 75671 84666
rect 75671 84644 75673 84666
rect 75617 84632 75673 84644
rect 75617 84610 75619 84632
rect 75619 84610 75671 84632
rect 75671 84610 75673 84632
rect 75617 84580 75619 84586
rect 75619 84580 75671 84586
rect 75671 84580 75673 84586
rect 75617 84568 75673 84580
rect 75617 84530 75619 84568
rect 75619 84530 75671 84568
rect 75671 84530 75673 84568
rect 75617 84504 75673 84506
rect 75617 84452 75619 84504
rect 75619 84452 75671 84504
rect 75671 84452 75673 84504
rect 75617 84450 75673 84452
rect 75617 84388 75619 84426
rect 75619 84388 75671 84426
rect 75671 84388 75673 84426
rect 75617 84376 75673 84388
rect 75617 84370 75619 84376
rect 75619 84370 75671 84376
rect 75671 84370 75673 84376
rect 75617 84324 75619 84346
rect 75619 84324 75671 84346
rect 75671 84324 75673 84346
rect 75617 84312 75673 84324
rect 75617 84290 75619 84312
rect 75619 84290 75671 84312
rect 75671 84290 75673 84312
rect 75617 84260 75619 84266
rect 75619 84260 75671 84266
rect 75671 84260 75673 84266
rect 75617 84248 75673 84260
rect 75617 84210 75619 84248
rect 75619 84210 75671 84248
rect 75671 84210 75673 84248
rect 76705 84708 76707 84746
rect 76707 84708 76759 84746
rect 76759 84708 76761 84746
rect 76705 84696 76761 84708
rect 76705 84690 76707 84696
rect 76707 84690 76759 84696
rect 76759 84690 76761 84696
rect 76705 84644 76707 84666
rect 76707 84644 76759 84666
rect 76759 84644 76761 84666
rect 76705 84632 76761 84644
rect 76705 84610 76707 84632
rect 76707 84610 76759 84632
rect 76759 84610 76761 84632
rect 76705 84580 76707 84586
rect 76707 84580 76759 84586
rect 76759 84580 76761 84586
rect 76705 84568 76761 84580
rect 76705 84530 76707 84568
rect 76707 84530 76759 84568
rect 76759 84530 76761 84568
rect 76705 84504 76761 84506
rect 76705 84452 76707 84504
rect 76707 84452 76759 84504
rect 76759 84452 76761 84504
rect 76705 84450 76761 84452
rect 76705 84388 76707 84426
rect 76707 84388 76759 84426
rect 76759 84388 76761 84426
rect 76705 84376 76761 84388
rect 76705 84370 76707 84376
rect 76707 84370 76759 84376
rect 76759 84370 76761 84376
rect 76705 84324 76707 84346
rect 76707 84324 76759 84346
rect 76759 84324 76761 84346
rect 76705 84312 76761 84324
rect 76705 84290 76707 84312
rect 76707 84290 76759 84312
rect 76759 84290 76761 84312
rect 76705 84260 76707 84266
rect 76707 84260 76759 84266
rect 76759 84260 76761 84266
rect 76705 84248 76761 84260
rect 76705 84210 76707 84248
rect 76707 84210 76759 84248
rect 76759 84210 76761 84248
rect 77793 84708 77795 84746
rect 77795 84708 77847 84746
rect 77847 84708 77849 84746
rect 77793 84696 77849 84708
rect 77793 84690 77795 84696
rect 77795 84690 77847 84696
rect 77847 84690 77849 84696
rect 77793 84644 77795 84666
rect 77795 84644 77847 84666
rect 77847 84644 77849 84666
rect 77793 84632 77849 84644
rect 77793 84610 77795 84632
rect 77795 84610 77847 84632
rect 77847 84610 77849 84632
rect 77793 84580 77795 84586
rect 77795 84580 77847 84586
rect 77847 84580 77849 84586
rect 77793 84568 77849 84580
rect 77793 84530 77795 84568
rect 77795 84530 77847 84568
rect 77847 84530 77849 84568
rect 77793 84504 77849 84506
rect 77793 84452 77795 84504
rect 77795 84452 77847 84504
rect 77847 84452 77849 84504
rect 77793 84450 77849 84452
rect 77793 84388 77795 84426
rect 77795 84388 77847 84426
rect 77847 84388 77849 84426
rect 77793 84376 77849 84388
rect 77793 84370 77795 84376
rect 77795 84370 77847 84376
rect 77847 84370 77849 84376
rect 77793 84324 77795 84346
rect 77795 84324 77847 84346
rect 77847 84324 77849 84346
rect 77793 84312 77849 84324
rect 77793 84290 77795 84312
rect 77795 84290 77847 84312
rect 77847 84290 77849 84312
rect 77793 84260 77795 84266
rect 77795 84260 77847 84266
rect 77847 84260 77849 84266
rect 77793 84248 77849 84260
rect 77793 84210 77795 84248
rect 77795 84210 77847 84248
rect 77847 84210 77849 84248
rect 78881 84708 78883 84746
rect 78883 84708 78935 84746
rect 78935 84708 78937 84746
rect 78881 84696 78937 84708
rect 78881 84690 78883 84696
rect 78883 84690 78935 84696
rect 78935 84690 78937 84696
rect 78881 84644 78883 84666
rect 78883 84644 78935 84666
rect 78935 84644 78937 84666
rect 78881 84632 78937 84644
rect 78881 84610 78883 84632
rect 78883 84610 78935 84632
rect 78935 84610 78937 84632
rect 78881 84580 78883 84586
rect 78883 84580 78935 84586
rect 78935 84580 78937 84586
rect 78881 84568 78937 84580
rect 78881 84530 78883 84568
rect 78883 84530 78935 84568
rect 78935 84530 78937 84568
rect 78881 84504 78937 84506
rect 78881 84452 78883 84504
rect 78883 84452 78935 84504
rect 78935 84452 78937 84504
rect 78881 84450 78937 84452
rect 78881 84388 78883 84426
rect 78883 84388 78935 84426
rect 78935 84388 78937 84426
rect 78881 84376 78937 84388
rect 78881 84370 78883 84376
rect 78883 84370 78935 84376
rect 78935 84370 78937 84376
rect 78881 84324 78883 84346
rect 78883 84324 78935 84346
rect 78935 84324 78937 84346
rect 78881 84312 78937 84324
rect 78881 84290 78883 84312
rect 78883 84290 78935 84312
rect 78935 84290 78937 84312
rect 78881 84260 78883 84266
rect 78883 84260 78935 84266
rect 78935 84260 78937 84266
rect 78881 84248 78937 84260
rect 78881 84210 78883 84248
rect 78883 84210 78935 84248
rect 78935 84210 78937 84248
rect 79969 84708 79971 84746
rect 79971 84708 80023 84746
rect 80023 84708 80025 84746
rect 79969 84696 80025 84708
rect 79969 84690 79971 84696
rect 79971 84690 80023 84696
rect 80023 84690 80025 84696
rect 79969 84644 79971 84666
rect 79971 84644 80023 84666
rect 80023 84644 80025 84666
rect 79969 84632 80025 84644
rect 79969 84610 79971 84632
rect 79971 84610 80023 84632
rect 80023 84610 80025 84632
rect 79969 84580 79971 84586
rect 79971 84580 80023 84586
rect 80023 84580 80025 84586
rect 79969 84568 80025 84580
rect 79969 84530 79971 84568
rect 79971 84530 80023 84568
rect 80023 84530 80025 84568
rect 79969 84504 80025 84506
rect 79969 84452 79971 84504
rect 79971 84452 80023 84504
rect 80023 84452 80025 84504
rect 79969 84450 80025 84452
rect 79969 84388 79971 84426
rect 79971 84388 80023 84426
rect 80023 84388 80025 84426
rect 79969 84376 80025 84388
rect 79969 84370 79971 84376
rect 79971 84370 80023 84376
rect 80023 84370 80025 84376
rect 79969 84324 79971 84346
rect 79971 84324 80023 84346
rect 80023 84324 80025 84346
rect 79969 84312 80025 84324
rect 79969 84290 79971 84312
rect 79971 84290 80023 84312
rect 80023 84290 80025 84312
rect 79969 84260 79971 84266
rect 79971 84260 80023 84266
rect 80023 84260 80025 84266
rect 79969 84248 80025 84260
rect 79969 84210 79971 84248
rect 79971 84210 80023 84248
rect 80023 84210 80025 84248
rect 81057 84708 81059 84746
rect 81059 84708 81111 84746
rect 81111 84708 81113 84746
rect 81057 84696 81113 84708
rect 81057 84690 81059 84696
rect 81059 84690 81111 84696
rect 81111 84690 81113 84696
rect 81057 84644 81059 84666
rect 81059 84644 81111 84666
rect 81111 84644 81113 84666
rect 81057 84632 81113 84644
rect 81057 84610 81059 84632
rect 81059 84610 81111 84632
rect 81111 84610 81113 84632
rect 81057 84580 81059 84586
rect 81059 84580 81111 84586
rect 81111 84580 81113 84586
rect 81057 84568 81113 84580
rect 81057 84530 81059 84568
rect 81059 84530 81111 84568
rect 81111 84530 81113 84568
rect 81057 84504 81113 84506
rect 81057 84452 81059 84504
rect 81059 84452 81111 84504
rect 81111 84452 81113 84504
rect 81057 84450 81113 84452
rect 81057 84388 81059 84426
rect 81059 84388 81111 84426
rect 81111 84388 81113 84426
rect 81057 84376 81113 84388
rect 81057 84370 81059 84376
rect 81059 84370 81111 84376
rect 81111 84370 81113 84376
rect 81057 84324 81059 84346
rect 81059 84324 81111 84346
rect 81111 84324 81113 84346
rect 81057 84312 81113 84324
rect 81057 84290 81059 84312
rect 81059 84290 81111 84312
rect 81111 84290 81113 84312
rect 81057 84260 81059 84266
rect 81059 84260 81111 84266
rect 81111 84260 81113 84266
rect 81057 84248 81113 84260
rect 81057 84210 81059 84248
rect 81059 84210 81111 84248
rect 81111 84210 81113 84248
rect 82145 84708 82147 84746
rect 82147 84708 82199 84746
rect 82199 84708 82201 84746
rect 82145 84696 82201 84708
rect 82145 84690 82147 84696
rect 82147 84690 82199 84696
rect 82199 84690 82201 84696
rect 82145 84644 82147 84666
rect 82147 84644 82199 84666
rect 82199 84644 82201 84666
rect 82145 84632 82201 84644
rect 82145 84610 82147 84632
rect 82147 84610 82199 84632
rect 82199 84610 82201 84632
rect 82145 84580 82147 84586
rect 82147 84580 82199 84586
rect 82199 84580 82201 84586
rect 82145 84568 82201 84580
rect 82145 84530 82147 84568
rect 82147 84530 82199 84568
rect 82199 84530 82201 84568
rect 82145 84504 82201 84506
rect 82145 84452 82147 84504
rect 82147 84452 82199 84504
rect 82199 84452 82201 84504
rect 82145 84450 82201 84452
rect 82145 84388 82147 84426
rect 82147 84388 82199 84426
rect 82199 84388 82201 84426
rect 82145 84376 82201 84388
rect 82145 84370 82147 84376
rect 82147 84370 82199 84376
rect 82199 84370 82201 84376
rect 82145 84324 82147 84346
rect 82147 84324 82199 84346
rect 82199 84324 82201 84346
rect 82145 84312 82201 84324
rect 82145 84290 82147 84312
rect 82147 84290 82199 84312
rect 82199 84290 82201 84312
rect 82145 84260 82147 84266
rect 82147 84260 82199 84266
rect 82199 84260 82201 84266
rect 82145 84248 82201 84260
rect 82145 84210 82147 84248
rect 82147 84210 82199 84248
rect 82199 84210 82201 84248
rect 83233 84708 83235 84746
rect 83235 84708 83287 84746
rect 83287 84708 83289 84746
rect 83233 84696 83289 84708
rect 83233 84690 83235 84696
rect 83235 84690 83287 84696
rect 83287 84690 83289 84696
rect 83233 84644 83235 84666
rect 83235 84644 83287 84666
rect 83287 84644 83289 84666
rect 83233 84632 83289 84644
rect 83233 84610 83235 84632
rect 83235 84610 83287 84632
rect 83287 84610 83289 84632
rect 83233 84580 83235 84586
rect 83235 84580 83287 84586
rect 83287 84580 83289 84586
rect 83233 84568 83289 84580
rect 83233 84530 83235 84568
rect 83235 84530 83287 84568
rect 83287 84530 83289 84568
rect 83233 84504 83289 84506
rect 83233 84452 83235 84504
rect 83235 84452 83287 84504
rect 83287 84452 83289 84504
rect 83233 84450 83289 84452
rect 83233 84388 83235 84426
rect 83235 84388 83287 84426
rect 83287 84388 83289 84426
rect 83233 84376 83289 84388
rect 83233 84370 83235 84376
rect 83235 84370 83287 84376
rect 83287 84370 83289 84376
rect 83233 84324 83235 84346
rect 83235 84324 83287 84346
rect 83287 84324 83289 84346
rect 83233 84312 83289 84324
rect 83233 84290 83235 84312
rect 83235 84290 83287 84312
rect 83287 84290 83289 84312
rect 83233 84260 83235 84266
rect 83235 84260 83287 84266
rect 83287 84260 83289 84266
rect 83233 84248 83289 84260
rect 83233 84210 83235 84248
rect 83235 84210 83287 84248
rect 83287 84210 83289 84248
rect 84321 84708 84323 84746
rect 84323 84708 84375 84746
rect 84375 84708 84377 84746
rect 84321 84696 84377 84708
rect 84321 84690 84323 84696
rect 84323 84690 84375 84696
rect 84375 84690 84377 84696
rect 84321 84644 84323 84666
rect 84323 84644 84375 84666
rect 84375 84644 84377 84666
rect 84321 84632 84377 84644
rect 84321 84610 84323 84632
rect 84323 84610 84375 84632
rect 84375 84610 84377 84632
rect 84321 84580 84323 84586
rect 84323 84580 84375 84586
rect 84375 84580 84377 84586
rect 84321 84568 84377 84580
rect 84321 84530 84323 84568
rect 84323 84530 84375 84568
rect 84375 84530 84377 84568
rect 84321 84504 84377 84506
rect 84321 84452 84323 84504
rect 84323 84452 84375 84504
rect 84375 84452 84377 84504
rect 84321 84450 84377 84452
rect 84321 84388 84323 84426
rect 84323 84388 84375 84426
rect 84375 84388 84377 84426
rect 84321 84376 84377 84388
rect 84321 84370 84323 84376
rect 84323 84370 84375 84376
rect 84375 84370 84377 84376
rect 84321 84324 84323 84346
rect 84323 84324 84375 84346
rect 84375 84324 84377 84346
rect 84321 84312 84377 84324
rect 84321 84290 84323 84312
rect 84323 84290 84375 84312
rect 84375 84290 84377 84312
rect 84321 84260 84323 84266
rect 84323 84260 84375 84266
rect 84375 84260 84377 84266
rect 84321 84248 84377 84260
rect 84321 84210 84323 84248
rect 84323 84210 84375 84248
rect 84375 84210 84377 84248
rect 85409 84708 85411 84746
rect 85411 84708 85463 84746
rect 85463 84708 85465 84746
rect 85409 84696 85465 84708
rect 85409 84690 85411 84696
rect 85411 84690 85463 84696
rect 85463 84690 85465 84696
rect 85409 84644 85411 84666
rect 85411 84644 85463 84666
rect 85463 84644 85465 84666
rect 85409 84632 85465 84644
rect 85409 84610 85411 84632
rect 85411 84610 85463 84632
rect 85463 84610 85465 84632
rect 85409 84580 85411 84586
rect 85411 84580 85463 84586
rect 85463 84580 85465 84586
rect 85409 84568 85465 84580
rect 85409 84530 85411 84568
rect 85411 84530 85463 84568
rect 85463 84530 85465 84568
rect 85409 84504 85465 84506
rect 85409 84452 85411 84504
rect 85411 84452 85463 84504
rect 85463 84452 85465 84504
rect 85409 84450 85465 84452
rect 85409 84388 85411 84426
rect 85411 84388 85463 84426
rect 85463 84388 85465 84426
rect 85409 84376 85465 84388
rect 85409 84370 85411 84376
rect 85411 84370 85463 84376
rect 85463 84370 85465 84376
rect 85409 84324 85411 84346
rect 85411 84324 85463 84346
rect 85463 84324 85465 84346
rect 85409 84312 85465 84324
rect 85409 84290 85411 84312
rect 85411 84290 85463 84312
rect 85463 84290 85465 84312
rect 85409 84260 85411 84266
rect 85411 84260 85463 84266
rect 85463 84260 85465 84266
rect 85409 84248 85465 84260
rect 85409 84210 85411 84248
rect 85411 84210 85463 84248
rect 85463 84210 85465 84248
rect 86497 84708 86499 84746
rect 86499 84708 86551 84746
rect 86551 84708 86553 84746
rect 86497 84696 86553 84708
rect 86497 84690 86499 84696
rect 86499 84690 86551 84696
rect 86551 84690 86553 84696
rect 86497 84644 86499 84666
rect 86499 84644 86551 84666
rect 86551 84644 86553 84666
rect 86497 84632 86553 84644
rect 86497 84610 86499 84632
rect 86499 84610 86551 84632
rect 86551 84610 86553 84632
rect 86497 84580 86499 84586
rect 86499 84580 86551 84586
rect 86551 84580 86553 84586
rect 86497 84568 86553 84580
rect 86497 84530 86499 84568
rect 86499 84530 86551 84568
rect 86551 84530 86553 84568
rect 86497 84504 86553 84506
rect 86497 84452 86499 84504
rect 86499 84452 86551 84504
rect 86551 84452 86553 84504
rect 86497 84450 86553 84452
rect 86497 84388 86499 84426
rect 86499 84388 86551 84426
rect 86551 84388 86553 84426
rect 86497 84376 86553 84388
rect 86497 84370 86499 84376
rect 86499 84370 86551 84376
rect 86551 84370 86553 84376
rect 86497 84324 86499 84346
rect 86499 84324 86551 84346
rect 86551 84324 86553 84346
rect 86497 84312 86553 84324
rect 86497 84290 86499 84312
rect 86499 84290 86551 84312
rect 86551 84290 86553 84312
rect 86497 84260 86499 84266
rect 86499 84260 86551 84266
rect 86551 84260 86553 84266
rect 86497 84248 86553 84260
rect 86497 84210 86499 84248
rect 86499 84210 86551 84248
rect 86551 84210 86553 84248
rect 87585 84708 87587 84746
rect 87587 84708 87639 84746
rect 87639 84708 87641 84746
rect 87585 84696 87641 84708
rect 87585 84690 87587 84696
rect 87587 84690 87639 84696
rect 87639 84690 87641 84696
rect 87585 84644 87587 84666
rect 87587 84644 87639 84666
rect 87639 84644 87641 84666
rect 87585 84632 87641 84644
rect 87585 84610 87587 84632
rect 87587 84610 87639 84632
rect 87639 84610 87641 84632
rect 87585 84580 87587 84586
rect 87587 84580 87639 84586
rect 87639 84580 87641 84586
rect 87585 84568 87641 84580
rect 87585 84530 87587 84568
rect 87587 84530 87639 84568
rect 87639 84530 87641 84568
rect 87585 84504 87641 84506
rect 87585 84452 87587 84504
rect 87587 84452 87639 84504
rect 87639 84452 87641 84504
rect 87585 84450 87641 84452
rect 87585 84388 87587 84426
rect 87587 84388 87639 84426
rect 87639 84388 87641 84426
rect 87585 84376 87641 84388
rect 87585 84370 87587 84376
rect 87587 84370 87639 84376
rect 87639 84370 87641 84376
rect 87585 84324 87587 84346
rect 87587 84324 87639 84346
rect 87639 84324 87641 84346
rect 87585 84312 87641 84324
rect 87585 84290 87587 84312
rect 87587 84290 87639 84312
rect 87639 84290 87641 84312
rect 87585 84260 87587 84266
rect 87587 84260 87639 84266
rect 87639 84260 87641 84266
rect 87585 84248 87641 84260
rect 87585 84210 87587 84248
rect 87587 84210 87639 84248
rect 87639 84210 87641 84248
rect 88673 84708 88675 84746
rect 88675 84708 88727 84746
rect 88727 84708 88729 84746
rect 88673 84696 88729 84708
rect 88673 84690 88675 84696
rect 88675 84690 88727 84696
rect 88727 84690 88729 84696
rect 88673 84644 88675 84666
rect 88675 84644 88727 84666
rect 88727 84644 88729 84666
rect 88673 84632 88729 84644
rect 88673 84610 88675 84632
rect 88675 84610 88727 84632
rect 88727 84610 88729 84632
rect 88673 84580 88675 84586
rect 88675 84580 88727 84586
rect 88727 84580 88729 84586
rect 88673 84568 88729 84580
rect 88673 84530 88675 84568
rect 88675 84530 88727 84568
rect 88727 84530 88729 84568
rect 88673 84504 88729 84506
rect 88673 84452 88675 84504
rect 88675 84452 88727 84504
rect 88727 84452 88729 84504
rect 88673 84450 88729 84452
rect 88673 84388 88675 84426
rect 88675 84388 88727 84426
rect 88727 84388 88729 84426
rect 88673 84376 88729 84388
rect 88673 84370 88675 84376
rect 88675 84370 88727 84376
rect 88727 84370 88729 84376
rect 88673 84324 88675 84346
rect 88675 84324 88727 84346
rect 88727 84324 88729 84346
rect 88673 84312 88729 84324
rect 88673 84290 88675 84312
rect 88675 84290 88727 84312
rect 88727 84290 88729 84312
rect 88673 84260 88675 84266
rect 88675 84260 88727 84266
rect 88727 84260 88729 84266
rect 88673 84248 88729 84260
rect 88673 84210 88675 84248
rect 88675 84210 88727 84248
rect 88727 84210 88729 84248
rect 75074 82705 75076 82743
rect 75076 82705 75128 82743
rect 75128 82705 75130 82743
rect 75074 82693 75130 82705
rect 75074 82687 75076 82693
rect 75076 82687 75128 82693
rect 75128 82687 75130 82693
rect 75074 82641 75076 82663
rect 75076 82641 75128 82663
rect 75128 82641 75130 82663
rect 75074 82629 75130 82641
rect 75074 82607 75076 82629
rect 75076 82607 75128 82629
rect 75128 82607 75130 82629
rect 75074 82577 75076 82583
rect 75076 82577 75128 82583
rect 75128 82577 75130 82583
rect 75074 82565 75130 82577
rect 75074 82527 75076 82565
rect 75076 82527 75128 82565
rect 75128 82527 75130 82565
rect 75074 82501 75130 82503
rect 75074 82449 75076 82501
rect 75076 82449 75128 82501
rect 75128 82449 75130 82501
rect 75074 82447 75130 82449
rect 75074 82385 75076 82423
rect 75076 82385 75128 82423
rect 75128 82385 75130 82423
rect 75074 82373 75130 82385
rect 75074 82367 75076 82373
rect 75076 82367 75128 82373
rect 75128 82367 75130 82373
rect 75074 82321 75076 82343
rect 75076 82321 75128 82343
rect 75128 82321 75130 82343
rect 75074 82309 75130 82321
rect 75074 82287 75076 82309
rect 75076 82287 75128 82309
rect 75128 82287 75130 82309
rect 75074 82257 75076 82263
rect 75076 82257 75128 82263
rect 75128 82257 75130 82263
rect 75074 82245 75130 82257
rect 75074 82207 75076 82245
rect 75076 82207 75128 82245
rect 75128 82207 75130 82245
rect 76162 82705 76164 82743
rect 76164 82705 76216 82743
rect 76216 82705 76218 82743
rect 76162 82693 76218 82705
rect 76162 82687 76164 82693
rect 76164 82687 76216 82693
rect 76216 82687 76218 82693
rect 76162 82641 76164 82663
rect 76164 82641 76216 82663
rect 76216 82641 76218 82663
rect 76162 82629 76218 82641
rect 76162 82607 76164 82629
rect 76164 82607 76216 82629
rect 76216 82607 76218 82629
rect 76162 82577 76164 82583
rect 76164 82577 76216 82583
rect 76216 82577 76218 82583
rect 76162 82565 76218 82577
rect 76162 82527 76164 82565
rect 76164 82527 76216 82565
rect 76216 82527 76218 82565
rect 76162 82501 76218 82503
rect 76162 82449 76164 82501
rect 76164 82449 76216 82501
rect 76216 82449 76218 82501
rect 76162 82447 76218 82449
rect 76162 82385 76164 82423
rect 76164 82385 76216 82423
rect 76216 82385 76218 82423
rect 76162 82373 76218 82385
rect 76162 82367 76164 82373
rect 76164 82367 76216 82373
rect 76216 82367 76218 82373
rect 76162 82321 76164 82343
rect 76164 82321 76216 82343
rect 76216 82321 76218 82343
rect 76162 82309 76218 82321
rect 76162 82287 76164 82309
rect 76164 82287 76216 82309
rect 76216 82287 76218 82309
rect 76162 82257 76164 82263
rect 76164 82257 76216 82263
rect 76216 82257 76218 82263
rect 76162 82245 76218 82257
rect 76162 82207 76164 82245
rect 76164 82207 76216 82245
rect 76216 82207 76218 82245
rect 77250 82705 77252 82743
rect 77252 82705 77304 82743
rect 77304 82705 77306 82743
rect 77250 82693 77306 82705
rect 77250 82687 77252 82693
rect 77252 82687 77304 82693
rect 77304 82687 77306 82693
rect 77250 82641 77252 82663
rect 77252 82641 77304 82663
rect 77304 82641 77306 82663
rect 77250 82629 77306 82641
rect 77250 82607 77252 82629
rect 77252 82607 77304 82629
rect 77304 82607 77306 82629
rect 77250 82577 77252 82583
rect 77252 82577 77304 82583
rect 77304 82577 77306 82583
rect 77250 82565 77306 82577
rect 77250 82527 77252 82565
rect 77252 82527 77304 82565
rect 77304 82527 77306 82565
rect 77250 82501 77306 82503
rect 77250 82449 77252 82501
rect 77252 82449 77304 82501
rect 77304 82449 77306 82501
rect 77250 82447 77306 82449
rect 77250 82385 77252 82423
rect 77252 82385 77304 82423
rect 77304 82385 77306 82423
rect 77250 82373 77306 82385
rect 77250 82367 77252 82373
rect 77252 82367 77304 82373
rect 77304 82367 77306 82373
rect 77250 82321 77252 82343
rect 77252 82321 77304 82343
rect 77304 82321 77306 82343
rect 77250 82309 77306 82321
rect 77250 82287 77252 82309
rect 77252 82287 77304 82309
rect 77304 82287 77306 82309
rect 77250 82257 77252 82263
rect 77252 82257 77304 82263
rect 77304 82257 77306 82263
rect 77250 82245 77306 82257
rect 77250 82207 77252 82245
rect 77252 82207 77304 82245
rect 77304 82207 77306 82245
rect 78338 82705 78340 82743
rect 78340 82705 78392 82743
rect 78392 82705 78394 82743
rect 78338 82693 78394 82705
rect 78338 82687 78340 82693
rect 78340 82687 78392 82693
rect 78392 82687 78394 82693
rect 78338 82641 78340 82663
rect 78340 82641 78392 82663
rect 78392 82641 78394 82663
rect 78338 82629 78394 82641
rect 78338 82607 78340 82629
rect 78340 82607 78392 82629
rect 78392 82607 78394 82629
rect 78338 82577 78340 82583
rect 78340 82577 78392 82583
rect 78392 82577 78394 82583
rect 78338 82565 78394 82577
rect 78338 82527 78340 82565
rect 78340 82527 78392 82565
rect 78392 82527 78394 82565
rect 78338 82501 78394 82503
rect 78338 82449 78340 82501
rect 78340 82449 78392 82501
rect 78392 82449 78394 82501
rect 78338 82447 78394 82449
rect 78338 82385 78340 82423
rect 78340 82385 78392 82423
rect 78392 82385 78394 82423
rect 78338 82373 78394 82385
rect 78338 82367 78340 82373
rect 78340 82367 78392 82373
rect 78392 82367 78394 82373
rect 78338 82321 78340 82343
rect 78340 82321 78392 82343
rect 78392 82321 78394 82343
rect 78338 82309 78394 82321
rect 78338 82287 78340 82309
rect 78340 82287 78392 82309
rect 78392 82287 78394 82309
rect 78338 82257 78340 82263
rect 78340 82257 78392 82263
rect 78392 82257 78394 82263
rect 78338 82245 78394 82257
rect 78338 82207 78340 82245
rect 78340 82207 78392 82245
rect 78392 82207 78394 82245
rect 79426 82705 79428 82743
rect 79428 82705 79480 82743
rect 79480 82705 79482 82743
rect 79426 82693 79482 82705
rect 79426 82687 79428 82693
rect 79428 82687 79480 82693
rect 79480 82687 79482 82693
rect 79426 82641 79428 82663
rect 79428 82641 79480 82663
rect 79480 82641 79482 82663
rect 79426 82629 79482 82641
rect 79426 82607 79428 82629
rect 79428 82607 79480 82629
rect 79480 82607 79482 82629
rect 79426 82577 79428 82583
rect 79428 82577 79480 82583
rect 79480 82577 79482 82583
rect 79426 82565 79482 82577
rect 79426 82527 79428 82565
rect 79428 82527 79480 82565
rect 79480 82527 79482 82565
rect 79426 82501 79482 82503
rect 79426 82449 79428 82501
rect 79428 82449 79480 82501
rect 79480 82449 79482 82501
rect 79426 82447 79482 82449
rect 79426 82385 79428 82423
rect 79428 82385 79480 82423
rect 79480 82385 79482 82423
rect 79426 82373 79482 82385
rect 79426 82367 79428 82373
rect 79428 82367 79480 82373
rect 79480 82367 79482 82373
rect 79426 82321 79428 82343
rect 79428 82321 79480 82343
rect 79480 82321 79482 82343
rect 79426 82309 79482 82321
rect 79426 82287 79428 82309
rect 79428 82287 79480 82309
rect 79480 82287 79482 82309
rect 79426 82257 79428 82263
rect 79428 82257 79480 82263
rect 79480 82257 79482 82263
rect 79426 82245 79482 82257
rect 79426 82207 79428 82245
rect 79428 82207 79480 82245
rect 79480 82207 79482 82245
rect 80514 82705 80516 82743
rect 80516 82705 80568 82743
rect 80568 82705 80570 82743
rect 80514 82693 80570 82705
rect 80514 82687 80516 82693
rect 80516 82687 80568 82693
rect 80568 82687 80570 82693
rect 80514 82641 80516 82663
rect 80516 82641 80568 82663
rect 80568 82641 80570 82663
rect 80514 82629 80570 82641
rect 80514 82607 80516 82629
rect 80516 82607 80568 82629
rect 80568 82607 80570 82629
rect 80514 82577 80516 82583
rect 80516 82577 80568 82583
rect 80568 82577 80570 82583
rect 80514 82565 80570 82577
rect 80514 82527 80516 82565
rect 80516 82527 80568 82565
rect 80568 82527 80570 82565
rect 80514 82501 80570 82503
rect 80514 82449 80516 82501
rect 80516 82449 80568 82501
rect 80568 82449 80570 82501
rect 80514 82447 80570 82449
rect 80514 82385 80516 82423
rect 80516 82385 80568 82423
rect 80568 82385 80570 82423
rect 80514 82373 80570 82385
rect 80514 82367 80516 82373
rect 80516 82367 80568 82373
rect 80568 82367 80570 82373
rect 80514 82321 80516 82343
rect 80516 82321 80568 82343
rect 80568 82321 80570 82343
rect 80514 82309 80570 82321
rect 80514 82287 80516 82309
rect 80516 82287 80568 82309
rect 80568 82287 80570 82309
rect 80514 82257 80516 82263
rect 80516 82257 80568 82263
rect 80568 82257 80570 82263
rect 80514 82245 80570 82257
rect 80514 82207 80516 82245
rect 80516 82207 80568 82245
rect 80568 82207 80570 82245
rect 81602 82705 81604 82743
rect 81604 82705 81656 82743
rect 81656 82705 81658 82743
rect 81602 82693 81658 82705
rect 81602 82687 81604 82693
rect 81604 82687 81656 82693
rect 81656 82687 81658 82693
rect 81602 82641 81604 82663
rect 81604 82641 81656 82663
rect 81656 82641 81658 82663
rect 81602 82629 81658 82641
rect 81602 82607 81604 82629
rect 81604 82607 81656 82629
rect 81656 82607 81658 82629
rect 81602 82577 81604 82583
rect 81604 82577 81656 82583
rect 81656 82577 81658 82583
rect 81602 82565 81658 82577
rect 81602 82527 81604 82565
rect 81604 82527 81656 82565
rect 81656 82527 81658 82565
rect 81602 82501 81658 82503
rect 81602 82449 81604 82501
rect 81604 82449 81656 82501
rect 81656 82449 81658 82501
rect 81602 82447 81658 82449
rect 81602 82385 81604 82423
rect 81604 82385 81656 82423
rect 81656 82385 81658 82423
rect 81602 82373 81658 82385
rect 81602 82367 81604 82373
rect 81604 82367 81656 82373
rect 81656 82367 81658 82373
rect 81602 82321 81604 82343
rect 81604 82321 81656 82343
rect 81656 82321 81658 82343
rect 81602 82309 81658 82321
rect 81602 82287 81604 82309
rect 81604 82287 81656 82309
rect 81656 82287 81658 82309
rect 81602 82257 81604 82263
rect 81604 82257 81656 82263
rect 81656 82257 81658 82263
rect 81602 82245 81658 82257
rect 81602 82207 81604 82245
rect 81604 82207 81656 82245
rect 81656 82207 81658 82245
rect 82690 82705 82692 82743
rect 82692 82705 82744 82743
rect 82744 82705 82746 82743
rect 82690 82693 82746 82705
rect 82690 82687 82692 82693
rect 82692 82687 82744 82693
rect 82744 82687 82746 82693
rect 82690 82641 82692 82663
rect 82692 82641 82744 82663
rect 82744 82641 82746 82663
rect 82690 82629 82746 82641
rect 82690 82607 82692 82629
rect 82692 82607 82744 82629
rect 82744 82607 82746 82629
rect 82690 82577 82692 82583
rect 82692 82577 82744 82583
rect 82744 82577 82746 82583
rect 82690 82565 82746 82577
rect 82690 82527 82692 82565
rect 82692 82527 82744 82565
rect 82744 82527 82746 82565
rect 82690 82501 82746 82503
rect 82690 82449 82692 82501
rect 82692 82449 82744 82501
rect 82744 82449 82746 82501
rect 82690 82447 82746 82449
rect 82690 82385 82692 82423
rect 82692 82385 82744 82423
rect 82744 82385 82746 82423
rect 82690 82373 82746 82385
rect 82690 82367 82692 82373
rect 82692 82367 82744 82373
rect 82744 82367 82746 82373
rect 82690 82321 82692 82343
rect 82692 82321 82744 82343
rect 82744 82321 82746 82343
rect 82690 82309 82746 82321
rect 82690 82287 82692 82309
rect 82692 82287 82744 82309
rect 82744 82287 82746 82309
rect 82690 82257 82692 82263
rect 82692 82257 82744 82263
rect 82744 82257 82746 82263
rect 82690 82245 82746 82257
rect 82690 82207 82692 82245
rect 82692 82207 82744 82245
rect 82744 82207 82746 82245
rect 83778 82705 83780 82743
rect 83780 82705 83832 82743
rect 83832 82705 83834 82743
rect 83778 82693 83834 82705
rect 83778 82687 83780 82693
rect 83780 82687 83832 82693
rect 83832 82687 83834 82693
rect 83778 82641 83780 82663
rect 83780 82641 83832 82663
rect 83832 82641 83834 82663
rect 83778 82629 83834 82641
rect 83778 82607 83780 82629
rect 83780 82607 83832 82629
rect 83832 82607 83834 82629
rect 83778 82577 83780 82583
rect 83780 82577 83832 82583
rect 83832 82577 83834 82583
rect 83778 82565 83834 82577
rect 83778 82527 83780 82565
rect 83780 82527 83832 82565
rect 83832 82527 83834 82565
rect 83778 82501 83834 82503
rect 83778 82449 83780 82501
rect 83780 82449 83832 82501
rect 83832 82449 83834 82501
rect 83778 82447 83834 82449
rect 83778 82385 83780 82423
rect 83780 82385 83832 82423
rect 83832 82385 83834 82423
rect 83778 82373 83834 82385
rect 83778 82367 83780 82373
rect 83780 82367 83832 82373
rect 83832 82367 83834 82373
rect 83778 82321 83780 82343
rect 83780 82321 83832 82343
rect 83832 82321 83834 82343
rect 83778 82309 83834 82321
rect 83778 82287 83780 82309
rect 83780 82287 83832 82309
rect 83832 82287 83834 82309
rect 83778 82257 83780 82263
rect 83780 82257 83832 82263
rect 83832 82257 83834 82263
rect 83778 82245 83834 82257
rect 83778 82207 83780 82245
rect 83780 82207 83832 82245
rect 83832 82207 83834 82245
rect 84866 82705 84868 82743
rect 84868 82705 84920 82743
rect 84920 82705 84922 82743
rect 84866 82693 84922 82705
rect 84866 82687 84868 82693
rect 84868 82687 84920 82693
rect 84920 82687 84922 82693
rect 84866 82641 84868 82663
rect 84868 82641 84920 82663
rect 84920 82641 84922 82663
rect 84866 82629 84922 82641
rect 84866 82607 84868 82629
rect 84868 82607 84920 82629
rect 84920 82607 84922 82629
rect 84866 82577 84868 82583
rect 84868 82577 84920 82583
rect 84920 82577 84922 82583
rect 84866 82565 84922 82577
rect 84866 82527 84868 82565
rect 84868 82527 84920 82565
rect 84920 82527 84922 82565
rect 84866 82501 84922 82503
rect 84866 82449 84868 82501
rect 84868 82449 84920 82501
rect 84920 82449 84922 82501
rect 84866 82447 84922 82449
rect 84866 82385 84868 82423
rect 84868 82385 84920 82423
rect 84920 82385 84922 82423
rect 84866 82373 84922 82385
rect 84866 82367 84868 82373
rect 84868 82367 84920 82373
rect 84920 82367 84922 82373
rect 84866 82321 84868 82343
rect 84868 82321 84920 82343
rect 84920 82321 84922 82343
rect 84866 82309 84922 82321
rect 84866 82287 84868 82309
rect 84868 82287 84920 82309
rect 84920 82287 84922 82309
rect 84866 82257 84868 82263
rect 84868 82257 84920 82263
rect 84920 82257 84922 82263
rect 84866 82245 84922 82257
rect 84866 82207 84868 82245
rect 84868 82207 84920 82245
rect 84920 82207 84922 82245
rect 85954 82705 85956 82743
rect 85956 82705 86008 82743
rect 86008 82705 86010 82743
rect 85954 82693 86010 82705
rect 85954 82687 85956 82693
rect 85956 82687 86008 82693
rect 86008 82687 86010 82693
rect 85954 82641 85956 82663
rect 85956 82641 86008 82663
rect 86008 82641 86010 82663
rect 85954 82629 86010 82641
rect 85954 82607 85956 82629
rect 85956 82607 86008 82629
rect 86008 82607 86010 82629
rect 85954 82577 85956 82583
rect 85956 82577 86008 82583
rect 86008 82577 86010 82583
rect 85954 82565 86010 82577
rect 85954 82527 85956 82565
rect 85956 82527 86008 82565
rect 86008 82527 86010 82565
rect 85954 82501 86010 82503
rect 85954 82449 85956 82501
rect 85956 82449 86008 82501
rect 86008 82449 86010 82501
rect 85954 82447 86010 82449
rect 85954 82385 85956 82423
rect 85956 82385 86008 82423
rect 86008 82385 86010 82423
rect 85954 82373 86010 82385
rect 85954 82367 85956 82373
rect 85956 82367 86008 82373
rect 86008 82367 86010 82373
rect 85954 82321 85956 82343
rect 85956 82321 86008 82343
rect 86008 82321 86010 82343
rect 85954 82309 86010 82321
rect 85954 82287 85956 82309
rect 85956 82287 86008 82309
rect 86008 82287 86010 82309
rect 85954 82257 85956 82263
rect 85956 82257 86008 82263
rect 86008 82257 86010 82263
rect 85954 82245 86010 82257
rect 85954 82207 85956 82245
rect 85956 82207 86008 82245
rect 86008 82207 86010 82245
rect 87042 82705 87044 82743
rect 87044 82705 87096 82743
rect 87096 82705 87098 82743
rect 87042 82693 87098 82705
rect 87042 82687 87044 82693
rect 87044 82687 87096 82693
rect 87096 82687 87098 82693
rect 87042 82641 87044 82663
rect 87044 82641 87096 82663
rect 87096 82641 87098 82663
rect 87042 82629 87098 82641
rect 87042 82607 87044 82629
rect 87044 82607 87096 82629
rect 87096 82607 87098 82629
rect 87042 82577 87044 82583
rect 87044 82577 87096 82583
rect 87096 82577 87098 82583
rect 87042 82565 87098 82577
rect 87042 82527 87044 82565
rect 87044 82527 87096 82565
rect 87096 82527 87098 82565
rect 87042 82501 87098 82503
rect 87042 82449 87044 82501
rect 87044 82449 87096 82501
rect 87096 82449 87098 82501
rect 87042 82447 87098 82449
rect 87042 82385 87044 82423
rect 87044 82385 87096 82423
rect 87096 82385 87098 82423
rect 87042 82373 87098 82385
rect 87042 82367 87044 82373
rect 87044 82367 87096 82373
rect 87096 82367 87098 82373
rect 87042 82321 87044 82343
rect 87044 82321 87096 82343
rect 87096 82321 87098 82343
rect 87042 82309 87098 82321
rect 87042 82287 87044 82309
rect 87044 82287 87096 82309
rect 87096 82287 87098 82309
rect 87042 82257 87044 82263
rect 87044 82257 87096 82263
rect 87096 82257 87098 82263
rect 87042 82245 87098 82257
rect 87042 82207 87044 82245
rect 87044 82207 87096 82245
rect 87096 82207 87098 82245
rect 88130 82705 88132 82743
rect 88132 82705 88184 82743
rect 88184 82705 88186 82743
rect 88130 82693 88186 82705
rect 88130 82687 88132 82693
rect 88132 82687 88184 82693
rect 88184 82687 88186 82693
rect 88130 82641 88132 82663
rect 88132 82641 88184 82663
rect 88184 82641 88186 82663
rect 88130 82629 88186 82641
rect 88130 82607 88132 82629
rect 88132 82607 88184 82629
rect 88184 82607 88186 82629
rect 88130 82577 88132 82583
rect 88132 82577 88184 82583
rect 88184 82577 88186 82583
rect 88130 82565 88186 82577
rect 88130 82527 88132 82565
rect 88132 82527 88184 82565
rect 88184 82527 88186 82565
rect 88130 82501 88186 82503
rect 88130 82449 88132 82501
rect 88132 82449 88184 82501
rect 88184 82449 88186 82501
rect 88130 82447 88186 82449
rect 88130 82385 88132 82423
rect 88132 82385 88184 82423
rect 88184 82385 88186 82423
rect 88130 82373 88186 82385
rect 88130 82367 88132 82373
rect 88132 82367 88184 82373
rect 88184 82367 88186 82373
rect 88130 82321 88132 82343
rect 88132 82321 88184 82343
rect 88184 82321 88186 82343
rect 88130 82309 88186 82321
rect 88130 82287 88132 82309
rect 88132 82287 88184 82309
rect 88184 82287 88186 82309
rect 88130 82257 88132 82263
rect 88132 82257 88184 82263
rect 88184 82257 88186 82263
rect 88130 82245 88186 82257
rect 88130 82207 88132 82245
rect 88132 82207 88184 82245
rect 88184 82207 88186 82245
rect 74529 80708 74531 80746
rect 74531 80708 74583 80746
rect 74583 80708 74585 80746
rect 74529 80696 74585 80708
rect 74529 80690 74531 80696
rect 74531 80690 74583 80696
rect 74583 80690 74585 80696
rect 74529 80644 74531 80666
rect 74531 80644 74583 80666
rect 74583 80644 74585 80666
rect 74529 80632 74585 80644
rect 74529 80610 74531 80632
rect 74531 80610 74583 80632
rect 74583 80610 74585 80632
rect 74529 80580 74531 80586
rect 74531 80580 74583 80586
rect 74583 80580 74585 80586
rect 74529 80568 74585 80580
rect 74529 80530 74531 80568
rect 74531 80530 74583 80568
rect 74583 80530 74585 80568
rect 74529 80504 74585 80506
rect 74529 80452 74531 80504
rect 74531 80452 74583 80504
rect 74583 80452 74585 80504
rect 74529 80450 74585 80452
rect 74529 80388 74531 80426
rect 74531 80388 74583 80426
rect 74583 80388 74585 80426
rect 74529 80376 74585 80388
rect 74529 80370 74531 80376
rect 74531 80370 74583 80376
rect 74583 80370 74585 80376
rect 74529 80324 74531 80346
rect 74531 80324 74583 80346
rect 74583 80324 74585 80346
rect 74529 80312 74585 80324
rect 74529 80290 74531 80312
rect 74531 80290 74583 80312
rect 74583 80290 74585 80312
rect 74529 80260 74531 80266
rect 74531 80260 74583 80266
rect 74583 80260 74585 80266
rect 74529 80248 74585 80260
rect 74529 80210 74531 80248
rect 74531 80210 74583 80248
rect 74583 80210 74585 80248
rect 75617 80708 75619 80746
rect 75619 80708 75671 80746
rect 75671 80708 75673 80746
rect 75617 80696 75673 80708
rect 75617 80690 75619 80696
rect 75619 80690 75671 80696
rect 75671 80690 75673 80696
rect 75617 80644 75619 80666
rect 75619 80644 75671 80666
rect 75671 80644 75673 80666
rect 75617 80632 75673 80644
rect 75617 80610 75619 80632
rect 75619 80610 75671 80632
rect 75671 80610 75673 80632
rect 75617 80580 75619 80586
rect 75619 80580 75671 80586
rect 75671 80580 75673 80586
rect 75617 80568 75673 80580
rect 75617 80530 75619 80568
rect 75619 80530 75671 80568
rect 75671 80530 75673 80568
rect 75617 80504 75673 80506
rect 75617 80452 75619 80504
rect 75619 80452 75671 80504
rect 75671 80452 75673 80504
rect 75617 80450 75673 80452
rect 75617 80388 75619 80426
rect 75619 80388 75671 80426
rect 75671 80388 75673 80426
rect 75617 80376 75673 80388
rect 75617 80370 75619 80376
rect 75619 80370 75671 80376
rect 75671 80370 75673 80376
rect 75617 80324 75619 80346
rect 75619 80324 75671 80346
rect 75671 80324 75673 80346
rect 75617 80312 75673 80324
rect 75617 80290 75619 80312
rect 75619 80290 75671 80312
rect 75671 80290 75673 80312
rect 75617 80260 75619 80266
rect 75619 80260 75671 80266
rect 75671 80260 75673 80266
rect 75617 80248 75673 80260
rect 75617 80210 75619 80248
rect 75619 80210 75671 80248
rect 75671 80210 75673 80248
rect 76705 80708 76707 80746
rect 76707 80708 76759 80746
rect 76759 80708 76761 80746
rect 76705 80696 76761 80708
rect 76705 80690 76707 80696
rect 76707 80690 76759 80696
rect 76759 80690 76761 80696
rect 76705 80644 76707 80666
rect 76707 80644 76759 80666
rect 76759 80644 76761 80666
rect 76705 80632 76761 80644
rect 76705 80610 76707 80632
rect 76707 80610 76759 80632
rect 76759 80610 76761 80632
rect 76705 80580 76707 80586
rect 76707 80580 76759 80586
rect 76759 80580 76761 80586
rect 76705 80568 76761 80580
rect 76705 80530 76707 80568
rect 76707 80530 76759 80568
rect 76759 80530 76761 80568
rect 76705 80504 76761 80506
rect 76705 80452 76707 80504
rect 76707 80452 76759 80504
rect 76759 80452 76761 80504
rect 76705 80450 76761 80452
rect 76705 80388 76707 80426
rect 76707 80388 76759 80426
rect 76759 80388 76761 80426
rect 76705 80376 76761 80388
rect 76705 80370 76707 80376
rect 76707 80370 76759 80376
rect 76759 80370 76761 80376
rect 76705 80324 76707 80346
rect 76707 80324 76759 80346
rect 76759 80324 76761 80346
rect 76705 80312 76761 80324
rect 76705 80290 76707 80312
rect 76707 80290 76759 80312
rect 76759 80290 76761 80312
rect 76705 80260 76707 80266
rect 76707 80260 76759 80266
rect 76759 80260 76761 80266
rect 76705 80248 76761 80260
rect 76705 80210 76707 80248
rect 76707 80210 76759 80248
rect 76759 80210 76761 80248
rect 77793 80708 77795 80746
rect 77795 80708 77847 80746
rect 77847 80708 77849 80746
rect 77793 80696 77849 80708
rect 77793 80690 77795 80696
rect 77795 80690 77847 80696
rect 77847 80690 77849 80696
rect 77793 80644 77795 80666
rect 77795 80644 77847 80666
rect 77847 80644 77849 80666
rect 77793 80632 77849 80644
rect 77793 80610 77795 80632
rect 77795 80610 77847 80632
rect 77847 80610 77849 80632
rect 77793 80580 77795 80586
rect 77795 80580 77847 80586
rect 77847 80580 77849 80586
rect 77793 80568 77849 80580
rect 77793 80530 77795 80568
rect 77795 80530 77847 80568
rect 77847 80530 77849 80568
rect 77793 80504 77849 80506
rect 77793 80452 77795 80504
rect 77795 80452 77847 80504
rect 77847 80452 77849 80504
rect 77793 80450 77849 80452
rect 77793 80388 77795 80426
rect 77795 80388 77847 80426
rect 77847 80388 77849 80426
rect 77793 80376 77849 80388
rect 77793 80370 77795 80376
rect 77795 80370 77847 80376
rect 77847 80370 77849 80376
rect 77793 80324 77795 80346
rect 77795 80324 77847 80346
rect 77847 80324 77849 80346
rect 77793 80312 77849 80324
rect 77793 80290 77795 80312
rect 77795 80290 77847 80312
rect 77847 80290 77849 80312
rect 77793 80260 77795 80266
rect 77795 80260 77847 80266
rect 77847 80260 77849 80266
rect 77793 80248 77849 80260
rect 77793 80210 77795 80248
rect 77795 80210 77847 80248
rect 77847 80210 77849 80248
rect 78881 80708 78883 80746
rect 78883 80708 78935 80746
rect 78935 80708 78937 80746
rect 78881 80696 78937 80708
rect 78881 80690 78883 80696
rect 78883 80690 78935 80696
rect 78935 80690 78937 80696
rect 78881 80644 78883 80666
rect 78883 80644 78935 80666
rect 78935 80644 78937 80666
rect 78881 80632 78937 80644
rect 78881 80610 78883 80632
rect 78883 80610 78935 80632
rect 78935 80610 78937 80632
rect 78881 80580 78883 80586
rect 78883 80580 78935 80586
rect 78935 80580 78937 80586
rect 78881 80568 78937 80580
rect 78881 80530 78883 80568
rect 78883 80530 78935 80568
rect 78935 80530 78937 80568
rect 78881 80504 78937 80506
rect 78881 80452 78883 80504
rect 78883 80452 78935 80504
rect 78935 80452 78937 80504
rect 78881 80450 78937 80452
rect 78881 80388 78883 80426
rect 78883 80388 78935 80426
rect 78935 80388 78937 80426
rect 78881 80376 78937 80388
rect 78881 80370 78883 80376
rect 78883 80370 78935 80376
rect 78935 80370 78937 80376
rect 78881 80324 78883 80346
rect 78883 80324 78935 80346
rect 78935 80324 78937 80346
rect 78881 80312 78937 80324
rect 78881 80290 78883 80312
rect 78883 80290 78935 80312
rect 78935 80290 78937 80312
rect 78881 80260 78883 80266
rect 78883 80260 78935 80266
rect 78935 80260 78937 80266
rect 78881 80248 78937 80260
rect 78881 80210 78883 80248
rect 78883 80210 78935 80248
rect 78935 80210 78937 80248
rect 79969 80708 79971 80746
rect 79971 80708 80023 80746
rect 80023 80708 80025 80746
rect 79969 80696 80025 80708
rect 79969 80690 79971 80696
rect 79971 80690 80023 80696
rect 80023 80690 80025 80696
rect 79969 80644 79971 80666
rect 79971 80644 80023 80666
rect 80023 80644 80025 80666
rect 79969 80632 80025 80644
rect 79969 80610 79971 80632
rect 79971 80610 80023 80632
rect 80023 80610 80025 80632
rect 79969 80580 79971 80586
rect 79971 80580 80023 80586
rect 80023 80580 80025 80586
rect 79969 80568 80025 80580
rect 79969 80530 79971 80568
rect 79971 80530 80023 80568
rect 80023 80530 80025 80568
rect 79969 80504 80025 80506
rect 79969 80452 79971 80504
rect 79971 80452 80023 80504
rect 80023 80452 80025 80504
rect 79969 80450 80025 80452
rect 79969 80388 79971 80426
rect 79971 80388 80023 80426
rect 80023 80388 80025 80426
rect 79969 80376 80025 80388
rect 79969 80370 79971 80376
rect 79971 80370 80023 80376
rect 80023 80370 80025 80376
rect 79969 80324 79971 80346
rect 79971 80324 80023 80346
rect 80023 80324 80025 80346
rect 79969 80312 80025 80324
rect 79969 80290 79971 80312
rect 79971 80290 80023 80312
rect 80023 80290 80025 80312
rect 79969 80260 79971 80266
rect 79971 80260 80023 80266
rect 80023 80260 80025 80266
rect 79969 80248 80025 80260
rect 79969 80210 79971 80248
rect 79971 80210 80023 80248
rect 80023 80210 80025 80248
rect 81057 80708 81059 80746
rect 81059 80708 81111 80746
rect 81111 80708 81113 80746
rect 81057 80696 81113 80708
rect 81057 80690 81059 80696
rect 81059 80690 81111 80696
rect 81111 80690 81113 80696
rect 81057 80644 81059 80666
rect 81059 80644 81111 80666
rect 81111 80644 81113 80666
rect 81057 80632 81113 80644
rect 81057 80610 81059 80632
rect 81059 80610 81111 80632
rect 81111 80610 81113 80632
rect 81057 80580 81059 80586
rect 81059 80580 81111 80586
rect 81111 80580 81113 80586
rect 81057 80568 81113 80580
rect 81057 80530 81059 80568
rect 81059 80530 81111 80568
rect 81111 80530 81113 80568
rect 81057 80504 81113 80506
rect 81057 80452 81059 80504
rect 81059 80452 81111 80504
rect 81111 80452 81113 80504
rect 81057 80450 81113 80452
rect 81057 80388 81059 80426
rect 81059 80388 81111 80426
rect 81111 80388 81113 80426
rect 81057 80376 81113 80388
rect 81057 80370 81059 80376
rect 81059 80370 81111 80376
rect 81111 80370 81113 80376
rect 81057 80324 81059 80346
rect 81059 80324 81111 80346
rect 81111 80324 81113 80346
rect 81057 80312 81113 80324
rect 81057 80290 81059 80312
rect 81059 80290 81111 80312
rect 81111 80290 81113 80312
rect 81057 80260 81059 80266
rect 81059 80260 81111 80266
rect 81111 80260 81113 80266
rect 81057 80248 81113 80260
rect 81057 80210 81059 80248
rect 81059 80210 81111 80248
rect 81111 80210 81113 80248
rect 82145 80708 82147 80746
rect 82147 80708 82199 80746
rect 82199 80708 82201 80746
rect 82145 80696 82201 80708
rect 82145 80690 82147 80696
rect 82147 80690 82199 80696
rect 82199 80690 82201 80696
rect 82145 80644 82147 80666
rect 82147 80644 82199 80666
rect 82199 80644 82201 80666
rect 82145 80632 82201 80644
rect 82145 80610 82147 80632
rect 82147 80610 82199 80632
rect 82199 80610 82201 80632
rect 82145 80580 82147 80586
rect 82147 80580 82199 80586
rect 82199 80580 82201 80586
rect 82145 80568 82201 80580
rect 82145 80530 82147 80568
rect 82147 80530 82199 80568
rect 82199 80530 82201 80568
rect 82145 80504 82201 80506
rect 82145 80452 82147 80504
rect 82147 80452 82199 80504
rect 82199 80452 82201 80504
rect 82145 80450 82201 80452
rect 82145 80388 82147 80426
rect 82147 80388 82199 80426
rect 82199 80388 82201 80426
rect 82145 80376 82201 80388
rect 82145 80370 82147 80376
rect 82147 80370 82199 80376
rect 82199 80370 82201 80376
rect 82145 80324 82147 80346
rect 82147 80324 82199 80346
rect 82199 80324 82201 80346
rect 82145 80312 82201 80324
rect 82145 80290 82147 80312
rect 82147 80290 82199 80312
rect 82199 80290 82201 80312
rect 82145 80260 82147 80266
rect 82147 80260 82199 80266
rect 82199 80260 82201 80266
rect 82145 80248 82201 80260
rect 82145 80210 82147 80248
rect 82147 80210 82199 80248
rect 82199 80210 82201 80248
rect 83233 80708 83235 80746
rect 83235 80708 83287 80746
rect 83287 80708 83289 80746
rect 83233 80696 83289 80708
rect 83233 80690 83235 80696
rect 83235 80690 83287 80696
rect 83287 80690 83289 80696
rect 83233 80644 83235 80666
rect 83235 80644 83287 80666
rect 83287 80644 83289 80666
rect 83233 80632 83289 80644
rect 83233 80610 83235 80632
rect 83235 80610 83287 80632
rect 83287 80610 83289 80632
rect 83233 80580 83235 80586
rect 83235 80580 83287 80586
rect 83287 80580 83289 80586
rect 83233 80568 83289 80580
rect 83233 80530 83235 80568
rect 83235 80530 83287 80568
rect 83287 80530 83289 80568
rect 83233 80504 83289 80506
rect 83233 80452 83235 80504
rect 83235 80452 83287 80504
rect 83287 80452 83289 80504
rect 83233 80450 83289 80452
rect 83233 80388 83235 80426
rect 83235 80388 83287 80426
rect 83287 80388 83289 80426
rect 83233 80376 83289 80388
rect 83233 80370 83235 80376
rect 83235 80370 83287 80376
rect 83287 80370 83289 80376
rect 83233 80324 83235 80346
rect 83235 80324 83287 80346
rect 83287 80324 83289 80346
rect 83233 80312 83289 80324
rect 83233 80290 83235 80312
rect 83235 80290 83287 80312
rect 83287 80290 83289 80312
rect 83233 80260 83235 80266
rect 83235 80260 83287 80266
rect 83287 80260 83289 80266
rect 83233 80248 83289 80260
rect 83233 80210 83235 80248
rect 83235 80210 83287 80248
rect 83287 80210 83289 80248
rect 84321 80708 84323 80746
rect 84323 80708 84375 80746
rect 84375 80708 84377 80746
rect 84321 80696 84377 80708
rect 84321 80690 84323 80696
rect 84323 80690 84375 80696
rect 84375 80690 84377 80696
rect 84321 80644 84323 80666
rect 84323 80644 84375 80666
rect 84375 80644 84377 80666
rect 84321 80632 84377 80644
rect 84321 80610 84323 80632
rect 84323 80610 84375 80632
rect 84375 80610 84377 80632
rect 84321 80580 84323 80586
rect 84323 80580 84375 80586
rect 84375 80580 84377 80586
rect 84321 80568 84377 80580
rect 84321 80530 84323 80568
rect 84323 80530 84375 80568
rect 84375 80530 84377 80568
rect 84321 80504 84377 80506
rect 84321 80452 84323 80504
rect 84323 80452 84375 80504
rect 84375 80452 84377 80504
rect 84321 80450 84377 80452
rect 84321 80388 84323 80426
rect 84323 80388 84375 80426
rect 84375 80388 84377 80426
rect 84321 80376 84377 80388
rect 84321 80370 84323 80376
rect 84323 80370 84375 80376
rect 84375 80370 84377 80376
rect 84321 80324 84323 80346
rect 84323 80324 84375 80346
rect 84375 80324 84377 80346
rect 84321 80312 84377 80324
rect 84321 80290 84323 80312
rect 84323 80290 84375 80312
rect 84375 80290 84377 80312
rect 84321 80260 84323 80266
rect 84323 80260 84375 80266
rect 84375 80260 84377 80266
rect 84321 80248 84377 80260
rect 84321 80210 84323 80248
rect 84323 80210 84375 80248
rect 84375 80210 84377 80248
rect 85409 80708 85411 80746
rect 85411 80708 85463 80746
rect 85463 80708 85465 80746
rect 85409 80696 85465 80708
rect 85409 80690 85411 80696
rect 85411 80690 85463 80696
rect 85463 80690 85465 80696
rect 85409 80644 85411 80666
rect 85411 80644 85463 80666
rect 85463 80644 85465 80666
rect 85409 80632 85465 80644
rect 85409 80610 85411 80632
rect 85411 80610 85463 80632
rect 85463 80610 85465 80632
rect 85409 80580 85411 80586
rect 85411 80580 85463 80586
rect 85463 80580 85465 80586
rect 85409 80568 85465 80580
rect 85409 80530 85411 80568
rect 85411 80530 85463 80568
rect 85463 80530 85465 80568
rect 85409 80504 85465 80506
rect 85409 80452 85411 80504
rect 85411 80452 85463 80504
rect 85463 80452 85465 80504
rect 85409 80450 85465 80452
rect 85409 80388 85411 80426
rect 85411 80388 85463 80426
rect 85463 80388 85465 80426
rect 85409 80376 85465 80388
rect 85409 80370 85411 80376
rect 85411 80370 85463 80376
rect 85463 80370 85465 80376
rect 85409 80324 85411 80346
rect 85411 80324 85463 80346
rect 85463 80324 85465 80346
rect 85409 80312 85465 80324
rect 85409 80290 85411 80312
rect 85411 80290 85463 80312
rect 85463 80290 85465 80312
rect 85409 80260 85411 80266
rect 85411 80260 85463 80266
rect 85463 80260 85465 80266
rect 85409 80248 85465 80260
rect 85409 80210 85411 80248
rect 85411 80210 85463 80248
rect 85463 80210 85465 80248
rect 86497 80708 86499 80746
rect 86499 80708 86551 80746
rect 86551 80708 86553 80746
rect 86497 80696 86553 80708
rect 86497 80690 86499 80696
rect 86499 80690 86551 80696
rect 86551 80690 86553 80696
rect 86497 80644 86499 80666
rect 86499 80644 86551 80666
rect 86551 80644 86553 80666
rect 86497 80632 86553 80644
rect 86497 80610 86499 80632
rect 86499 80610 86551 80632
rect 86551 80610 86553 80632
rect 86497 80580 86499 80586
rect 86499 80580 86551 80586
rect 86551 80580 86553 80586
rect 86497 80568 86553 80580
rect 86497 80530 86499 80568
rect 86499 80530 86551 80568
rect 86551 80530 86553 80568
rect 86497 80504 86553 80506
rect 86497 80452 86499 80504
rect 86499 80452 86551 80504
rect 86551 80452 86553 80504
rect 86497 80450 86553 80452
rect 86497 80388 86499 80426
rect 86499 80388 86551 80426
rect 86551 80388 86553 80426
rect 86497 80376 86553 80388
rect 86497 80370 86499 80376
rect 86499 80370 86551 80376
rect 86551 80370 86553 80376
rect 86497 80324 86499 80346
rect 86499 80324 86551 80346
rect 86551 80324 86553 80346
rect 86497 80312 86553 80324
rect 86497 80290 86499 80312
rect 86499 80290 86551 80312
rect 86551 80290 86553 80312
rect 86497 80260 86499 80266
rect 86499 80260 86551 80266
rect 86551 80260 86553 80266
rect 86497 80248 86553 80260
rect 86497 80210 86499 80248
rect 86499 80210 86551 80248
rect 86551 80210 86553 80248
rect 87585 80708 87587 80746
rect 87587 80708 87639 80746
rect 87639 80708 87641 80746
rect 87585 80696 87641 80708
rect 87585 80690 87587 80696
rect 87587 80690 87639 80696
rect 87639 80690 87641 80696
rect 87585 80644 87587 80666
rect 87587 80644 87639 80666
rect 87639 80644 87641 80666
rect 87585 80632 87641 80644
rect 87585 80610 87587 80632
rect 87587 80610 87639 80632
rect 87639 80610 87641 80632
rect 87585 80580 87587 80586
rect 87587 80580 87639 80586
rect 87639 80580 87641 80586
rect 87585 80568 87641 80580
rect 87585 80530 87587 80568
rect 87587 80530 87639 80568
rect 87639 80530 87641 80568
rect 87585 80504 87641 80506
rect 87585 80452 87587 80504
rect 87587 80452 87639 80504
rect 87639 80452 87641 80504
rect 87585 80450 87641 80452
rect 87585 80388 87587 80426
rect 87587 80388 87639 80426
rect 87639 80388 87641 80426
rect 87585 80376 87641 80388
rect 87585 80370 87587 80376
rect 87587 80370 87639 80376
rect 87639 80370 87641 80376
rect 87585 80324 87587 80346
rect 87587 80324 87639 80346
rect 87639 80324 87641 80346
rect 87585 80312 87641 80324
rect 87585 80290 87587 80312
rect 87587 80290 87639 80312
rect 87639 80290 87641 80312
rect 87585 80260 87587 80266
rect 87587 80260 87639 80266
rect 87639 80260 87641 80266
rect 87585 80248 87641 80260
rect 87585 80210 87587 80248
rect 87587 80210 87639 80248
rect 87639 80210 87641 80248
rect 88673 80708 88675 80746
rect 88675 80708 88727 80746
rect 88727 80708 88729 80746
rect 88673 80696 88729 80708
rect 88673 80690 88675 80696
rect 88675 80690 88727 80696
rect 88727 80690 88729 80696
rect 88673 80644 88675 80666
rect 88675 80644 88727 80666
rect 88727 80644 88729 80666
rect 88673 80632 88729 80644
rect 88673 80610 88675 80632
rect 88675 80610 88727 80632
rect 88727 80610 88729 80632
rect 88673 80580 88675 80586
rect 88675 80580 88727 80586
rect 88727 80580 88729 80586
rect 88673 80568 88729 80580
rect 88673 80530 88675 80568
rect 88675 80530 88727 80568
rect 88727 80530 88729 80568
rect 88673 80504 88729 80506
rect 88673 80452 88675 80504
rect 88675 80452 88727 80504
rect 88727 80452 88729 80504
rect 88673 80450 88729 80452
rect 88673 80388 88675 80426
rect 88675 80388 88727 80426
rect 88727 80388 88729 80426
rect 88673 80376 88729 80388
rect 88673 80370 88675 80376
rect 88675 80370 88727 80376
rect 88727 80370 88729 80376
rect 88673 80324 88675 80346
rect 88675 80324 88727 80346
rect 88727 80324 88729 80346
rect 88673 80312 88729 80324
rect 88673 80290 88675 80312
rect 88675 80290 88727 80312
rect 88727 80290 88729 80312
rect 88673 80260 88675 80266
rect 88675 80260 88727 80266
rect 88727 80260 88729 80266
rect 88673 80248 88729 80260
rect 88673 80210 88675 80248
rect 88675 80210 88727 80248
rect 88727 80210 88729 80248
rect 75074 78705 75076 78743
rect 75076 78705 75128 78743
rect 75128 78705 75130 78743
rect 75074 78693 75130 78705
rect 75074 78687 75076 78693
rect 75076 78687 75128 78693
rect 75128 78687 75130 78693
rect 75074 78641 75076 78663
rect 75076 78641 75128 78663
rect 75128 78641 75130 78663
rect 75074 78629 75130 78641
rect 75074 78607 75076 78629
rect 75076 78607 75128 78629
rect 75128 78607 75130 78629
rect 75074 78577 75076 78583
rect 75076 78577 75128 78583
rect 75128 78577 75130 78583
rect 75074 78565 75130 78577
rect 75074 78527 75076 78565
rect 75076 78527 75128 78565
rect 75128 78527 75130 78565
rect 75074 78501 75130 78503
rect 75074 78449 75076 78501
rect 75076 78449 75128 78501
rect 75128 78449 75130 78501
rect 75074 78447 75130 78449
rect 75074 78385 75076 78423
rect 75076 78385 75128 78423
rect 75128 78385 75130 78423
rect 75074 78373 75130 78385
rect 75074 78367 75076 78373
rect 75076 78367 75128 78373
rect 75128 78367 75130 78373
rect 75074 78321 75076 78343
rect 75076 78321 75128 78343
rect 75128 78321 75130 78343
rect 75074 78309 75130 78321
rect 75074 78287 75076 78309
rect 75076 78287 75128 78309
rect 75128 78287 75130 78309
rect 75074 78257 75076 78263
rect 75076 78257 75128 78263
rect 75128 78257 75130 78263
rect 75074 78245 75130 78257
rect 75074 78207 75076 78245
rect 75076 78207 75128 78245
rect 75128 78207 75130 78245
rect 76162 78705 76164 78743
rect 76164 78705 76216 78743
rect 76216 78705 76218 78743
rect 76162 78693 76218 78705
rect 76162 78687 76164 78693
rect 76164 78687 76216 78693
rect 76216 78687 76218 78693
rect 76162 78641 76164 78663
rect 76164 78641 76216 78663
rect 76216 78641 76218 78663
rect 76162 78629 76218 78641
rect 76162 78607 76164 78629
rect 76164 78607 76216 78629
rect 76216 78607 76218 78629
rect 76162 78577 76164 78583
rect 76164 78577 76216 78583
rect 76216 78577 76218 78583
rect 76162 78565 76218 78577
rect 76162 78527 76164 78565
rect 76164 78527 76216 78565
rect 76216 78527 76218 78565
rect 76162 78501 76218 78503
rect 76162 78449 76164 78501
rect 76164 78449 76216 78501
rect 76216 78449 76218 78501
rect 76162 78447 76218 78449
rect 76162 78385 76164 78423
rect 76164 78385 76216 78423
rect 76216 78385 76218 78423
rect 76162 78373 76218 78385
rect 76162 78367 76164 78373
rect 76164 78367 76216 78373
rect 76216 78367 76218 78373
rect 76162 78321 76164 78343
rect 76164 78321 76216 78343
rect 76216 78321 76218 78343
rect 76162 78309 76218 78321
rect 76162 78287 76164 78309
rect 76164 78287 76216 78309
rect 76216 78287 76218 78309
rect 76162 78257 76164 78263
rect 76164 78257 76216 78263
rect 76216 78257 76218 78263
rect 76162 78245 76218 78257
rect 76162 78207 76164 78245
rect 76164 78207 76216 78245
rect 76216 78207 76218 78245
rect 77250 78705 77252 78743
rect 77252 78705 77304 78743
rect 77304 78705 77306 78743
rect 77250 78693 77306 78705
rect 77250 78687 77252 78693
rect 77252 78687 77304 78693
rect 77304 78687 77306 78693
rect 77250 78641 77252 78663
rect 77252 78641 77304 78663
rect 77304 78641 77306 78663
rect 77250 78629 77306 78641
rect 77250 78607 77252 78629
rect 77252 78607 77304 78629
rect 77304 78607 77306 78629
rect 77250 78577 77252 78583
rect 77252 78577 77304 78583
rect 77304 78577 77306 78583
rect 77250 78565 77306 78577
rect 77250 78527 77252 78565
rect 77252 78527 77304 78565
rect 77304 78527 77306 78565
rect 77250 78501 77306 78503
rect 77250 78449 77252 78501
rect 77252 78449 77304 78501
rect 77304 78449 77306 78501
rect 77250 78447 77306 78449
rect 77250 78385 77252 78423
rect 77252 78385 77304 78423
rect 77304 78385 77306 78423
rect 77250 78373 77306 78385
rect 77250 78367 77252 78373
rect 77252 78367 77304 78373
rect 77304 78367 77306 78373
rect 77250 78321 77252 78343
rect 77252 78321 77304 78343
rect 77304 78321 77306 78343
rect 77250 78309 77306 78321
rect 77250 78287 77252 78309
rect 77252 78287 77304 78309
rect 77304 78287 77306 78309
rect 77250 78257 77252 78263
rect 77252 78257 77304 78263
rect 77304 78257 77306 78263
rect 77250 78245 77306 78257
rect 77250 78207 77252 78245
rect 77252 78207 77304 78245
rect 77304 78207 77306 78245
rect 78338 78705 78340 78743
rect 78340 78705 78392 78743
rect 78392 78705 78394 78743
rect 78338 78693 78394 78705
rect 78338 78687 78340 78693
rect 78340 78687 78392 78693
rect 78392 78687 78394 78693
rect 78338 78641 78340 78663
rect 78340 78641 78392 78663
rect 78392 78641 78394 78663
rect 78338 78629 78394 78641
rect 78338 78607 78340 78629
rect 78340 78607 78392 78629
rect 78392 78607 78394 78629
rect 78338 78577 78340 78583
rect 78340 78577 78392 78583
rect 78392 78577 78394 78583
rect 78338 78565 78394 78577
rect 78338 78527 78340 78565
rect 78340 78527 78392 78565
rect 78392 78527 78394 78565
rect 78338 78501 78394 78503
rect 78338 78449 78340 78501
rect 78340 78449 78392 78501
rect 78392 78449 78394 78501
rect 78338 78447 78394 78449
rect 78338 78385 78340 78423
rect 78340 78385 78392 78423
rect 78392 78385 78394 78423
rect 78338 78373 78394 78385
rect 78338 78367 78340 78373
rect 78340 78367 78392 78373
rect 78392 78367 78394 78373
rect 78338 78321 78340 78343
rect 78340 78321 78392 78343
rect 78392 78321 78394 78343
rect 78338 78309 78394 78321
rect 78338 78287 78340 78309
rect 78340 78287 78392 78309
rect 78392 78287 78394 78309
rect 78338 78257 78340 78263
rect 78340 78257 78392 78263
rect 78392 78257 78394 78263
rect 78338 78245 78394 78257
rect 78338 78207 78340 78245
rect 78340 78207 78392 78245
rect 78392 78207 78394 78245
rect 79426 78705 79428 78743
rect 79428 78705 79480 78743
rect 79480 78705 79482 78743
rect 79426 78693 79482 78705
rect 79426 78687 79428 78693
rect 79428 78687 79480 78693
rect 79480 78687 79482 78693
rect 79426 78641 79428 78663
rect 79428 78641 79480 78663
rect 79480 78641 79482 78663
rect 79426 78629 79482 78641
rect 79426 78607 79428 78629
rect 79428 78607 79480 78629
rect 79480 78607 79482 78629
rect 79426 78577 79428 78583
rect 79428 78577 79480 78583
rect 79480 78577 79482 78583
rect 79426 78565 79482 78577
rect 79426 78527 79428 78565
rect 79428 78527 79480 78565
rect 79480 78527 79482 78565
rect 79426 78501 79482 78503
rect 79426 78449 79428 78501
rect 79428 78449 79480 78501
rect 79480 78449 79482 78501
rect 79426 78447 79482 78449
rect 79426 78385 79428 78423
rect 79428 78385 79480 78423
rect 79480 78385 79482 78423
rect 79426 78373 79482 78385
rect 79426 78367 79428 78373
rect 79428 78367 79480 78373
rect 79480 78367 79482 78373
rect 79426 78321 79428 78343
rect 79428 78321 79480 78343
rect 79480 78321 79482 78343
rect 79426 78309 79482 78321
rect 79426 78287 79428 78309
rect 79428 78287 79480 78309
rect 79480 78287 79482 78309
rect 79426 78257 79428 78263
rect 79428 78257 79480 78263
rect 79480 78257 79482 78263
rect 79426 78245 79482 78257
rect 79426 78207 79428 78245
rect 79428 78207 79480 78245
rect 79480 78207 79482 78245
rect 80514 78705 80516 78743
rect 80516 78705 80568 78743
rect 80568 78705 80570 78743
rect 80514 78693 80570 78705
rect 80514 78687 80516 78693
rect 80516 78687 80568 78693
rect 80568 78687 80570 78693
rect 80514 78641 80516 78663
rect 80516 78641 80568 78663
rect 80568 78641 80570 78663
rect 80514 78629 80570 78641
rect 80514 78607 80516 78629
rect 80516 78607 80568 78629
rect 80568 78607 80570 78629
rect 80514 78577 80516 78583
rect 80516 78577 80568 78583
rect 80568 78577 80570 78583
rect 80514 78565 80570 78577
rect 80514 78527 80516 78565
rect 80516 78527 80568 78565
rect 80568 78527 80570 78565
rect 80514 78501 80570 78503
rect 80514 78449 80516 78501
rect 80516 78449 80568 78501
rect 80568 78449 80570 78501
rect 80514 78447 80570 78449
rect 80514 78385 80516 78423
rect 80516 78385 80568 78423
rect 80568 78385 80570 78423
rect 80514 78373 80570 78385
rect 80514 78367 80516 78373
rect 80516 78367 80568 78373
rect 80568 78367 80570 78373
rect 80514 78321 80516 78343
rect 80516 78321 80568 78343
rect 80568 78321 80570 78343
rect 80514 78309 80570 78321
rect 80514 78287 80516 78309
rect 80516 78287 80568 78309
rect 80568 78287 80570 78309
rect 80514 78257 80516 78263
rect 80516 78257 80568 78263
rect 80568 78257 80570 78263
rect 80514 78245 80570 78257
rect 80514 78207 80516 78245
rect 80516 78207 80568 78245
rect 80568 78207 80570 78245
rect 81602 78705 81604 78743
rect 81604 78705 81656 78743
rect 81656 78705 81658 78743
rect 81602 78693 81658 78705
rect 81602 78687 81604 78693
rect 81604 78687 81656 78693
rect 81656 78687 81658 78693
rect 81602 78641 81604 78663
rect 81604 78641 81656 78663
rect 81656 78641 81658 78663
rect 81602 78629 81658 78641
rect 81602 78607 81604 78629
rect 81604 78607 81656 78629
rect 81656 78607 81658 78629
rect 81602 78577 81604 78583
rect 81604 78577 81656 78583
rect 81656 78577 81658 78583
rect 81602 78565 81658 78577
rect 81602 78527 81604 78565
rect 81604 78527 81656 78565
rect 81656 78527 81658 78565
rect 81602 78501 81658 78503
rect 81602 78449 81604 78501
rect 81604 78449 81656 78501
rect 81656 78449 81658 78501
rect 81602 78447 81658 78449
rect 81602 78385 81604 78423
rect 81604 78385 81656 78423
rect 81656 78385 81658 78423
rect 81602 78373 81658 78385
rect 81602 78367 81604 78373
rect 81604 78367 81656 78373
rect 81656 78367 81658 78373
rect 81602 78321 81604 78343
rect 81604 78321 81656 78343
rect 81656 78321 81658 78343
rect 81602 78309 81658 78321
rect 81602 78287 81604 78309
rect 81604 78287 81656 78309
rect 81656 78287 81658 78309
rect 81602 78257 81604 78263
rect 81604 78257 81656 78263
rect 81656 78257 81658 78263
rect 81602 78245 81658 78257
rect 81602 78207 81604 78245
rect 81604 78207 81656 78245
rect 81656 78207 81658 78245
rect 82690 78705 82692 78743
rect 82692 78705 82744 78743
rect 82744 78705 82746 78743
rect 82690 78693 82746 78705
rect 82690 78687 82692 78693
rect 82692 78687 82744 78693
rect 82744 78687 82746 78693
rect 82690 78641 82692 78663
rect 82692 78641 82744 78663
rect 82744 78641 82746 78663
rect 82690 78629 82746 78641
rect 82690 78607 82692 78629
rect 82692 78607 82744 78629
rect 82744 78607 82746 78629
rect 82690 78577 82692 78583
rect 82692 78577 82744 78583
rect 82744 78577 82746 78583
rect 82690 78565 82746 78577
rect 82690 78527 82692 78565
rect 82692 78527 82744 78565
rect 82744 78527 82746 78565
rect 82690 78501 82746 78503
rect 82690 78449 82692 78501
rect 82692 78449 82744 78501
rect 82744 78449 82746 78501
rect 82690 78447 82746 78449
rect 82690 78385 82692 78423
rect 82692 78385 82744 78423
rect 82744 78385 82746 78423
rect 82690 78373 82746 78385
rect 82690 78367 82692 78373
rect 82692 78367 82744 78373
rect 82744 78367 82746 78373
rect 82690 78321 82692 78343
rect 82692 78321 82744 78343
rect 82744 78321 82746 78343
rect 82690 78309 82746 78321
rect 82690 78287 82692 78309
rect 82692 78287 82744 78309
rect 82744 78287 82746 78309
rect 82690 78257 82692 78263
rect 82692 78257 82744 78263
rect 82744 78257 82746 78263
rect 82690 78245 82746 78257
rect 82690 78207 82692 78245
rect 82692 78207 82744 78245
rect 82744 78207 82746 78245
rect 83778 78705 83780 78743
rect 83780 78705 83832 78743
rect 83832 78705 83834 78743
rect 83778 78693 83834 78705
rect 83778 78687 83780 78693
rect 83780 78687 83832 78693
rect 83832 78687 83834 78693
rect 83778 78641 83780 78663
rect 83780 78641 83832 78663
rect 83832 78641 83834 78663
rect 83778 78629 83834 78641
rect 83778 78607 83780 78629
rect 83780 78607 83832 78629
rect 83832 78607 83834 78629
rect 83778 78577 83780 78583
rect 83780 78577 83832 78583
rect 83832 78577 83834 78583
rect 83778 78565 83834 78577
rect 83778 78527 83780 78565
rect 83780 78527 83832 78565
rect 83832 78527 83834 78565
rect 83778 78501 83834 78503
rect 83778 78449 83780 78501
rect 83780 78449 83832 78501
rect 83832 78449 83834 78501
rect 83778 78447 83834 78449
rect 83778 78385 83780 78423
rect 83780 78385 83832 78423
rect 83832 78385 83834 78423
rect 83778 78373 83834 78385
rect 83778 78367 83780 78373
rect 83780 78367 83832 78373
rect 83832 78367 83834 78373
rect 83778 78321 83780 78343
rect 83780 78321 83832 78343
rect 83832 78321 83834 78343
rect 83778 78309 83834 78321
rect 83778 78287 83780 78309
rect 83780 78287 83832 78309
rect 83832 78287 83834 78309
rect 83778 78257 83780 78263
rect 83780 78257 83832 78263
rect 83832 78257 83834 78263
rect 83778 78245 83834 78257
rect 83778 78207 83780 78245
rect 83780 78207 83832 78245
rect 83832 78207 83834 78245
rect 84866 78705 84868 78743
rect 84868 78705 84920 78743
rect 84920 78705 84922 78743
rect 84866 78693 84922 78705
rect 84866 78687 84868 78693
rect 84868 78687 84920 78693
rect 84920 78687 84922 78693
rect 84866 78641 84868 78663
rect 84868 78641 84920 78663
rect 84920 78641 84922 78663
rect 84866 78629 84922 78641
rect 84866 78607 84868 78629
rect 84868 78607 84920 78629
rect 84920 78607 84922 78629
rect 84866 78577 84868 78583
rect 84868 78577 84920 78583
rect 84920 78577 84922 78583
rect 84866 78565 84922 78577
rect 84866 78527 84868 78565
rect 84868 78527 84920 78565
rect 84920 78527 84922 78565
rect 84866 78501 84922 78503
rect 84866 78449 84868 78501
rect 84868 78449 84920 78501
rect 84920 78449 84922 78501
rect 84866 78447 84922 78449
rect 84866 78385 84868 78423
rect 84868 78385 84920 78423
rect 84920 78385 84922 78423
rect 84866 78373 84922 78385
rect 84866 78367 84868 78373
rect 84868 78367 84920 78373
rect 84920 78367 84922 78373
rect 84866 78321 84868 78343
rect 84868 78321 84920 78343
rect 84920 78321 84922 78343
rect 84866 78309 84922 78321
rect 84866 78287 84868 78309
rect 84868 78287 84920 78309
rect 84920 78287 84922 78309
rect 84866 78257 84868 78263
rect 84868 78257 84920 78263
rect 84920 78257 84922 78263
rect 84866 78245 84922 78257
rect 84866 78207 84868 78245
rect 84868 78207 84920 78245
rect 84920 78207 84922 78245
rect 85954 78705 85956 78743
rect 85956 78705 86008 78743
rect 86008 78705 86010 78743
rect 85954 78693 86010 78705
rect 85954 78687 85956 78693
rect 85956 78687 86008 78693
rect 86008 78687 86010 78693
rect 85954 78641 85956 78663
rect 85956 78641 86008 78663
rect 86008 78641 86010 78663
rect 85954 78629 86010 78641
rect 85954 78607 85956 78629
rect 85956 78607 86008 78629
rect 86008 78607 86010 78629
rect 85954 78577 85956 78583
rect 85956 78577 86008 78583
rect 86008 78577 86010 78583
rect 85954 78565 86010 78577
rect 85954 78527 85956 78565
rect 85956 78527 86008 78565
rect 86008 78527 86010 78565
rect 85954 78501 86010 78503
rect 85954 78449 85956 78501
rect 85956 78449 86008 78501
rect 86008 78449 86010 78501
rect 85954 78447 86010 78449
rect 85954 78385 85956 78423
rect 85956 78385 86008 78423
rect 86008 78385 86010 78423
rect 85954 78373 86010 78385
rect 85954 78367 85956 78373
rect 85956 78367 86008 78373
rect 86008 78367 86010 78373
rect 85954 78321 85956 78343
rect 85956 78321 86008 78343
rect 86008 78321 86010 78343
rect 85954 78309 86010 78321
rect 85954 78287 85956 78309
rect 85956 78287 86008 78309
rect 86008 78287 86010 78309
rect 85954 78257 85956 78263
rect 85956 78257 86008 78263
rect 86008 78257 86010 78263
rect 85954 78245 86010 78257
rect 85954 78207 85956 78245
rect 85956 78207 86008 78245
rect 86008 78207 86010 78245
rect 87042 78705 87044 78743
rect 87044 78705 87096 78743
rect 87096 78705 87098 78743
rect 87042 78693 87098 78705
rect 87042 78687 87044 78693
rect 87044 78687 87096 78693
rect 87096 78687 87098 78693
rect 87042 78641 87044 78663
rect 87044 78641 87096 78663
rect 87096 78641 87098 78663
rect 87042 78629 87098 78641
rect 87042 78607 87044 78629
rect 87044 78607 87096 78629
rect 87096 78607 87098 78629
rect 87042 78577 87044 78583
rect 87044 78577 87096 78583
rect 87096 78577 87098 78583
rect 87042 78565 87098 78577
rect 87042 78527 87044 78565
rect 87044 78527 87096 78565
rect 87096 78527 87098 78565
rect 87042 78501 87098 78503
rect 87042 78449 87044 78501
rect 87044 78449 87096 78501
rect 87096 78449 87098 78501
rect 87042 78447 87098 78449
rect 87042 78385 87044 78423
rect 87044 78385 87096 78423
rect 87096 78385 87098 78423
rect 87042 78373 87098 78385
rect 87042 78367 87044 78373
rect 87044 78367 87096 78373
rect 87096 78367 87098 78373
rect 87042 78321 87044 78343
rect 87044 78321 87096 78343
rect 87096 78321 87098 78343
rect 87042 78309 87098 78321
rect 87042 78287 87044 78309
rect 87044 78287 87096 78309
rect 87096 78287 87098 78309
rect 87042 78257 87044 78263
rect 87044 78257 87096 78263
rect 87096 78257 87098 78263
rect 87042 78245 87098 78257
rect 87042 78207 87044 78245
rect 87044 78207 87096 78245
rect 87096 78207 87098 78245
rect 88130 78705 88132 78743
rect 88132 78705 88184 78743
rect 88184 78705 88186 78743
rect 88130 78693 88186 78705
rect 88130 78687 88132 78693
rect 88132 78687 88184 78693
rect 88184 78687 88186 78693
rect 88130 78641 88132 78663
rect 88132 78641 88184 78663
rect 88184 78641 88186 78663
rect 88130 78629 88186 78641
rect 88130 78607 88132 78629
rect 88132 78607 88184 78629
rect 88184 78607 88186 78629
rect 88130 78577 88132 78583
rect 88132 78577 88184 78583
rect 88184 78577 88186 78583
rect 88130 78565 88186 78577
rect 88130 78527 88132 78565
rect 88132 78527 88184 78565
rect 88184 78527 88186 78565
rect 88130 78501 88186 78503
rect 88130 78449 88132 78501
rect 88132 78449 88184 78501
rect 88184 78449 88186 78501
rect 88130 78447 88186 78449
rect 88130 78385 88132 78423
rect 88132 78385 88184 78423
rect 88184 78385 88186 78423
rect 88130 78373 88186 78385
rect 88130 78367 88132 78373
rect 88132 78367 88184 78373
rect 88184 78367 88186 78373
rect 88130 78321 88132 78343
rect 88132 78321 88184 78343
rect 88184 78321 88186 78343
rect 88130 78309 88186 78321
rect 88130 78287 88132 78309
rect 88132 78287 88184 78309
rect 88184 78287 88186 78309
rect 88130 78257 88132 78263
rect 88132 78257 88184 78263
rect 88184 78257 88186 78263
rect 88130 78245 88186 78257
rect 88130 78207 88132 78245
rect 88132 78207 88184 78245
rect 88184 78207 88186 78245
rect 74529 76708 74531 76746
rect 74531 76708 74583 76746
rect 74583 76708 74585 76746
rect 74529 76696 74585 76708
rect 74529 76690 74531 76696
rect 74531 76690 74583 76696
rect 74583 76690 74585 76696
rect 74529 76644 74531 76666
rect 74531 76644 74583 76666
rect 74583 76644 74585 76666
rect 74529 76632 74585 76644
rect 74529 76610 74531 76632
rect 74531 76610 74583 76632
rect 74583 76610 74585 76632
rect 74529 76580 74531 76586
rect 74531 76580 74583 76586
rect 74583 76580 74585 76586
rect 74529 76568 74585 76580
rect 74529 76530 74531 76568
rect 74531 76530 74583 76568
rect 74583 76530 74585 76568
rect 74529 76504 74585 76506
rect 74529 76452 74531 76504
rect 74531 76452 74583 76504
rect 74583 76452 74585 76504
rect 74529 76450 74585 76452
rect 74529 76388 74531 76426
rect 74531 76388 74583 76426
rect 74583 76388 74585 76426
rect 74529 76376 74585 76388
rect 74529 76370 74531 76376
rect 74531 76370 74583 76376
rect 74583 76370 74585 76376
rect 74529 76324 74531 76346
rect 74531 76324 74583 76346
rect 74583 76324 74585 76346
rect 74529 76312 74585 76324
rect 74529 76290 74531 76312
rect 74531 76290 74583 76312
rect 74583 76290 74585 76312
rect 74529 76260 74531 76266
rect 74531 76260 74583 76266
rect 74583 76260 74585 76266
rect 74529 76248 74585 76260
rect 74529 76210 74531 76248
rect 74531 76210 74583 76248
rect 74583 76210 74585 76248
rect 75617 76708 75619 76746
rect 75619 76708 75671 76746
rect 75671 76708 75673 76746
rect 75617 76696 75673 76708
rect 75617 76690 75619 76696
rect 75619 76690 75671 76696
rect 75671 76690 75673 76696
rect 75617 76644 75619 76666
rect 75619 76644 75671 76666
rect 75671 76644 75673 76666
rect 75617 76632 75673 76644
rect 75617 76610 75619 76632
rect 75619 76610 75671 76632
rect 75671 76610 75673 76632
rect 75617 76580 75619 76586
rect 75619 76580 75671 76586
rect 75671 76580 75673 76586
rect 75617 76568 75673 76580
rect 75617 76530 75619 76568
rect 75619 76530 75671 76568
rect 75671 76530 75673 76568
rect 75617 76504 75673 76506
rect 75617 76452 75619 76504
rect 75619 76452 75671 76504
rect 75671 76452 75673 76504
rect 75617 76450 75673 76452
rect 75617 76388 75619 76426
rect 75619 76388 75671 76426
rect 75671 76388 75673 76426
rect 75617 76376 75673 76388
rect 75617 76370 75619 76376
rect 75619 76370 75671 76376
rect 75671 76370 75673 76376
rect 75617 76324 75619 76346
rect 75619 76324 75671 76346
rect 75671 76324 75673 76346
rect 75617 76312 75673 76324
rect 75617 76290 75619 76312
rect 75619 76290 75671 76312
rect 75671 76290 75673 76312
rect 75617 76260 75619 76266
rect 75619 76260 75671 76266
rect 75671 76260 75673 76266
rect 75617 76248 75673 76260
rect 75617 76210 75619 76248
rect 75619 76210 75671 76248
rect 75671 76210 75673 76248
rect 76705 76708 76707 76746
rect 76707 76708 76759 76746
rect 76759 76708 76761 76746
rect 76705 76696 76761 76708
rect 76705 76690 76707 76696
rect 76707 76690 76759 76696
rect 76759 76690 76761 76696
rect 76705 76644 76707 76666
rect 76707 76644 76759 76666
rect 76759 76644 76761 76666
rect 76705 76632 76761 76644
rect 76705 76610 76707 76632
rect 76707 76610 76759 76632
rect 76759 76610 76761 76632
rect 76705 76580 76707 76586
rect 76707 76580 76759 76586
rect 76759 76580 76761 76586
rect 76705 76568 76761 76580
rect 76705 76530 76707 76568
rect 76707 76530 76759 76568
rect 76759 76530 76761 76568
rect 76705 76504 76761 76506
rect 76705 76452 76707 76504
rect 76707 76452 76759 76504
rect 76759 76452 76761 76504
rect 76705 76450 76761 76452
rect 76705 76388 76707 76426
rect 76707 76388 76759 76426
rect 76759 76388 76761 76426
rect 76705 76376 76761 76388
rect 76705 76370 76707 76376
rect 76707 76370 76759 76376
rect 76759 76370 76761 76376
rect 76705 76324 76707 76346
rect 76707 76324 76759 76346
rect 76759 76324 76761 76346
rect 76705 76312 76761 76324
rect 76705 76290 76707 76312
rect 76707 76290 76759 76312
rect 76759 76290 76761 76312
rect 76705 76260 76707 76266
rect 76707 76260 76759 76266
rect 76759 76260 76761 76266
rect 76705 76248 76761 76260
rect 76705 76210 76707 76248
rect 76707 76210 76759 76248
rect 76759 76210 76761 76248
rect 77793 76708 77795 76746
rect 77795 76708 77847 76746
rect 77847 76708 77849 76746
rect 77793 76696 77849 76708
rect 77793 76690 77795 76696
rect 77795 76690 77847 76696
rect 77847 76690 77849 76696
rect 77793 76644 77795 76666
rect 77795 76644 77847 76666
rect 77847 76644 77849 76666
rect 77793 76632 77849 76644
rect 77793 76610 77795 76632
rect 77795 76610 77847 76632
rect 77847 76610 77849 76632
rect 77793 76580 77795 76586
rect 77795 76580 77847 76586
rect 77847 76580 77849 76586
rect 77793 76568 77849 76580
rect 77793 76530 77795 76568
rect 77795 76530 77847 76568
rect 77847 76530 77849 76568
rect 77793 76504 77849 76506
rect 77793 76452 77795 76504
rect 77795 76452 77847 76504
rect 77847 76452 77849 76504
rect 77793 76450 77849 76452
rect 77793 76388 77795 76426
rect 77795 76388 77847 76426
rect 77847 76388 77849 76426
rect 77793 76376 77849 76388
rect 77793 76370 77795 76376
rect 77795 76370 77847 76376
rect 77847 76370 77849 76376
rect 77793 76324 77795 76346
rect 77795 76324 77847 76346
rect 77847 76324 77849 76346
rect 77793 76312 77849 76324
rect 77793 76290 77795 76312
rect 77795 76290 77847 76312
rect 77847 76290 77849 76312
rect 77793 76260 77795 76266
rect 77795 76260 77847 76266
rect 77847 76260 77849 76266
rect 77793 76248 77849 76260
rect 77793 76210 77795 76248
rect 77795 76210 77847 76248
rect 77847 76210 77849 76248
rect 78881 76708 78883 76746
rect 78883 76708 78935 76746
rect 78935 76708 78937 76746
rect 78881 76696 78937 76708
rect 78881 76690 78883 76696
rect 78883 76690 78935 76696
rect 78935 76690 78937 76696
rect 78881 76644 78883 76666
rect 78883 76644 78935 76666
rect 78935 76644 78937 76666
rect 78881 76632 78937 76644
rect 78881 76610 78883 76632
rect 78883 76610 78935 76632
rect 78935 76610 78937 76632
rect 78881 76580 78883 76586
rect 78883 76580 78935 76586
rect 78935 76580 78937 76586
rect 78881 76568 78937 76580
rect 78881 76530 78883 76568
rect 78883 76530 78935 76568
rect 78935 76530 78937 76568
rect 78881 76504 78937 76506
rect 78881 76452 78883 76504
rect 78883 76452 78935 76504
rect 78935 76452 78937 76504
rect 78881 76450 78937 76452
rect 78881 76388 78883 76426
rect 78883 76388 78935 76426
rect 78935 76388 78937 76426
rect 78881 76376 78937 76388
rect 78881 76370 78883 76376
rect 78883 76370 78935 76376
rect 78935 76370 78937 76376
rect 78881 76324 78883 76346
rect 78883 76324 78935 76346
rect 78935 76324 78937 76346
rect 78881 76312 78937 76324
rect 78881 76290 78883 76312
rect 78883 76290 78935 76312
rect 78935 76290 78937 76312
rect 78881 76260 78883 76266
rect 78883 76260 78935 76266
rect 78935 76260 78937 76266
rect 78881 76248 78937 76260
rect 78881 76210 78883 76248
rect 78883 76210 78935 76248
rect 78935 76210 78937 76248
rect 79969 76708 79971 76746
rect 79971 76708 80023 76746
rect 80023 76708 80025 76746
rect 79969 76696 80025 76708
rect 79969 76690 79971 76696
rect 79971 76690 80023 76696
rect 80023 76690 80025 76696
rect 79969 76644 79971 76666
rect 79971 76644 80023 76666
rect 80023 76644 80025 76666
rect 79969 76632 80025 76644
rect 79969 76610 79971 76632
rect 79971 76610 80023 76632
rect 80023 76610 80025 76632
rect 79969 76580 79971 76586
rect 79971 76580 80023 76586
rect 80023 76580 80025 76586
rect 79969 76568 80025 76580
rect 79969 76530 79971 76568
rect 79971 76530 80023 76568
rect 80023 76530 80025 76568
rect 79969 76504 80025 76506
rect 79969 76452 79971 76504
rect 79971 76452 80023 76504
rect 80023 76452 80025 76504
rect 79969 76450 80025 76452
rect 79969 76388 79971 76426
rect 79971 76388 80023 76426
rect 80023 76388 80025 76426
rect 79969 76376 80025 76388
rect 79969 76370 79971 76376
rect 79971 76370 80023 76376
rect 80023 76370 80025 76376
rect 79969 76324 79971 76346
rect 79971 76324 80023 76346
rect 80023 76324 80025 76346
rect 79969 76312 80025 76324
rect 79969 76290 79971 76312
rect 79971 76290 80023 76312
rect 80023 76290 80025 76312
rect 79969 76260 79971 76266
rect 79971 76260 80023 76266
rect 80023 76260 80025 76266
rect 79969 76248 80025 76260
rect 79969 76210 79971 76248
rect 79971 76210 80023 76248
rect 80023 76210 80025 76248
rect 81057 76708 81059 76746
rect 81059 76708 81111 76746
rect 81111 76708 81113 76746
rect 81057 76696 81113 76708
rect 81057 76690 81059 76696
rect 81059 76690 81111 76696
rect 81111 76690 81113 76696
rect 81057 76644 81059 76666
rect 81059 76644 81111 76666
rect 81111 76644 81113 76666
rect 81057 76632 81113 76644
rect 81057 76610 81059 76632
rect 81059 76610 81111 76632
rect 81111 76610 81113 76632
rect 81057 76580 81059 76586
rect 81059 76580 81111 76586
rect 81111 76580 81113 76586
rect 81057 76568 81113 76580
rect 81057 76530 81059 76568
rect 81059 76530 81111 76568
rect 81111 76530 81113 76568
rect 81057 76504 81113 76506
rect 81057 76452 81059 76504
rect 81059 76452 81111 76504
rect 81111 76452 81113 76504
rect 81057 76450 81113 76452
rect 81057 76388 81059 76426
rect 81059 76388 81111 76426
rect 81111 76388 81113 76426
rect 81057 76376 81113 76388
rect 81057 76370 81059 76376
rect 81059 76370 81111 76376
rect 81111 76370 81113 76376
rect 81057 76324 81059 76346
rect 81059 76324 81111 76346
rect 81111 76324 81113 76346
rect 81057 76312 81113 76324
rect 81057 76290 81059 76312
rect 81059 76290 81111 76312
rect 81111 76290 81113 76312
rect 81057 76260 81059 76266
rect 81059 76260 81111 76266
rect 81111 76260 81113 76266
rect 81057 76248 81113 76260
rect 81057 76210 81059 76248
rect 81059 76210 81111 76248
rect 81111 76210 81113 76248
rect 82145 76708 82147 76746
rect 82147 76708 82199 76746
rect 82199 76708 82201 76746
rect 82145 76696 82201 76708
rect 82145 76690 82147 76696
rect 82147 76690 82199 76696
rect 82199 76690 82201 76696
rect 82145 76644 82147 76666
rect 82147 76644 82199 76666
rect 82199 76644 82201 76666
rect 82145 76632 82201 76644
rect 82145 76610 82147 76632
rect 82147 76610 82199 76632
rect 82199 76610 82201 76632
rect 82145 76580 82147 76586
rect 82147 76580 82199 76586
rect 82199 76580 82201 76586
rect 82145 76568 82201 76580
rect 82145 76530 82147 76568
rect 82147 76530 82199 76568
rect 82199 76530 82201 76568
rect 82145 76504 82201 76506
rect 82145 76452 82147 76504
rect 82147 76452 82199 76504
rect 82199 76452 82201 76504
rect 82145 76450 82201 76452
rect 82145 76388 82147 76426
rect 82147 76388 82199 76426
rect 82199 76388 82201 76426
rect 82145 76376 82201 76388
rect 82145 76370 82147 76376
rect 82147 76370 82199 76376
rect 82199 76370 82201 76376
rect 82145 76324 82147 76346
rect 82147 76324 82199 76346
rect 82199 76324 82201 76346
rect 82145 76312 82201 76324
rect 82145 76290 82147 76312
rect 82147 76290 82199 76312
rect 82199 76290 82201 76312
rect 82145 76260 82147 76266
rect 82147 76260 82199 76266
rect 82199 76260 82201 76266
rect 82145 76248 82201 76260
rect 82145 76210 82147 76248
rect 82147 76210 82199 76248
rect 82199 76210 82201 76248
rect 83233 76708 83235 76746
rect 83235 76708 83287 76746
rect 83287 76708 83289 76746
rect 83233 76696 83289 76708
rect 83233 76690 83235 76696
rect 83235 76690 83287 76696
rect 83287 76690 83289 76696
rect 83233 76644 83235 76666
rect 83235 76644 83287 76666
rect 83287 76644 83289 76666
rect 83233 76632 83289 76644
rect 83233 76610 83235 76632
rect 83235 76610 83287 76632
rect 83287 76610 83289 76632
rect 83233 76580 83235 76586
rect 83235 76580 83287 76586
rect 83287 76580 83289 76586
rect 83233 76568 83289 76580
rect 83233 76530 83235 76568
rect 83235 76530 83287 76568
rect 83287 76530 83289 76568
rect 83233 76504 83289 76506
rect 83233 76452 83235 76504
rect 83235 76452 83287 76504
rect 83287 76452 83289 76504
rect 83233 76450 83289 76452
rect 83233 76388 83235 76426
rect 83235 76388 83287 76426
rect 83287 76388 83289 76426
rect 83233 76376 83289 76388
rect 83233 76370 83235 76376
rect 83235 76370 83287 76376
rect 83287 76370 83289 76376
rect 83233 76324 83235 76346
rect 83235 76324 83287 76346
rect 83287 76324 83289 76346
rect 83233 76312 83289 76324
rect 83233 76290 83235 76312
rect 83235 76290 83287 76312
rect 83287 76290 83289 76312
rect 83233 76260 83235 76266
rect 83235 76260 83287 76266
rect 83287 76260 83289 76266
rect 83233 76248 83289 76260
rect 83233 76210 83235 76248
rect 83235 76210 83287 76248
rect 83287 76210 83289 76248
rect 84321 76708 84323 76746
rect 84323 76708 84375 76746
rect 84375 76708 84377 76746
rect 84321 76696 84377 76708
rect 84321 76690 84323 76696
rect 84323 76690 84375 76696
rect 84375 76690 84377 76696
rect 84321 76644 84323 76666
rect 84323 76644 84375 76666
rect 84375 76644 84377 76666
rect 84321 76632 84377 76644
rect 84321 76610 84323 76632
rect 84323 76610 84375 76632
rect 84375 76610 84377 76632
rect 84321 76580 84323 76586
rect 84323 76580 84375 76586
rect 84375 76580 84377 76586
rect 84321 76568 84377 76580
rect 84321 76530 84323 76568
rect 84323 76530 84375 76568
rect 84375 76530 84377 76568
rect 84321 76504 84377 76506
rect 84321 76452 84323 76504
rect 84323 76452 84375 76504
rect 84375 76452 84377 76504
rect 84321 76450 84377 76452
rect 84321 76388 84323 76426
rect 84323 76388 84375 76426
rect 84375 76388 84377 76426
rect 84321 76376 84377 76388
rect 84321 76370 84323 76376
rect 84323 76370 84375 76376
rect 84375 76370 84377 76376
rect 84321 76324 84323 76346
rect 84323 76324 84375 76346
rect 84375 76324 84377 76346
rect 84321 76312 84377 76324
rect 84321 76290 84323 76312
rect 84323 76290 84375 76312
rect 84375 76290 84377 76312
rect 84321 76260 84323 76266
rect 84323 76260 84375 76266
rect 84375 76260 84377 76266
rect 84321 76248 84377 76260
rect 84321 76210 84323 76248
rect 84323 76210 84375 76248
rect 84375 76210 84377 76248
rect 85409 76708 85411 76746
rect 85411 76708 85463 76746
rect 85463 76708 85465 76746
rect 85409 76696 85465 76708
rect 85409 76690 85411 76696
rect 85411 76690 85463 76696
rect 85463 76690 85465 76696
rect 85409 76644 85411 76666
rect 85411 76644 85463 76666
rect 85463 76644 85465 76666
rect 85409 76632 85465 76644
rect 85409 76610 85411 76632
rect 85411 76610 85463 76632
rect 85463 76610 85465 76632
rect 85409 76580 85411 76586
rect 85411 76580 85463 76586
rect 85463 76580 85465 76586
rect 85409 76568 85465 76580
rect 85409 76530 85411 76568
rect 85411 76530 85463 76568
rect 85463 76530 85465 76568
rect 85409 76504 85465 76506
rect 85409 76452 85411 76504
rect 85411 76452 85463 76504
rect 85463 76452 85465 76504
rect 85409 76450 85465 76452
rect 85409 76388 85411 76426
rect 85411 76388 85463 76426
rect 85463 76388 85465 76426
rect 85409 76376 85465 76388
rect 85409 76370 85411 76376
rect 85411 76370 85463 76376
rect 85463 76370 85465 76376
rect 85409 76324 85411 76346
rect 85411 76324 85463 76346
rect 85463 76324 85465 76346
rect 85409 76312 85465 76324
rect 85409 76290 85411 76312
rect 85411 76290 85463 76312
rect 85463 76290 85465 76312
rect 85409 76260 85411 76266
rect 85411 76260 85463 76266
rect 85463 76260 85465 76266
rect 85409 76248 85465 76260
rect 85409 76210 85411 76248
rect 85411 76210 85463 76248
rect 85463 76210 85465 76248
rect 86497 76708 86499 76746
rect 86499 76708 86551 76746
rect 86551 76708 86553 76746
rect 86497 76696 86553 76708
rect 86497 76690 86499 76696
rect 86499 76690 86551 76696
rect 86551 76690 86553 76696
rect 86497 76644 86499 76666
rect 86499 76644 86551 76666
rect 86551 76644 86553 76666
rect 86497 76632 86553 76644
rect 86497 76610 86499 76632
rect 86499 76610 86551 76632
rect 86551 76610 86553 76632
rect 86497 76580 86499 76586
rect 86499 76580 86551 76586
rect 86551 76580 86553 76586
rect 86497 76568 86553 76580
rect 86497 76530 86499 76568
rect 86499 76530 86551 76568
rect 86551 76530 86553 76568
rect 86497 76504 86553 76506
rect 86497 76452 86499 76504
rect 86499 76452 86551 76504
rect 86551 76452 86553 76504
rect 86497 76450 86553 76452
rect 86497 76388 86499 76426
rect 86499 76388 86551 76426
rect 86551 76388 86553 76426
rect 86497 76376 86553 76388
rect 86497 76370 86499 76376
rect 86499 76370 86551 76376
rect 86551 76370 86553 76376
rect 86497 76324 86499 76346
rect 86499 76324 86551 76346
rect 86551 76324 86553 76346
rect 86497 76312 86553 76324
rect 86497 76290 86499 76312
rect 86499 76290 86551 76312
rect 86551 76290 86553 76312
rect 86497 76260 86499 76266
rect 86499 76260 86551 76266
rect 86551 76260 86553 76266
rect 86497 76248 86553 76260
rect 86497 76210 86499 76248
rect 86499 76210 86551 76248
rect 86551 76210 86553 76248
rect 87585 76708 87587 76746
rect 87587 76708 87639 76746
rect 87639 76708 87641 76746
rect 87585 76696 87641 76708
rect 87585 76690 87587 76696
rect 87587 76690 87639 76696
rect 87639 76690 87641 76696
rect 87585 76644 87587 76666
rect 87587 76644 87639 76666
rect 87639 76644 87641 76666
rect 87585 76632 87641 76644
rect 87585 76610 87587 76632
rect 87587 76610 87639 76632
rect 87639 76610 87641 76632
rect 87585 76580 87587 76586
rect 87587 76580 87639 76586
rect 87639 76580 87641 76586
rect 87585 76568 87641 76580
rect 87585 76530 87587 76568
rect 87587 76530 87639 76568
rect 87639 76530 87641 76568
rect 87585 76504 87641 76506
rect 87585 76452 87587 76504
rect 87587 76452 87639 76504
rect 87639 76452 87641 76504
rect 87585 76450 87641 76452
rect 87585 76388 87587 76426
rect 87587 76388 87639 76426
rect 87639 76388 87641 76426
rect 87585 76376 87641 76388
rect 87585 76370 87587 76376
rect 87587 76370 87639 76376
rect 87639 76370 87641 76376
rect 87585 76324 87587 76346
rect 87587 76324 87639 76346
rect 87639 76324 87641 76346
rect 87585 76312 87641 76324
rect 87585 76290 87587 76312
rect 87587 76290 87639 76312
rect 87639 76290 87641 76312
rect 87585 76260 87587 76266
rect 87587 76260 87639 76266
rect 87639 76260 87641 76266
rect 87585 76248 87641 76260
rect 87585 76210 87587 76248
rect 87587 76210 87639 76248
rect 87639 76210 87641 76248
rect 88673 76708 88675 76746
rect 88675 76708 88727 76746
rect 88727 76708 88729 76746
rect 88673 76696 88729 76708
rect 88673 76690 88675 76696
rect 88675 76690 88727 76696
rect 88727 76690 88729 76696
rect 88673 76644 88675 76666
rect 88675 76644 88727 76666
rect 88727 76644 88729 76666
rect 88673 76632 88729 76644
rect 88673 76610 88675 76632
rect 88675 76610 88727 76632
rect 88727 76610 88729 76632
rect 88673 76580 88675 76586
rect 88675 76580 88727 76586
rect 88727 76580 88729 76586
rect 88673 76568 88729 76580
rect 88673 76530 88675 76568
rect 88675 76530 88727 76568
rect 88727 76530 88729 76568
rect 88673 76504 88729 76506
rect 88673 76452 88675 76504
rect 88675 76452 88727 76504
rect 88727 76452 88729 76504
rect 88673 76450 88729 76452
rect 88673 76388 88675 76426
rect 88675 76388 88727 76426
rect 88727 76388 88729 76426
rect 88673 76376 88729 76388
rect 88673 76370 88675 76376
rect 88675 76370 88727 76376
rect 88727 76370 88729 76376
rect 88673 76324 88675 76346
rect 88675 76324 88727 76346
rect 88727 76324 88729 76346
rect 88673 76312 88729 76324
rect 88673 76290 88675 76312
rect 88675 76290 88727 76312
rect 88727 76290 88729 76312
rect 88673 76260 88675 76266
rect 88675 76260 88727 76266
rect 88727 76260 88729 76266
rect 88673 76248 88729 76260
rect 88673 76210 88675 76248
rect 88675 76210 88727 76248
rect 88727 76210 88729 76248
rect 75074 74705 75076 74743
rect 75076 74705 75128 74743
rect 75128 74705 75130 74743
rect 75074 74693 75130 74705
rect 75074 74687 75076 74693
rect 75076 74687 75128 74693
rect 75128 74687 75130 74693
rect 75074 74641 75076 74663
rect 75076 74641 75128 74663
rect 75128 74641 75130 74663
rect 75074 74629 75130 74641
rect 75074 74607 75076 74629
rect 75076 74607 75128 74629
rect 75128 74607 75130 74629
rect 75074 74577 75076 74583
rect 75076 74577 75128 74583
rect 75128 74577 75130 74583
rect 75074 74565 75130 74577
rect 75074 74527 75076 74565
rect 75076 74527 75128 74565
rect 75128 74527 75130 74565
rect 75074 74501 75130 74503
rect 75074 74449 75076 74501
rect 75076 74449 75128 74501
rect 75128 74449 75130 74501
rect 75074 74447 75130 74449
rect 75074 74385 75076 74423
rect 75076 74385 75128 74423
rect 75128 74385 75130 74423
rect 75074 74373 75130 74385
rect 75074 74367 75076 74373
rect 75076 74367 75128 74373
rect 75128 74367 75130 74373
rect 75074 74321 75076 74343
rect 75076 74321 75128 74343
rect 75128 74321 75130 74343
rect 75074 74309 75130 74321
rect 75074 74287 75076 74309
rect 75076 74287 75128 74309
rect 75128 74287 75130 74309
rect 75074 74257 75076 74263
rect 75076 74257 75128 74263
rect 75128 74257 75130 74263
rect 75074 74245 75130 74257
rect 75074 74207 75076 74245
rect 75076 74207 75128 74245
rect 75128 74207 75130 74245
rect 77250 74705 77252 74743
rect 77252 74705 77304 74743
rect 77304 74705 77306 74743
rect 77250 74693 77306 74705
rect 77250 74687 77252 74693
rect 77252 74687 77304 74693
rect 77304 74687 77306 74693
rect 77250 74641 77252 74663
rect 77252 74641 77304 74663
rect 77304 74641 77306 74663
rect 77250 74629 77306 74641
rect 77250 74607 77252 74629
rect 77252 74607 77304 74629
rect 77304 74607 77306 74629
rect 77250 74577 77252 74583
rect 77252 74577 77304 74583
rect 77304 74577 77306 74583
rect 77250 74565 77306 74577
rect 77250 74527 77252 74565
rect 77252 74527 77304 74565
rect 77304 74527 77306 74565
rect 77250 74501 77306 74503
rect 77250 74449 77252 74501
rect 77252 74449 77304 74501
rect 77304 74449 77306 74501
rect 77250 74447 77306 74449
rect 77250 74385 77252 74423
rect 77252 74385 77304 74423
rect 77304 74385 77306 74423
rect 77250 74373 77306 74385
rect 77250 74367 77252 74373
rect 77252 74367 77304 74373
rect 77304 74367 77306 74373
rect 77250 74321 77252 74343
rect 77252 74321 77304 74343
rect 77304 74321 77306 74343
rect 77250 74309 77306 74321
rect 77250 74287 77252 74309
rect 77252 74287 77304 74309
rect 77304 74287 77306 74309
rect 77250 74257 77252 74263
rect 77252 74257 77304 74263
rect 77304 74257 77306 74263
rect 77250 74245 77306 74257
rect 77250 74207 77252 74245
rect 77252 74207 77304 74245
rect 77304 74207 77306 74245
rect 78338 74705 78340 74743
rect 78340 74705 78392 74743
rect 78392 74705 78394 74743
rect 78338 74693 78394 74705
rect 78338 74687 78340 74693
rect 78340 74687 78392 74693
rect 78392 74687 78394 74693
rect 78338 74641 78340 74663
rect 78340 74641 78392 74663
rect 78392 74641 78394 74663
rect 78338 74629 78394 74641
rect 78338 74607 78340 74629
rect 78340 74607 78392 74629
rect 78392 74607 78394 74629
rect 78338 74577 78340 74583
rect 78340 74577 78392 74583
rect 78392 74577 78394 74583
rect 78338 74565 78394 74577
rect 78338 74527 78340 74565
rect 78340 74527 78392 74565
rect 78392 74527 78394 74565
rect 78338 74501 78394 74503
rect 78338 74449 78340 74501
rect 78340 74449 78392 74501
rect 78392 74449 78394 74501
rect 78338 74447 78394 74449
rect 78338 74385 78340 74423
rect 78340 74385 78392 74423
rect 78392 74385 78394 74423
rect 78338 74373 78394 74385
rect 78338 74367 78340 74373
rect 78340 74367 78392 74373
rect 78392 74367 78394 74373
rect 78338 74321 78340 74343
rect 78340 74321 78392 74343
rect 78392 74321 78394 74343
rect 78338 74309 78394 74321
rect 78338 74287 78340 74309
rect 78340 74287 78392 74309
rect 78392 74287 78394 74309
rect 78338 74257 78340 74263
rect 78340 74257 78392 74263
rect 78392 74257 78394 74263
rect 78338 74245 78394 74257
rect 78338 74207 78340 74245
rect 78340 74207 78392 74245
rect 78392 74207 78394 74245
rect 80514 74705 80516 74743
rect 80516 74705 80568 74743
rect 80568 74705 80570 74743
rect 80514 74693 80570 74705
rect 80514 74687 80516 74693
rect 80516 74687 80568 74693
rect 80568 74687 80570 74693
rect 80514 74641 80516 74663
rect 80516 74641 80568 74663
rect 80568 74641 80570 74663
rect 80514 74629 80570 74641
rect 80514 74607 80516 74629
rect 80516 74607 80568 74629
rect 80568 74607 80570 74629
rect 80514 74577 80516 74583
rect 80516 74577 80568 74583
rect 80568 74577 80570 74583
rect 80514 74565 80570 74577
rect 80514 74527 80516 74565
rect 80516 74527 80568 74565
rect 80568 74527 80570 74565
rect 80514 74501 80570 74503
rect 80514 74449 80516 74501
rect 80516 74449 80568 74501
rect 80568 74449 80570 74501
rect 80514 74447 80570 74449
rect 80514 74385 80516 74423
rect 80516 74385 80568 74423
rect 80568 74385 80570 74423
rect 80514 74373 80570 74385
rect 80514 74367 80516 74373
rect 80516 74367 80568 74373
rect 80568 74367 80570 74373
rect 80514 74321 80516 74343
rect 80516 74321 80568 74343
rect 80568 74321 80570 74343
rect 80514 74309 80570 74321
rect 80514 74287 80516 74309
rect 80516 74287 80568 74309
rect 80568 74287 80570 74309
rect 80514 74257 80516 74263
rect 80516 74257 80568 74263
rect 80568 74257 80570 74263
rect 80514 74245 80570 74257
rect 80514 74207 80516 74245
rect 80516 74207 80568 74245
rect 80568 74207 80570 74245
rect 81602 74705 81604 74743
rect 81604 74705 81656 74743
rect 81656 74705 81658 74743
rect 81602 74693 81658 74705
rect 81602 74687 81604 74693
rect 81604 74687 81656 74693
rect 81656 74687 81658 74693
rect 81602 74641 81604 74663
rect 81604 74641 81656 74663
rect 81656 74641 81658 74663
rect 81602 74629 81658 74641
rect 81602 74607 81604 74629
rect 81604 74607 81656 74629
rect 81656 74607 81658 74629
rect 81602 74577 81604 74583
rect 81604 74577 81656 74583
rect 81656 74577 81658 74583
rect 81602 74565 81658 74577
rect 81602 74527 81604 74565
rect 81604 74527 81656 74565
rect 81656 74527 81658 74565
rect 81602 74501 81658 74503
rect 81602 74449 81604 74501
rect 81604 74449 81656 74501
rect 81656 74449 81658 74501
rect 81602 74447 81658 74449
rect 81602 74385 81604 74423
rect 81604 74385 81656 74423
rect 81656 74385 81658 74423
rect 81602 74373 81658 74385
rect 81602 74367 81604 74373
rect 81604 74367 81656 74373
rect 81656 74367 81658 74373
rect 81602 74321 81604 74343
rect 81604 74321 81656 74343
rect 81656 74321 81658 74343
rect 81602 74309 81658 74321
rect 81602 74287 81604 74309
rect 81604 74287 81656 74309
rect 81656 74287 81658 74309
rect 81602 74257 81604 74263
rect 81604 74257 81656 74263
rect 81656 74257 81658 74263
rect 81602 74245 81658 74257
rect 81602 74207 81604 74245
rect 81604 74207 81656 74245
rect 81656 74207 81658 74245
rect 82690 74705 82692 74743
rect 82692 74705 82744 74743
rect 82744 74705 82746 74743
rect 82690 74693 82746 74705
rect 82690 74687 82692 74693
rect 82692 74687 82744 74693
rect 82744 74687 82746 74693
rect 82690 74641 82692 74663
rect 82692 74641 82744 74663
rect 82744 74641 82746 74663
rect 82690 74629 82746 74641
rect 82690 74607 82692 74629
rect 82692 74607 82744 74629
rect 82744 74607 82746 74629
rect 82690 74577 82692 74583
rect 82692 74577 82744 74583
rect 82744 74577 82746 74583
rect 82690 74565 82746 74577
rect 82690 74527 82692 74565
rect 82692 74527 82744 74565
rect 82744 74527 82746 74565
rect 82690 74501 82746 74503
rect 82690 74449 82692 74501
rect 82692 74449 82744 74501
rect 82744 74449 82746 74501
rect 82690 74447 82746 74449
rect 82690 74385 82692 74423
rect 82692 74385 82744 74423
rect 82744 74385 82746 74423
rect 82690 74373 82746 74385
rect 82690 74367 82692 74373
rect 82692 74367 82744 74373
rect 82744 74367 82746 74373
rect 82690 74321 82692 74343
rect 82692 74321 82744 74343
rect 82744 74321 82746 74343
rect 82690 74309 82746 74321
rect 82690 74287 82692 74309
rect 82692 74287 82744 74309
rect 82744 74287 82746 74309
rect 82690 74257 82692 74263
rect 82692 74257 82744 74263
rect 82744 74257 82746 74263
rect 82690 74245 82746 74257
rect 82690 74207 82692 74245
rect 82692 74207 82744 74245
rect 82744 74207 82746 74245
rect 84866 74705 84868 74743
rect 84868 74705 84920 74743
rect 84920 74705 84922 74743
rect 84866 74693 84922 74705
rect 84866 74687 84868 74693
rect 84868 74687 84920 74693
rect 84920 74687 84922 74693
rect 84866 74641 84868 74663
rect 84868 74641 84920 74663
rect 84920 74641 84922 74663
rect 84866 74629 84922 74641
rect 84866 74607 84868 74629
rect 84868 74607 84920 74629
rect 84920 74607 84922 74629
rect 84866 74577 84868 74583
rect 84868 74577 84920 74583
rect 84920 74577 84922 74583
rect 84866 74565 84922 74577
rect 84866 74527 84868 74565
rect 84868 74527 84920 74565
rect 84920 74527 84922 74565
rect 84866 74501 84922 74503
rect 84866 74449 84868 74501
rect 84868 74449 84920 74501
rect 84920 74449 84922 74501
rect 84866 74447 84922 74449
rect 84866 74385 84868 74423
rect 84868 74385 84920 74423
rect 84920 74385 84922 74423
rect 84866 74373 84922 74385
rect 84866 74367 84868 74373
rect 84868 74367 84920 74373
rect 84920 74367 84922 74373
rect 84866 74321 84868 74343
rect 84868 74321 84920 74343
rect 84920 74321 84922 74343
rect 84866 74309 84922 74321
rect 84866 74287 84868 74309
rect 84868 74287 84920 74309
rect 84920 74287 84922 74309
rect 84866 74257 84868 74263
rect 84868 74257 84920 74263
rect 84920 74257 84922 74263
rect 84866 74245 84922 74257
rect 84866 74207 84868 74245
rect 84868 74207 84920 74245
rect 84920 74207 84922 74245
rect 85954 74705 85956 74743
rect 85956 74705 86008 74743
rect 86008 74705 86010 74743
rect 85954 74693 86010 74705
rect 85954 74687 85956 74693
rect 85956 74687 86008 74693
rect 86008 74687 86010 74693
rect 85954 74641 85956 74663
rect 85956 74641 86008 74663
rect 86008 74641 86010 74663
rect 85954 74629 86010 74641
rect 85954 74607 85956 74629
rect 85956 74607 86008 74629
rect 86008 74607 86010 74629
rect 85954 74577 85956 74583
rect 85956 74577 86008 74583
rect 86008 74577 86010 74583
rect 85954 74565 86010 74577
rect 85954 74527 85956 74565
rect 85956 74527 86008 74565
rect 86008 74527 86010 74565
rect 85954 74501 86010 74503
rect 85954 74449 85956 74501
rect 85956 74449 86008 74501
rect 86008 74449 86010 74501
rect 85954 74447 86010 74449
rect 85954 74385 85956 74423
rect 85956 74385 86008 74423
rect 86008 74385 86010 74423
rect 85954 74373 86010 74385
rect 85954 74367 85956 74373
rect 85956 74367 86008 74373
rect 86008 74367 86010 74373
rect 85954 74321 85956 74343
rect 85956 74321 86008 74343
rect 86008 74321 86010 74343
rect 85954 74309 86010 74321
rect 85954 74287 85956 74309
rect 85956 74287 86008 74309
rect 86008 74287 86010 74309
rect 85954 74257 85956 74263
rect 85956 74257 86008 74263
rect 86008 74257 86010 74263
rect 85954 74245 86010 74257
rect 85954 74207 85956 74245
rect 85956 74207 86008 74245
rect 86008 74207 86010 74245
rect 88130 74705 88132 74743
rect 88132 74705 88184 74743
rect 88184 74705 88186 74743
rect 88130 74693 88186 74705
rect 88130 74687 88132 74693
rect 88132 74687 88184 74693
rect 88184 74687 88186 74693
rect 88130 74641 88132 74663
rect 88132 74641 88184 74663
rect 88184 74641 88186 74663
rect 88130 74629 88186 74641
rect 88130 74607 88132 74629
rect 88132 74607 88184 74629
rect 88184 74607 88186 74629
rect 88130 74577 88132 74583
rect 88132 74577 88184 74583
rect 88184 74577 88186 74583
rect 88130 74565 88186 74577
rect 88130 74527 88132 74565
rect 88132 74527 88184 74565
rect 88184 74527 88186 74565
rect 88130 74501 88186 74503
rect 88130 74449 88132 74501
rect 88132 74449 88184 74501
rect 88184 74449 88186 74501
rect 88130 74447 88186 74449
rect 88130 74385 88132 74423
rect 88132 74385 88184 74423
rect 88184 74385 88186 74423
rect 88130 74373 88186 74385
rect 88130 74367 88132 74373
rect 88132 74367 88184 74373
rect 88184 74367 88186 74373
rect 88130 74321 88132 74343
rect 88132 74321 88184 74343
rect 88184 74321 88186 74343
rect 88130 74309 88186 74321
rect 88130 74287 88132 74309
rect 88132 74287 88184 74309
rect 88184 74287 88186 74309
rect 88130 74257 88132 74263
rect 88132 74257 88184 74263
rect 88184 74257 88186 74263
rect 88130 74245 88186 74257
rect 88130 74207 88132 74245
rect 88132 74207 88184 74245
rect 88184 74207 88186 74245
rect 74529 72708 74531 72746
rect 74531 72708 74583 72746
rect 74583 72708 74585 72746
rect 74529 72696 74585 72708
rect 74529 72690 74531 72696
rect 74531 72690 74583 72696
rect 74583 72690 74585 72696
rect 74529 72644 74531 72666
rect 74531 72644 74583 72666
rect 74583 72644 74585 72666
rect 74529 72632 74585 72644
rect 74529 72610 74531 72632
rect 74531 72610 74583 72632
rect 74583 72610 74585 72632
rect 74529 72580 74531 72586
rect 74531 72580 74583 72586
rect 74583 72580 74585 72586
rect 74529 72568 74585 72580
rect 74529 72530 74531 72568
rect 74531 72530 74583 72568
rect 74583 72530 74585 72568
rect 74529 72504 74585 72506
rect 74529 72452 74531 72504
rect 74531 72452 74583 72504
rect 74583 72452 74585 72504
rect 74529 72450 74585 72452
rect 74529 72388 74531 72426
rect 74531 72388 74583 72426
rect 74583 72388 74585 72426
rect 74529 72376 74585 72388
rect 74529 72370 74531 72376
rect 74531 72370 74583 72376
rect 74583 72370 74585 72376
rect 74529 72324 74531 72346
rect 74531 72324 74583 72346
rect 74583 72324 74585 72346
rect 74529 72312 74585 72324
rect 74529 72290 74531 72312
rect 74531 72290 74583 72312
rect 74583 72290 74585 72312
rect 74529 72260 74531 72266
rect 74531 72260 74583 72266
rect 74583 72260 74585 72266
rect 74529 72248 74585 72260
rect 74529 72210 74531 72248
rect 74531 72210 74583 72248
rect 74583 72210 74585 72248
rect 75617 72708 75619 72746
rect 75619 72708 75671 72746
rect 75671 72708 75673 72746
rect 75617 72696 75673 72708
rect 75617 72690 75619 72696
rect 75619 72690 75671 72696
rect 75671 72690 75673 72696
rect 75617 72644 75619 72666
rect 75619 72644 75671 72666
rect 75671 72644 75673 72666
rect 75617 72632 75673 72644
rect 75617 72610 75619 72632
rect 75619 72610 75671 72632
rect 75671 72610 75673 72632
rect 75617 72580 75619 72586
rect 75619 72580 75671 72586
rect 75671 72580 75673 72586
rect 75617 72568 75673 72580
rect 75617 72530 75619 72568
rect 75619 72530 75671 72568
rect 75671 72530 75673 72568
rect 75617 72504 75673 72506
rect 75617 72452 75619 72504
rect 75619 72452 75671 72504
rect 75671 72452 75673 72504
rect 75617 72450 75673 72452
rect 75617 72388 75619 72426
rect 75619 72388 75671 72426
rect 75671 72388 75673 72426
rect 75617 72376 75673 72388
rect 75617 72370 75619 72376
rect 75619 72370 75671 72376
rect 75671 72370 75673 72376
rect 75617 72324 75619 72346
rect 75619 72324 75671 72346
rect 75671 72324 75673 72346
rect 75617 72312 75673 72324
rect 75617 72290 75619 72312
rect 75619 72290 75671 72312
rect 75671 72290 75673 72312
rect 75617 72260 75619 72266
rect 75619 72260 75671 72266
rect 75671 72260 75673 72266
rect 75617 72248 75673 72260
rect 75617 72210 75619 72248
rect 75619 72210 75671 72248
rect 75671 72210 75673 72248
rect 76705 72708 76707 72746
rect 76707 72708 76759 72746
rect 76759 72708 76761 72746
rect 76705 72696 76761 72708
rect 76705 72690 76707 72696
rect 76707 72690 76759 72696
rect 76759 72690 76761 72696
rect 76705 72644 76707 72666
rect 76707 72644 76759 72666
rect 76759 72644 76761 72666
rect 76705 72632 76761 72644
rect 76705 72610 76707 72632
rect 76707 72610 76759 72632
rect 76759 72610 76761 72632
rect 76705 72580 76707 72586
rect 76707 72580 76759 72586
rect 76759 72580 76761 72586
rect 76705 72568 76761 72580
rect 76705 72530 76707 72568
rect 76707 72530 76759 72568
rect 76759 72530 76761 72568
rect 76705 72504 76761 72506
rect 76705 72452 76707 72504
rect 76707 72452 76759 72504
rect 76759 72452 76761 72504
rect 76705 72450 76761 72452
rect 76705 72388 76707 72426
rect 76707 72388 76759 72426
rect 76759 72388 76761 72426
rect 76705 72376 76761 72388
rect 76705 72370 76707 72376
rect 76707 72370 76759 72376
rect 76759 72370 76761 72376
rect 76705 72324 76707 72346
rect 76707 72324 76759 72346
rect 76759 72324 76761 72346
rect 76705 72312 76761 72324
rect 76705 72290 76707 72312
rect 76707 72290 76759 72312
rect 76759 72290 76761 72312
rect 76705 72260 76707 72266
rect 76707 72260 76759 72266
rect 76759 72260 76761 72266
rect 76705 72248 76761 72260
rect 76705 72210 76707 72248
rect 76707 72210 76759 72248
rect 76759 72210 76761 72248
rect 77793 72708 77795 72746
rect 77795 72708 77847 72746
rect 77847 72708 77849 72746
rect 77793 72696 77849 72708
rect 77793 72690 77795 72696
rect 77795 72690 77847 72696
rect 77847 72690 77849 72696
rect 77793 72644 77795 72666
rect 77795 72644 77847 72666
rect 77847 72644 77849 72666
rect 77793 72632 77849 72644
rect 77793 72610 77795 72632
rect 77795 72610 77847 72632
rect 77847 72610 77849 72632
rect 77793 72580 77795 72586
rect 77795 72580 77847 72586
rect 77847 72580 77849 72586
rect 77793 72568 77849 72580
rect 77793 72530 77795 72568
rect 77795 72530 77847 72568
rect 77847 72530 77849 72568
rect 77793 72504 77849 72506
rect 77793 72452 77795 72504
rect 77795 72452 77847 72504
rect 77847 72452 77849 72504
rect 77793 72450 77849 72452
rect 77793 72388 77795 72426
rect 77795 72388 77847 72426
rect 77847 72388 77849 72426
rect 77793 72376 77849 72388
rect 77793 72370 77795 72376
rect 77795 72370 77847 72376
rect 77847 72370 77849 72376
rect 77793 72324 77795 72346
rect 77795 72324 77847 72346
rect 77847 72324 77849 72346
rect 77793 72312 77849 72324
rect 77793 72290 77795 72312
rect 77795 72290 77847 72312
rect 77847 72290 77849 72312
rect 77793 72260 77795 72266
rect 77795 72260 77847 72266
rect 77847 72260 77849 72266
rect 77793 72248 77849 72260
rect 77793 72210 77795 72248
rect 77795 72210 77847 72248
rect 77847 72210 77849 72248
rect 78881 72708 78883 72746
rect 78883 72708 78935 72746
rect 78935 72708 78937 72746
rect 78881 72696 78937 72708
rect 78881 72690 78883 72696
rect 78883 72690 78935 72696
rect 78935 72690 78937 72696
rect 78881 72644 78883 72666
rect 78883 72644 78935 72666
rect 78935 72644 78937 72666
rect 78881 72632 78937 72644
rect 78881 72610 78883 72632
rect 78883 72610 78935 72632
rect 78935 72610 78937 72632
rect 78881 72580 78883 72586
rect 78883 72580 78935 72586
rect 78935 72580 78937 72586
rect 78881 72568 78937 72580
rect 78881 72530 78883 72568
rect 78883 72530 78935 72568
rect 78935 72530 78937 72568
rect 78881 72504 78937 72506
rect 78881 72452 78883 72504
rect 78883 72452 78935 72504
rect 78935 72452 78937 72504
rect 78881 72450 78937 72452
rect 78881 72388 78883 72426
rect 78883 72388 78935 72426
rect 78935 72388 78937 72426
rect 78881 72376 78937 72388
rect 78881 72370 78883 72376
rect 78883 72370 78935 72376
rect 78935 72370 78937 72376
rect 78881 72324 78883 72346
rect 78883 72324 78935 72346
rect 78935 72324 78937 72346
rect 78881 72312 78937 72324
rect 78881 72290 78883 72312
rect 78883 72290 78935 72312
rect 78935 72290 78937 72312
rect 78881 72260 78883 72266
rect 78883 72260 78935 72266
rect 78935 72260 78937 72266
rect 78881 72248 78937 72260
rect 78881 72210 78883 72248
rect 78883 72210 78935 72248
rect 78935 72210 78937 72248
rect 79969 72708 79971 72746
rect 79971 72708 80023 72746
rect 80023 72708 80025 72746
rect 79969 72696 80025 72708
rect 79969 72690 79971 72696
rect 79971 72690 80023 72696
rect 80023 72690 80025 72696
rect 79969 72644 79971 72666
rect 79971 72644 80023 72666
rect 80023 72644 80025 72666
rect 79969 72632 80025 72644
rect 79969 72610 79971 72632
rect 79971 72610 80023 72632
rect 80023 72610 80025 72632
rect 79969 72580 79971 72586
rect 79971 72580 80023 72586
rect 80023 72580 80025 72586
rect 79969 72568 80025 72580
rect 79969 72530 79971 72568
rect 79971 72530 80023 72568
rect 80023 72530 80025 72568
rect 79969 72504 80025 72506
rect 79969 72452 79971 72504
rect 79971 72452 80023 72504
rect 80023 72452 80025 72504
rect 79969 72450 80025 72452
rect 79969 72388 79971 72426
rect 79971 72388 80023 72426
rect 80023 72388 80025 72426
rect 79969 72376 80025 72388
rect 79969 72370 79971 72376
rect 79971 72370 80023 72376
rect 80023 72370 80025 72376
rect 79969 72324 79971 72346
rect 79971 72324 80023 72346
rect 80023 72324 80025 72346
rect 79969 72312 80025 72324
rect 79969 72290 79971 72312
rect 79971 72290 80023 72312
rect 80023 72290 80025 72312
rect 79969 72260 79971 72266
rect 79971 72260 80023 72266
rect 80023 72260 80025 72266
rect 79969 72248 80025 72260
rect 79969 72210 79971 72248
rect 79971 72210 80023 72248
rect 80023 72210 80025 72248
rect 81057 72708 81059 72746
rect 81059 72708 81111 72746
rect 81111 72708 81113 72746
rect 81057 72696 81113 72708
rect 81057 72690 81059 72696
rect 81059 72690 81111 72696
rect 81111 72690 81113 72696
rect 81057 72644 81059 72666
rect 81059 72644 81111 72666
rect 81111 72644 81113 72666
rect 81057 72632 81113 72644
rect 81057 72610 81059 72632
rect 81059 72610 81111 72632
rect 81111 72610 81113 72632
rect 81057 72580 81059 72586
rect 81059 72580 81111 72586
rect 81111 72580 81113 72586
rect 81057 72568 81113 72580
rect 81057 72530 81059 72568
rect 81059 72530 81111 72568
rect 81111 72530 81113 72568
rect 81057 72504 81113 72506
rect 81057 72452 81059 72504
rect 81059 72452 81111 72504
rect 81111 72452 81113 72504
rect 81057 72450 81113 72452
rect 81057 72388 81059 72426
rect 81059 72388 81111 72426
rect 81111 72388 81113 72426
rect 81057 72376 81113 72388
rect 81057 72370 81059 72376
rect 81059 72370 81111 72376
rect 81111 72370 81113 72376
rect 81057 72324 81059 72346
rect 81059 72324 81111 72346
rect 81111 72324 81113 72346
rect 81057 72312 81113 72324
rect 81057 72290 81059 72312
rect 81059 72290 81111 72312
rect 81111 72290 81113 72312
rect 81057 72260 81059 72266
rect 81059 72260 81111 72266
rect 81111 72260 81113 72266
rect 81057 72248 81113 72260
rect 81057 72210 81059 72248
rect 81059 72210 81111 72248
rect 81111 72210 81113 72248
rect 86497 72708 86499 72746
rect 86499 72708 86551 72746
rect 86551 72708 86553 72746
rect 86497 72696 86553 72708
rect 86497 72690 86499 72696
rect 86499 72690 86551 72696
rect 86551 72690 86553 72696
rect 86497 72644 86499 72666
rect 86499 72644 86551 72666
rect 86551 72644 86553 72666
rect 86497 72632 86553 72644
rect 86497 72610 86499 72632
rect 86499 72610 86551 72632
rect 86551 72610 86553 72632
rect 86497 72580 86499 72586
rect 86499 72580 86551 72586
rect 86551 72580 86553 72586
rect 86497 72568 86553 72580
rect 86497 72530 86499 72568
rect 86499 72530 86551 72568
rect 86551 72530 86553 72568
rect 86497 72504 86553 72506
rect 86497 72452 86499 72504
rect 86499 72452 86551 72504
rect 86551 72452 86553 72504
rect 86497 72450 86553 72452
rect 86497 72388 86499 72426
rect 86499 72388 86551 72426
rect 86551 72388 86553 72426
rect 86497 72376 86553 72388
rect 86497 72370 86499 72376
rect 86499 72370 86551 72376
rect 86551 72370 86553 72376
rect 86497 72324 86499 72346
rect 86499 72324 86551 72346
rect 86551 72324 86553 72346
rect 86497 72312 86553 72324
rect 86497 72290 86499 72312
rect 86499 72290 86551 72312
rect 86551 72290 86553 72312
rect 86497 72260 86499 72266
rect 86499 72260 86551 72266
rect 86551 72260 86553 72266
rect 86497 72248 86553 72260
rect 86497 72210 86499 72248
rect 86499 72210 86551 72248
rect 86551 72210 86553 72248
rect 87585 72708 87587 72746
rect 87587 72708 87639 72746
rect 87639 72708 87641 72746
rect 87585 72696 87641 72708
rect 87585 72690 87587 72696
rect 87587 72690 87639 72696
rect 87639 72690 87641 72696
rect 87585 72644 87587 72666
rect 87587 72644 87639 72666
rect 87639 72644 87641 72666
rect 87585 72632 87641 72644
rect 87585 72610 87587 72632
rect 87587 72610 87639 72632
rect 87639 72610 87641 72632
rect 87585 72580 87587 72586
rect 87587 72580 87639 72586
rect 87639 72580 87641 72586
rect 87585 72568 87641 72580
rect 87585 72530 87587 72568
rect 87587 72530 87639 72568
rect 87639 72530 87641 72568
rect 87585 72504 87641 72506
rect 87585 72452 87587 72504
rect 87587 72452 87639 72504
rect 87639 72452 87641 72504
rect 87585 72450 87641 72452
rect 87585 72388 87587 72426
rect 87587 72388 87639 72426
rect 87639 72388 87641 72426
rect 87585 72376 87641 72388
rect 87585 72370 87587 72376
rect 87587 72370 87639 72376
rect 87639 72370 87641 72376
rect 87585 72324 87587 72346
rect 87587 72324 87639 72346
rect 87639 72324 87641 72346
rect 87585 72312 87641 72324
rect 87585 72290 87587 72312
rect 87587 72290 87639 72312
rect 87639 72290 87641 72312
rect 87585 72260 87587 72266
rect 87587 72260 87639 72266
rect 87639 72260 87641 72266
rect 87585 72248 87641 72260
rect 87585 72210 87587 72248
rect 87587 72210 87639 72248
rect 87639 72210 87641 72248
rect 88673 72708 88675 72746
rect 88675 72708 88727 72746
rect 88727 72708 88729 72746
rect 88673 72696 88729 72708
rect 88673 72690 88675 72696
rect 88675 72690 88727 72696
rect 88727 72690 88729 72696
rect 88673 72644 88675 72666
rect 88675 72644 88727 72666
rect 88727 72644 88729 72666
rect 88673 72632 88729 72644
rect 88673 72610 88675 72632
rect 88675 72610 88727 72632
rect 88727 72610 88729 72632
rect 88673 72580 88675 72586
rect 88675 72580 88727 72586
rect 88727 72580 88729 72586
rect 88673 72568 88729 72580
rect 88673 72530 88675 72568
rect 88675 72530 88727 72568
rect 88727 72530 88729 72568
rect 88673 72504 88729 72506
rect 88673 72452 88675 72504
rect 88675 72452 88727 72504
rect 88727 72452 88729 72504
rect 88673 72450 88729 72452
rect 88673 72388 88675 72426
rect 88675 72388 88727 72426
rect 88727 72388 88729 72426
rect 88673 72376 88729 72388
rect 88673 72370 88675 72376
rect 88675 72370 88727 72376
rect 88727 72370 88729 72376
rect 88673 72324 88675 72346
rect 88675 72324 88727 72346
rect 88727 72324 88729 72346
rect 88673 72312 88729 72324
rect 88673 72290 88675 72312
rect 88675 72290 88727 72312
rect 88727 72290 88729 72312
rect 88673 72260 88675 72266
rect 88675 72260 88727 72266
rect 88727 72260 88729 72266
rect 88673 72248 88729 72260
rect 88673 72210 88675 72248
rect 88675 72210 88727 72248
rect 88727 72210 88729 72248
rect 67310 71660 67606 71662
rect 75074 70705 75076 70743
rect 75076 70705 75128 70743
rect 75128 70705 75130 70743
rect 75074 70693 75130 70705
rect 75074 70687 75076 70693
rect 75076 70687 75128 70693
rect 75128 70687 75130 70693
rect 75074 70641 75076 70663
rect 75076 70641 75128 70663
rect 75128 70641 75130 70663
rect 75074 70629 75130 70641
rect 75074 70607 75076 70629
rect 75076 70607 75128 70629
rect 75128 70607 75130 70629
rect 75074 70577 75076 70583
rect 75076 70577 75128 70583
rect 75128 70577 75130 70583
rect 75074 70565 75130 70577
rect 75074 70527 75076 70565
rect 75076 70527 75128 70565
rect 75128 70527 75130 70565
rect 75074 70501 75130 70503
rect 75074 70449 75076 70501
rect 75076 70449 75128 70501
rect 75128 70449 75130 70501
rect 75074 70447 75130 70449
rect 75074 70385 75076 70423
rect 75076 70385 75128 70423
rect 75128 70385 75130 70423
rect 75074 70373 75130 70385
rect 75074 70367 75076 70373
rect 75076 70367 75128 70373
rect 75128 70367 75130 70373
rect 51203 63880 51339 70256
rect 75074 70321 75076 70343
rect 75076 70321 75128 70343
rect 75128 70321 75130 70343
rect 75074 70309 75130 70321
rect 75074 70287 75076 70309
rect 75076 70287 75128 70309
rect 75128 70287 75130 70309
rect 75074 70257 75076 70263
rect 75076 70257 75128 70263
rect 75128 70257 75130 70263
rect 75074 70245 75130 70257
rect 75074 70207 75076 70245
rect 75076 70207 75128 70245
rect 75128 70207 75130 70245
rect 76162 70705 76164 70743
rect 76164 70705 76216 70743
rect 76216 70705 76218 70743
rect 76162 70693 76218 70705
rect 76162 70687 76164 70693
rect 76164 70687 76216 70693
rect 76216 70687 76218 70693
rect 76162 70641 76164 70663
rect 76164 70641 76216 70663
rect 76216 70641 76218 70663
rect 76162 70629 76218 70641
rect 76162 70607 76164 70629
rect 76164 70607 76216 70629
rect 76216 70607 76218 70629
rect 76162 70577 76164 70583
rect 76164 70577 76216 70583
rect 76216 70577 76218 70583
rect 76162 70565 76218 70577
rect 76162 70527 76164 70565
rect 76164 70527 76216 70565
rect 76216 70527 76218 70565
rect 76162 70501 76218 70503
rect 76162 70449 76164 70501
rect 76164 70449 76216 70501
rect 76216 70449 76218 70501
rect 76162 70447 76218 70449
rect 76162 70385 76164 70423
rect 76164 70385 76216 70423
rect 76216 70385 76218 70423
rect 76162 70373 76218 70385
rect 76162 70367 76164 70373
rect 76164 70367 76216 70373
rect 76216 70367 76218 70373
rect 76162 70321 76164 70343
rect 76164 70321 76216 70343
rect 76216 70321 76218 70343
rect 76162 70309 76218 70321
rect 76162 70287 76164 70309
rect 76164 70287 76216 70309
rect 76216 70287 76218 70309
rect 76162 70257 76164 70263
rect 76164 70257 76216 70263
rect 76216 70257 76218 70263
rect 76162 70245 76218 70257
rect 76162 70207 76164 70245
rect 76164 70207 76216 70245
rect 76216 70207 76218 70245
rect 77250 70705 77252 70743
rect 77252 70705 77304 70743
rect 77304 70705 77306 70743
rect 77250 70693 77306 70705
rect 77250 70687 77252 70693
rect 77252 70687 77304 70693
rect 77304 70687 77306 70693
rect 77250 70641 77252 70663
rect 77252 70641 77304 70663
rect 77304 70641 77306 70663
rect 77250 70629 77306 70641
rect 77250 70607 77252 70629
rect 77252 70607 77304 70629
rect 77304 70607 77306 70629
rect 77250 70577 77252 70583
rect 77252 70577 77304 70583
rect 77304 70577 77306 70583
rect 77250 70565 77306 70577
rect 77250 70527 77252 70565
rect 77252 70527 77304 70565
rect 77304 70527 77306 70565
rect 77250 70501 77306 70503
rect 77250 70449 77252 70501
rect 77252 70449 77304 70501
rect 77304 70449 77306 70501
rect 77250 70447 77306 70449
rect 77250 70385 77252 70423
rect 77252 70385 77304 70423
rect 77304 70385 77306 70423
rect 77250 70373 77306 70385
rect 77250 70367 77252 70373
rect 77252 70367 77304 70373
rect 77304 70367 77306 70373
rect 77250 70321 77252 70343
rect 77252 70321 77304 70343
rect 77304 70321 77306 70343
rect 77250 70309 77306 70321
rect 77250 70287 77252 70309
rect 77252 70287 77304 70309
rect 77304 70287 77306 70309
rect 77250 70257 77252 70263
rect 77252 70257 77304 70263
rect 77304 70257 77306 70263
rect 77250 70245 77306 70257
rect 77250 70207 77252 70245
rect 77252 70207 77304 70245
rect 77304 70207 77306 70245
rect 78338 70705 78340 70743
rect 78340 70705 78392 70743
rect 78392 70705 78394 70743
rect 78338 70693 78394 70705
rect 78338 70687 78340 70693
rect 78340 70687 78392 70693
rect 78392 70687 78394 70693
rect 78338 70641 78340 70663
rect 78340 70641 78392 70663
rect 78392 70641 78394 70663
rect 78338 70629 78394 70641
rect 78338 70607 78340 70629
rect 78340 70607 78392 70629
rect 78392 70607 78394 70629
rect 78338 70577 78340 70583
rect 78340 70577 78392 70583
rect 78392 70577 78394 70583
rect 78338 70565 78394 70577
rect 78338 70527 78340 70565
rect 78340 70527 78392 70565
rect 78392 70527 78394 70565
rect 78338 70501 78394 70503
rect 78338 70449 78340 70501
rect 78340 70449 78392 70501
rect 78392 70449 78394 70501
rect 78338 70447 78394 70449
rect 78338 70385 78340 70423
rect 78340 70385 78392 70423
rect 78392 70385 78394 70423
rect 78338 70373 78394 70385
rect 78338 70367 78340 70373
rect 78340 70367 78392 70373
rect 78392 70367 78394 70373
rect 78338 70321 78340 70343
rect 78340 70321 78392 70343
rect 78392 70321 78394 70343
rect 78338 70309 78394 70321
rect 78338 70287 78340 70309
rect 78340 70287 78392 70309
rect 78392 70287 78394 70309
rect 78338 70257 78340 70263
rect 78340 70257 78392 70263
rect 78392 70257 78394 70263
rect 78338 70245 78394 70257
rect 78338 70207 78340 70245
rect 78340 70207 78392 70245
rect 78392 70207 78394 70245
rect 79426 70705 79428 70743
rect 79428 70705 79480 70743
rect 79480 70705 79482 70743
rect 79426 70693 79482 70705
rect 79426 70687 79428 70693
rect 79428 70687 79480 70693
rect 79480 70687 79482 70693
rect 79426 70641 79428 70663
rect 79428 70641 79480 70663
rect 79480 70641 79482 70663
rect 79426 70629 79482 70641
rect 79426 70607 79428 70629
rect 79428 70607 79480 70629
rect 79480 70607 79482 70629
rect 79426 70577 79428 70583
rect 79428 70577 79480 70583
rect 79480 70577 79482 70583
rect 79426 70565 79482 70577
rect 79426 70527 79428 70565
rect 79428 70527 79480 70565
rect 79480 70527 79482 70565
rect 79426 70501 79482 70503
rect 79426 70449 79428 70501
rect 79428 70449 79480 70501
rect 79480 70449 79482 70501
rect 79426 70447 79482 70449
rect 79426 70385 79428 70423
rect 79428 70385 79480 70423
rect 79480 70385 79482 70423
rect 79426 70373 79482 70385
rect 79426 70367 79428 70373
rect 79428 70367 79480 70373
rect 79480 70367 79482 70373
rect 79426 70321 79428 70343
rect 79428 70321 79480 70343
rect 79480 70321 79482 70343
rect 79426 70309 79482 70321
rect 79426 70287 79428 70309
rect 79428 70287 79480 70309
rect 79480 70287 79482 70309
rect 79426 70257 79428 70263
rect 79428 70257 79480 70263
rect 79480 70257 79482 70263
rect 79426 70245 79482 70257
rect 79426 70207 79428 70245
rect 79428 70207 79480 70245
rect 79480 70207 79482 70245
rect 81602 70705 81604 70743
rect 81604 70705 81656 70743
rect 81656 70705 81658 70743
rect 81602 70693 81658 70705
rect 81602 70687 81604 70693
rect 81604 70687 81656 70693
rect 81656 70687 81658 70693
rect 81602 70641 81604 70663
rect 81604 70641 81656 70663
rect 81656 70641 81658 70663
rect 81602 70629 81658 70641
rect 81602 70607 81604 70629
rect 81604 70607 81656 70629
rect 81656 70607 81658 70629
rect 81602 70577 81604 70583
rect 81604 70577 81656 70583
rect 81656 70577 81658 70583
rect 81602 70565 81658 70577
rect 81602 70527 81604 70565
rect 81604 70527 81656 70565
rect 81656 70527 81658 70565
rect 81602 70501 81658 70503
rect 81602 70449 81604 70501
rect 81604 70449 81656 70501
rect 81656 70449 81658 70501
rect 81602 70447 81658 70449
rect 81602 70385 81604 70423
rect 81604 70385 81656 70423
rect 81656 70385 81658 70423
rect 81602 70373 81658 70385
rect 81602 70367 81604 70373
rect 81604 70367 81656 70373
rect 81656 70367 81658 70373
rect 81602 70321 81604 70343
rect 81604 70321 81656 70343
rect 81656 70321 81658 70343
rect 81602 70309 81658 70321
rect 81602 70287 81604 70309
rect 81604 70287 81656 70309
rect 81656 70287 81658 70309
rect 81602 70257 81604 70263
rect 81604 70257 81656 70263
rect 81656 70257 81658 70263
rect 81602 70245 81658 70257
rect 81602 70207 81604 70245
rect 81604 70207 81656 70245
rect 81656 70207 81658 70245
rect 82690 70705 82692 70743
rect 82692 70705 82744 70743
rect 82744 70705 82746 70743
rect 82690 70693 82746 70705
rect 82690 70687 82692 70693
rect 82692 70687 82744 70693
rect 82744 70687 82746 70693
rect 82690 70641 82692 70663
rect 82692 70641 82744 70663
rect 82744 70641 82746 70663
rect 82690 70629 82746 70641
rect 82690 70607 82692 70629
rect 82692 70607 82744 70629
rect 82744 70607 82746 70629
rect 82690 70577 82692 70583
rect 82692 70577 82744 70583
rect 82744 70577 82746 70583
rect 82690 70565 82746 70577
rect 82690 70527 82692 70565
rect 82692 70527 82744 70565
rect 82744 70527 82746 70565
rect 82690 70501 82746 70503
rect 82690 70449 82692 70501
rect 82692 70449 82744 70501
rect 82744 70449 82746 70501
rect 82690 70447 82746 70449
rect 82690 70385 82692 70423
rect 82692 70385 82744 70423
rect 82744 70385 82746 70423
rect 82690 70373 82746 70385
rect 82690 70367 82692 70373
rect 82692 70367 82744 70373
rect 82744 70367 82746 70373
rect 82690 70321 82692 70343
rect 82692 70321 82744 70343
rect 82744 70321 82746 70343
rect 82690 70309 82746 70321
rect 82690 70287 82692 70309
rect 82692 70287 82744 70309
rect 82744 70287 82746 70309
rect 82690 70257 82692 70263
rect 82692 70257 82744 70263
rect 82744 70257 82746 70263
rect 82690 70245 82746 70257
rect 82690 70207 82692 70245
rect 82692 70207 82744 70245
rect 82744 70207 82746 70245
rect 83778 70705 83780 70743
rect 83780 70705 83832 70743
rect 83832 70705 83834 70743
rect 83778 70693 83834 70705
rect 83778 70687 83780 70693
rect 83780 70687 83832 70693
rect 83832 70687 83834 70693
rect 83778 70641 83780 70663
rect 83780 70641 83832 70663
rect 83832 70641 83834 70663
rect 83778 70629 83834 70641
rect 83778 70607 83780 70629
rect 83780 70607 83832 70629
rect 83832 70607 83834 70629
rect 83778 70577 83780 70583
rect 83780 70577 83832 70583
rect 83832 70577 83834 70583
rect 83778 70565 83834 70577
rect 83778 70527 83780 70565
rect 83780 70527 83832 70565
rect 83832 70527 83834 70565
rect 83778 70501 83834 70503
rect 83778 70449 83780 70501
rect 83780 70449 83832 70501
rect 83832 70449 83834 70501
rect 83778 70447 83834 70449
rect 83778 70385 83780 70423
rect 83780 70385 83832 70423
rect 83832 70385 83834 70423
rect 83778 70373 83834 70385
rect 83778 70367 83780 70373
rect 83780 70367 83832 70373
rect 83832 70367 83834 70373
rect 83778 70321 83780 70343
rect 83780 70321 83832 70343
rect 83832 70321 83834 70343
rect 83778 70309 83834 70321
rect 83778 70287 83780 70309
rect 83780 70287 83832 70309
rect 83832 70287 83834 70309
rect 83778 70257 83780 70263
rect 83780 70257 83832 70263
rect 83832 70257 83834 70263
rect 83778 70245 83834 70257
rect 83778 70207 83780 70245
rect 83780 70207 83832 70245
rect 83832 70207 83834 70245
rect 84866 70705 84868 70743
rect 84868 70705 84920 70743
rect 84920 70705 84922 70743
rect 84866 70693 84922 70705
rect 84866 70687 84868 70693
rect 84868 70687 84920 70693
rect 84920 70687 84922 70693
rect 84866 70641 84868 70663
rect 84868 70641 84920 70663
rect 84920 70641 84922 70663
rect 84866 70629 84922 70641
rect 84866 70607 84868 70629
rect 84868 70607 84920 70629
rect 84920 70607 84922 70629
rect 84866 70577 84868 70583
rect 84868 70577 84920 70583
rect 84920 70577 84922 70583
rect 84866 70565 84922 70577
rect 84866 70527 84868 70565
rect 84868 70527 84920 70565
rect 84920 70527 84922 70565
rect 84866 70501 84922 70503
rect 84866 70449 84868 70501
rect 84868 70449 84920 70501
rect 84920 70449 84922 70501
rect 84866 70447 84922 70449
rect 84866 70385 84868 70423
rect 84868 70385 84920 70423
rect 84920 70385 84922 70423
rect 84866 70373 84922 70385
rect 84866 70367 84868 70373
rect 84868 70367 84920 70373
rect 84920 70367 84922 70373
rect 84866 70321 84868 70343
rect 84868 70321 84920 70343
rect 84920 70321 84922 70343
rect 84866 70309 84922 70321
rect 84866 70287 84868 70309
rect 84868 70287 84920 70309
rect 84920 70287 84922 70309
rect 84866 70257 84868 70263
rect 84868 70257 84920 70263
rect 84920 70257 84922 70263
rect 84866 70245 84922 70257
rect 84866 70207 84868 70245
rect 84868 70207 84920 70245
rect 84920 70207 84922 70245
rect 85954 70705 85956 70743
rect 85956 70705 86008 70743
rect 86008 70705 86010 70743
rect 85954 70693 86010 70705
rect 85954 70687 85956 70693
rect 85956 70687 86008 70693
rect 86008 70687 86010 70693
rect 85954 70641 85956 70663
rect 85956 70641 86008 70663
rect 86008 70641 86010 70663
rect 85954 70629 86010 70641
rect 85954 70607 85956 70629
rect 85956 70607 86008 70629
rect 86008 70607 86010 70629
rect 85954 70577 85956 70583
rect 85956 70577 86008 70583
rect 86008 70577 86010 70583
rect 85954 70565 86010 70577
rect 85954 70527 85956 70565
rect 85956 70527 86008 70565
rect 86008 70527 86010 70565
rect 85954 70501 86010 70503
rect 85954 70449 85956 70501
rect 85956 70449 86008 70501
rect 86008 70449 86010 70501
rect 85954 70447 86010 70449
rect 85954 70385 85956 70423
rect 85956 70385 86008 70423
rect 86008 70385 86010 70423
rect 85954 70373 86010 70385
rect 85954 70367 85956 70373
rect 85956 70367 86008 70373
rect 86008 70367 86010 70373
rect 85954 70321 85956 70343
rect 85956 70321 86008 70343
rect 86008 70321 86010 70343
rect 85954 70309 86010 70321
rect 85954 70287 85956 70309
rect 85956 70287 86008 70309
rect 86008 70287 86010 70309
rect 85954 70257 85956 70263
rect 85956 70257 86008 70263
rect 86008 70257 86010 70263
rect 85954 70245 86010 70257
rect 85954 70207 85956 70245
rect 85956 70207 86008 70245
rect 86008 70207 86010 70245
rect 87042 70705 87044 70743
rect 87044 70705 87096 70743
rect 87096 70705 87098 70743
rect 87042 70693 87098 70705
rect 87042 70687 87044 70693
rect 87044 70687 87096 70693
rect 87096 70687 87098 70693
rect 87042 70641 87044 70663
rect 87044 70641 87096 70663
rect 87096 70641 87098 70663
rect 87042 70629 87098 70641
rect 87042 70607 87044 70629
rect 87044 70607 87096 70629
rect 87096 70607 87098 70629
rect 87042 70577 87044 70583
rect 87044 70577 87096 70583
rect 87096 70577 87098 70583
rect 87042 70565 87098 70577
rect 87042 70527 87044 70565
rect 87044 70527 87096 70565
rect 87096 70527 87098 70565
rect 87042 70501 87098 70503
rect 87042 70449 87044 70501
rect 87044 70449 87096 70501
rect 87096 70449 87098 70501
rect 87042 70447 87098 70449
rect 87042 70385 87044 70423
rect 87044 70385 87096 70423
rect 87096 70385 87098 70423
rect 87042 70373 87098 70385
rect 87042 70367 87044 70373
rect 87044 70367 87096 70373
rect 87096 70367 87098 70373
rect 87042 70321 87044 70343
rect 87044 70321 87096 70343
rect 87096 70321 87098 70343
rect 87042 70309 87098 70321
rect 87042 70287 87044 70309
rect 87044 70287 87096 70309
rect 87096 70287 87098 70309
rect 87042 70257 87044 70263
rect 87044 70257 87096 70263
rect 87096 70257 87098 70263
rect 87042 70245 87098 70257
rect 87042 70207 87044 70245
rect 87044 70207 87096 70245
rect 87096 70207 87098 70245
rect 88130 70705 88132 70743
rect 88132 70705 88184 70743
rect 88184 70705 88186 70743
rect 88130 70693 88186 70705
rect 88130 70687 88132 70693
rect 88132 70687 88184 70693
rect 88184 70687 88186 70693
rect 88130 70641 88132 70663
rect 88132 70641 88184 70663
rect 88184 70641 88186 70663
rect 88130 70629 88186 70641
rect 88130 70607 88132 70629
rect 88132 70607 88184 70629
rect 88184 70607 88186 70629
rect 88130 70577 88132 70583
rect 88132 70577 88184 70583
rect 88184 70577 88186 70583
rect 88130 70565 88186 70577
rect 88130 70527 88132 70565
rect 88132 70527 88184 70565
rect 88184 70527 88186 70565
rect 88130 70501 88186 70503
rect 88130 70449 88132 70501
rect 88132 70449 88184 70501
rect 88184 70449 88186 70501
rect 88130 70447 88186 70449
rect 88130 70385 88132 70423
rect 88132 70385 88184 70423
rect 88184 70385 88186 70423
rect 88130 70373 88186 70385
rect 88130 70367 88132 70373
rect 88132 70367 88184 70373
rect 88184 70367 88186 70373
rect 88130 70321 88132 70343
rect 88132 70321 88184 70343
rect 88184 70321 88186 70343
rect 88130 70309 88186 70321
rect 88130 70287 88132 70309
rect 88132 70287 88184 70309
rect 88184 70287 88186 70309
rect 97687 70337 97743 70393
rect 88130 70257 88132 70263
rect 88132 70257 88184 70263
rect 88184 70257 88186 70263
rect 88130 70245 88186 70257
rect 88130 70207 88132 70245
rect 88132 70207 88184 70245
rect 88184 70207 88186 70245
rect 57477 68355 57613 69851
rect 57458 63893 57468 65389
rect 57468 63893 57584 65389
rect 57584 63893 57594 65389
rect 67311 63911 67607 70127
rect 75343 69764 75399 69766
rect 75343 69712 75345 69764
rect 75345 69712 75397 69764
rect 75397 69712 75399 69764
rect 75343 69710 75399 69712
rect 75889 69764 75945 69766
rect 75889 69712 75891 69764
rect 75891 69712 75943 69764
rect 75943 69712 75945 69764
rect 75889 69710 75945 69712
rect 76435 69755 76491 69757
rect 76435 69703 76437 69755
rect 76437 69703 76489 69755
rect 76489 69703 76491 69755
rect 76435 69701 76491 69703
rect 76980 69754 77036 69756
rect 76980 69702 76982 69754
rect 76982 69702 77034 69754
rect 77034 69702 77036 69754
rect 76980 69700 77036 69702
rect 78611 69742 78667 69744
rect 78611 69690 78613 69742
rect 78613 69690 78665 69742
rect 78665 69690 78667 69742
rect 78611 69688 78667 69690
rect 79154 69739 79210 69741
rect 79154 69687 79156 69739
rect 79156 69687 79208 69739
rect 79208 69687 79210 69739
rect 79154 69685 79210 69687
rect 79696 69738 79752 69740
rect 79696 69686 79698 69738
rect 79698 69686 79750 69738
rect 79750 69686 79752 69738
rect 79696 69684 79752 69686
rect 80243 69743 80299 69745
rect 80243 69691 80245 69743
rect 80245 69691 80297 69743
rect 80297 69691 80299 69743
rect 80243 69689 80299 69691
rect 82961 69754 83017 69756
rect 82961 69702 82963 69754
rect 82963 69702 83015 69754
rect 83015 69702 83017 69754
rect 82961 69700 83017 69702
rect 83504 69758 83560 69760
rect 83504 69706 83506 69758
rect 83506 69706 83558 69758
rect 83558 69706 83560 69758
rect 83504 69704 83560 69706
rect 84046 69752 84102 69754
rect 84046 69700 84048 69752
rect 84048 69700 84100 69752
rect 84100 69700 84102 69752
rect 84046 69698 84102 69700
rect 84603 69743 84659 69745
rect 84603 69691 84605 69743
rect 84605 69691 84657 69743
rect 84657 69691 84659 69743
rect 84603 69689 84659 69691
rect 86227 69754 86283 69756
rect 86227 69702 86229 69754
rect 86229 69702 86281 69754
rect 86281 69702 86283 69754
rect 86227 69700 86283 69702
rect 86771 69747 86827 69749
rect 86771 69695 86773 69747
rect 86773 69695 86825 69747
rect 86825 69695 86827 69747
rect 86771 69693 86827 69695
rect 87321 69751 87377 69753
rect 87321 69699 87323 69751
rect 87323 69699 87375 69751
rect 87375 69699 87377 69751
rect 87321 69697 87377 69699
rect 87854 69751 87910 69753
rect 87854 69699 87856 69751
rect 87856 69699 87908 69751
rect 87908 69699 87910 69751
rect 87854 69697 87910 69699
rect 96655 68907 96711 68909
rect 96655 68855 96657 68907
rect 96657 68855 96709 68907
rect 96709 68855 96711 68907
rect 96655 68853 96711 68855
rect 98244 69781 98300 69837
rect 98086 68953 98142 69009
rect 96655 68717 96711 68719
rect 96655 68665 96657 68717
rect 96657 68665 96709 68717
rect 96709 68665 96711 68717
rect 96655 68663 96711 68665
rect 96655 67757 96711 67759
rect 96655 67705 96657 67757
rect 96657 67705 96709 67757
rect 96709 67705 96711 67757
rect 96655 67703 96711 67705
rect 101856 69088 101912 69090
rect 101936 69088 101992 69090
rect 102016 69088 102072 69090
rect 102096 69088 102152 69090
rect 102176 69088 102232 69090
rect 102256 69088 102312 69090
rect 102336 69088 102392 69090
rect 101856 69036 101874 69088
rect 101874 69036 101912 69088
rect 101936 69036 101938 69088
rect 101938 69036 101990 69088
rect 101990 69036 101992 69088
rect 102016 69036 102054 69088
rect 102054 69036 102066 69088
rect 102066 69036 102072 69088
rect 102096 69036 102118 69088
rect 102118 69036 102130 69088
rect 102130 69036 102152 69088
rect 102176 69036 102182 69088
rect 102182 69036 102194 69088
rect 102194 69036 102232 69088
rect 102256 69036 102258 69088
rect 102258 69036 102310 69088
rect 102310 69036 102312 69088
rect 102336 69036 102374 69088
rect 102374 69036 102392 69088
rect 101856 69034 101912 69036
rect 101936 69034 101992 69036
rect 102016 69034 102072 69036
rect 102096 69034 102152 69036
rect 102176 69034 102232 69036
rect 102256 69034 102312 69036
rect 102336 69034 102392 69036
rect 97986 68569 98042 68625
rect 98086 67803 98142 67859
rect 96655 67567 96711 67569
rect 96655 67515 96657 67567
rect 96657 67515 96709 67567
rect 96709 67515 96711 67567
rect 96655 67513 96711 67515
rect 103398 68933 103614 68951
rect 103398 68753 103416 68933
rect 103416 68753 103596 68933
rect 103596 68753 103614 68933
rect 103398 68735 103614 68753
rect 98641 68542 98697 68544
rect 98721 68542 98777 68544
rect 98801 68542 98857 68544
rect 98881 68542 98937 68544
rect 98641 68490 98687 68542
rect 98687 68490 98697 68542
rect 98721 68490 98751 68542
rect 98751 68490 98763 68542
rect 98763 68490 98777 68542
rect 98801 68490 98815 68542
rect 98815 68490 98827 68542
rect 98827 68490 98857 68542
rect 98881 68490 98891 68542
rect 98891 68490 98937 68542
rect 98641 68488 98697 68490
rect 98721 68488 98777 68490
rect 98801 68488 98857 68490
rect 98881 68488 98937 68490
rect 101895 67937 101951 67939
rect 101975 67937 102031 67939
rect 102055 67937 102111 67939
rect 102135 67937 102191 67939
rect 102215 67937 102271 67939
rect 102295 67937 102351 67939
rect 101895 67885 101925 67937
rect 101925 67885 101937 67937
rect 101937 67885 101951 67937
rect 101975 67885 101989 67937
rect 101989 67885 102001 67937
rect 102001 67885 102031 67937
rect 102055 67885 102065 67937
rect 102065 67885 102111 67937
rect 102135 67885 102181 67937
rect 102181 67885 102191 67937
rect 102215 67885 102245 67937
rect 102245 67885 102257 67937
rect 102257 67885 102271 67937
rect 102295 67885 102309 67937
rect 102309 67885 102321 67937
rect 102321 67885 102351 67937
rect 101895 67883 101951 67885
rect 101975 67883 102031 67885
rect 102055 67883 102111 67885
rect 102135 67883 102191 67885
rect 102215 67883 102271 67885
rect 102295 67883 102351 67885
rect 103386 67782 103602 67800
rect 103386 67602 103404 67782
rect 103404 67602 103584 67782
rect 103584 67602 103602 67782
rect 103386 67584 103602 67602
rect 97986 67419 98042 67475
rect 98639 67392 98695 67394
rect 98719 67392 98775 67394
rect 98799 67392 98855 67394
rect 98879 67392 98935 67394
rect 98639 67340 98685 67392
rect 98685 67340 98695 67392
rect 98719 67340 98749 67392
rect 98749 67340 98761 67392
rect 98761 67340 98775 67392
rect 98799 67340 98813 67392
rect 98813 67340 98825 67392
rect 98825 67340 98855 67392
rect 98879 67340 98889 67392
rect 98889 67340 98935 67392
rect 98639 67338 98695 67340
rect 98719 67338 98775 67340
rect 98799 67338 98855 67340
rect 98879 67338 98935 67340
rect 97687 66647 97743 66703
rect 96655 65217 96711 65219
rect 96655 65165 96657 65217
rect 96657 65165 96709 65217
rect 96709 65165 96711 65217
rect 96655 65163 96711 65165
rect 98244 66091 98300 66147
rect 98086 65263 98142 65319
rect 96655 65027 96711 65029
rect 96655 64975 96657 65027
rect 96657 64975 96709 65027
rect 96709 64975 96711 65027
rect 96655 64973 96711 64975
rect 96655 63947 96711 63949
rect 96655 63895 96657 63947
rect 96657 63895 96709 63947
rect 96709 63895 96711 63947
rect 96655 63893 96711 63895
rect 101885 65395 101941 65397
rect 101965 65395 102021 65397
rect 102045 65395 102101 65397
rect 102125 65395 102181 65397
rect 102205 65395 102261 65397
rect 102285 65395 102341 65397
rect 101885 65343 101915 65395
rect 101915 65343 101927 65395
rect 101927 65343 101941 65395
rect 101965 65343 101979 65395
rect 101979 65343 101991 65395
rect 101991 65343 102021 65395
rect 102045 65343 102055 65395
rect 102055 65343 102101 65395
rect 102125 65343 102171 65395
rect 102171 65343 102181 65395
rect 102205 65343 102235 65395
rect 102235 65343 102247 65395
rect 102247 65343 102261 65395
rect 102285 65343 102299 65395
rect 102299 65343 102311 65395
rect 102311 65343 102341 65395
rect 101885 65341 101941 65343
rect 101965 65341 102021 65343
rect 102045 65341 102101 65343
rect 102125 65341 102181 65343
rect 102205 65341 102261 65343
rect 102285 65341 102341 65343
rect 97986 64879 98042 64935
rect 98086 63993 98142 64049
rect 30032 63703 30034 63749
rect 30034 63703 30086 63749
rect 30086 63703 30088 63749
rect 30032 63693 30088 63703
rect 51430 63710 51432 63846
rect 51432 63710 56924 63846
rect 56924 63710 56926 63846
rect 96655 63757 96711 63759
rect 96655 63705 96657 63757
rect 96657 63705 96709 63757
rect 96709 63705 96711 63757
rect 96655 63703 96711 63705
rect 103244 65250 103460 65268
rect 103244 65070 103262 65250
rect 103262 65070 103442 65250
rect 103442 65070 103460 65250
rect 103244 65052 103460 65070
rect 98557 64851 98613 64853
rect 98637 64851 98693 64853
rect 98717 64851 98773 64853
rect 98797 64851 98853 64853
rect 98557 64799 98603 64851
rect 98603 64799 98613 64851
rect 98637 64799 98667 64851
rect 98667 64799 98679 64851
rect 98679 64799 98693 64851
rect 98717 64799 98731 64851
rect 98731 64799 98743 64851
rect 98743 64799 98773 64851
rect 98797 64799 98807 64851
rect 98807 64799 98853 64851
rect 98557 64797 98613 64799
rect 98637 64797 98693 64799
rect 98717 64797 98773 64799
rect 98797 64797 98853 64799
rect 101885 64125 101941 64127
rect 101965 64125 102021 64127
rect 102045 64125 102101 64127
rect 102125 64125 102181 64127
rect 102205 64125 102261 64127
rect 102285 64125 102341 64127
rect 101885 64073 101915 64125
rect 101915 64073 101927 64125
rect 101927 64073 101941 64125
rect 101965 64073 101979 64125
rect 101979 64073 101991 64125
rect 101991 64073 102021 64125
rect 102045 64073 102055 64125
rect 102055 64073 102101 64125
rect 102125 64073 102171 64125
rect 102171 64073 102181 64125
rect 102205 64073 102235 64125
rect 102235 64073 102247 64125
rect 102247 64073 102261 64125
rect 102285 64073 102299 64125
rect 102299 64073 102311 64125
rect 102311 64073 102341 64125
rect 101885 64071 101941 64073
rect 101965 64071 102021 64073
rect 102045 64071 102101 64073
rect 102125 64071 102181 64073
rect 102205 64071 102261 64073
rect 102285 64071 102341 64073
rect 103215 63960 103431 63978
rect 103215 63780 103233 63960
rect 103233 63780 103413 63960
rect 103413 63780 103431 63960
rect 103215 63762 103431 63780
rect 30032 63639 30034 63669
rect 30034 63639 30086 63669
rect 30086 63639 30088 63669
rect 30032 63627 30088 63639
rect 30032 63613 30034 63627
rect 30034 63613 30086 63627
rect 30086 63613 30088 63627
rect 97986 63609 98042 63665
rect 30032 63575 30034 63589
rect 30034 63575 30086 63589
rect 30086 63575 30088 63589
rect 30032 63563 30088 63575
rect 30032 63533 30034 63563
rect 30034 63533 30086 63563
rect 30086 63533 30088 63563
rect 98555 63582 98611 63584
rect 98635 63582 98691 63584
rect 98715 63582 98771 63584
rect 98795 63582 98851 63584
rect 38221 63490 38223 63520
rect 38223 63490 38275 63520
rect 38275 63490 38277 63520
rect 38221 63478 38277 63490
rect 38221 63464 38223 63478
rect 38223 63464 38275 63478
rect 38275 63464 38277 63478
rect 98555 63530 98601 63582
rect 98601 63530 98611 63582
rect 98635 63530 98665 63582
rect 98665 63530 98677 63582
rect 98677 63530 98691 63582
rect 98715 63530 98729 63582
rect 98729 63530 98741 63582
rect 98741 63530 98771 63582
rect 98795 63530 98805 63582
rect 98805 63530 98851 63582
rect 98555 63528 98611 63530
rect 98635 63528 98691 63530
rect 98715 63528 98771 63530
rect 98795 63528 98851 63530
rect 38221 63426 38223 63440
rect 38223 63426 38275 63440
rect 38275 63426 38277 63440
rect 38221 63414 38277 63426
rect 38221 63384 38223 63414
rect 38223 63384 38275 63414
rect 38275 63384 38277 63414
rect 38221 63350 38277 63360
rect 38221 63304 38223 63350
rect 38223 63304 38275 63350
rect 38275 63304 38277 63350
rect 38221 63234 38223 63280
rect 38223 63234 38275 63280
rect 38275 63234 38277 63280
rect 38221 63224 38277 63234
rect 25286 63120 25288 63166
rect 25288 63120 25340 63166
rect 25340 63120 25342 63166
rect 25286 63110 25342 63120
rect 25286 63056 25288 63086
rect 25288 63056 25340 63086
rect 25340 63056 25342 63086
rect 25286 63044 25342 63056
rect 25286 63030 25288 63044
rect 25288 63030 25340 63044
rect 25340 63030 25342 63044
rect 25286 62992 25288 63006
rect 25288 62992 25340 63006
rect 25340 62992 25342 63006
rect 25286 62980 25342 62992
rect 25286 62950 25288 62980
rect 25288 62950 25340 62980
rect 25340 62950 25342 62980
rect 25286 62916 25342 62926
rect 25286 62870 25288 62916
rect 25288 62870 25340 62916
rect 25340 62870 25342 62916
rect 30026 63088 30028 63126
rect 30028 63088 30080 63126
rect 30080 63088 30082 63126
rect 30026 63076 30082 63088
rect 30026 63070 30028 63076
rect 30028 63070 30080 63076
rect 30080 63070 30082 63076
rect 30026 63024 30028 63046
rect 30028 63024 30080 63046
rect 30080 63024 30082 63046
rect 30026 63012 30082 63024
rect 30026 62990 30028 63012
rect 30028 62990 30080 63012
rect 30080 62990 30082 63012
rect 30026 62960 30028 62966
rect 30028 62960 30080 62966
rect 30080 62960 30082 62966
rect 30026 62948 30082 62960
rect 30026 62910 30028 62948
rect 30028 62910 30080 62948
rect 30080 62910 30082 62948
rect 30026 62884 30082 62886
rect 30026 62832 30028 62884
rect 30028 62832 30080 62884
rect 30080 62832 30082 62884
rect 30026 62830 30082 62832
rect 30026 62768 30028 62806
rect 30028 62768 30080 62806
rect 30080 62768 30082 62806
rect 30026 62756 30082 62768
rect 30026 62750 30028 62756
rect 30028 62750 30080 62756
rect 30080 62750 30082 62756
rect 30026 62704 30028 62726
rect 30028 62704 30080 62726
rect 30080 62704 30082 62726
rect 30026 62692 30082 62704
rect 30026 62670 30028 62692
rect 30028 62670 30080 62692
rect 30080 62670 30082 62692
rect 25287 62617 25343 62627
rect 25287 62571 25289 62617
rect 25289 62571 25341 62617
rect 25341 62571 25343 62617
rect 25287 62501 25289 62547
rect 25289 62501 25341 62547
rect 25341 62501 25343 62547
rect 25287 62491 25343 62501
rect 25287 62437 25289 62467
rect 25289 62437 25341 62467
rect 25341 62437 25343 62467
rect 25287 62425 25343 62437
rect 25287 62411 25289 62425
rect 25289 62411 25341 62425
rect 25341 62411 25343 62425
rect 30026 62640 30028 62646
rect 30028 62640 30080 62646
rect 30080 62640 30082 62646
rect 30026 62628 30082 62640
rect 30026 62590 30028 62628
rect 30028 62590 30080 62628
rect 30080 62590 30082 62628
rect 30026 62564 30082 62566
rect 30026 62512 30028 62564
rect 30028 62512 30080 62564
rect 30080 62512 30082 62564
rect 30026 62510 30082 62512
rect 25287 62373 25289 62387
rect 25289 62373 25341 62387
rect 25341 62373 25343 62387
rect 25287 62361 25343 62373
rect 25287 62331 25289 62361
rect 25289 62331 25341 62361
rect 25341 62331 25343 62361
rect 27484 62429 27540 62431
rect 27564 62429 27620 62431
rect 27644 62429 27700 62431
rect 27724 62429 27780 62431
rect 27804 62429 27860 62431
rect 27884 62429 27940 62431
rect 27484 62377 27494 62429
rect 27494 62377 27540 62429
rect 27564 62377 27610 62429
rect 27610 62377 27620 62429
rect 27644 62377 27674 62429
rect 27674 62377 27686 62429
rect 27686 62377 27700 62429
rect 27724 62377 27738 62429
rect 27738 62377 27750 62429
rect 27750 62377 27780 62429
rect 27804 62377 27814 62429
rect 27814 62377 27860 62429
rect 27884 62377 27930 62429
rect 27930 62377 27940 62429
rect 27484 62375 27540 62377
rect 27564 62375 27620 62377
rect 27644 62375 27700 62377
rect 27724 62375 27780 62377
rect 27804 62375 27860 62377
rect 27884 62375 27940 62377
rect 30026 62448 30028 62486
rect 30028 62448 30080 62486
rect 30080 62448 30082 62486
rect 30026 62436 30082 62448
rect 30026 62430 30028 62436
rect 30028 62430 30080 62436
rect 30080 62430 30082 62436
rect 25287 62297 25343 62307
rect 25287 62251 25289 62297
rect 25289 62251 25341 62297
rect 25341 62251 25343 62297
rect 30026 62384 30028 62406
rect 30028 62384 30080 62406
rect 30080 62384 30082 62406
rect 30026 62372 30082 62384
rect 30026 62350 30028 62372
rect 30028 62350 30080 62372
rect 30080 62350 30082 62372
rect 25287 62181 25289 62227
rect 25289 62181 25341 62227
rect 25341 62181 25343 62227
rect 25287 62171 25343 62181
rect 30026 62320 30028 62326
rect 30028 62320 30080 62326
rect 30080 62320 30082 62326
rect 30026 62308 30082 62320
rect 30026 62270 30028 62308
rect 30028 62270 30080 62308
rect 30080 62270 30082 62308
rect 38221 63170 38223 63200
rect 38223 63170 38275 63200
rect 38275 63170 38277 63200
rect 38221 63158 38277 63170
rect 38221 63144 38223 63158
rect 38223 63144 38275 63158
rect 38275 63144 38277 63158
rect 38221 63106 38223 63120
rect 38223 63106 38275 63120
rect 38275 63106 38277 63120
rect 38221 63094 38277 63106
rect 38221 63064 38223 63094
rect 38223 63064 38275 63094
rect 38275 63064 38277 63094
rect 38221 63030 38277 63040
rect 38221 62984 38223 63030
rect 38223 62984 38275 63030
rect 38275 62984 38277 63030
rect 38221 62914 38223 62960
rect 38223 62914 38275 62960
rect 38275 62914 38277 62960
rect 38221 62904 38277 62914
rect 38221 62850 38223 62880
rect 38223 62850 38275 62880
rect 38275 62850 38277 62880
rect 38221 62838 38277 62850
rect 38221 62824 38223 62838
rect 38223 62824 38275 62838
rect 38275 62824 38277 62838
rect 58571 62840 58627 62896
rect 59620 62873 59676 62891
rect 59620 62835 59622 62873
rect 59622 62835 59674 62873
rect 59674 62835 59676 62873
rect 38221 62786 38223 62800
rect 38223 62786 38275 62800
rect 38275 62786 38277 62800
rect 38221 62774 38277 62786
rect 38221 62744 38223 62774
rect 38223 62744 38275 62774
rect 38275 62744 38277 62774
rect 38221 62710 38277 62720
rect 38221 62664 38223 62710
rect 38223 62664 38275 62710
rect 38275 62664 38277 62710
rect 59620 62809 59676 62811
rect 59620 62757 59622 62809
rect 59622 62757 59674 62809
rect 59674 62757 59676 62809
rect 59620 62755 59676 62757
rect 59620 62693 59622 62731
rect 59622 62693 59674 62731
rect 59674 62693 59676 62731
rect 59620 62675 59676 62693
rect 38221 62594 38223 62640
rect 38223 62594 38275 62640
rect 38275 62594 38277 62640
rect 38221 62584 38277 62594
rect 38221 62530 38223 62560
rect 38223 62530 38275 62560
rect 38275 62530 38277 62560
rect 38221 62518 38277 62530
rect 38221 62504 38223 62518
rect 38223 62504 38275 62518
rect 38275 62504 38277 62518
rect 38221 62466 38223 62480
rect 38223 62466 38275 62480
rect 38275 62466 38277 62480
rect 38221 62454 38277 62466
rect 38221 62424 38223 62454
rect 38223 62424 38275 62454
rect 38275 62424 38277 62454
rect 38221 62390 38277 62400
rect 38221 62344 38223 62390
rect 38223 62344 38275 62390
rect 38275 62344 38277 62390
rect 38221 62274 38223 62320
rect 38223 62274 38275 62320
rect 38275 62274 38277 62320
rect 38221 62264 38277 62274
rect 21586 61562 21802 61580
rect 21586 61382 21604 61562
rect 21604 61382 21784 61562
rect 21784 61382 21802 61562
rect 21586 61364 21802 61382
rect 38221 62210 38223 62240
rect 38223 62210 38275 62240
rect 38275 62210 38277 62240
rect 38221 62198 38277 62210
rect 38221 62184 38223 62198
rect 38223 62184 38275 62198
rect 38275 62184 38277 62198
rect 38221 62146 38223 62160
rect 38223 62146 38275 62160
rect 38275 62146 38277 62160
rect 38221 62134 38277 62146
rect 38221 62104 38223 62134
rect 38223 62104 38275 62134
rect 38275 62104 38277 62134
rect 59630 62416 59686 62418
rect 59630 62364 59632 62416
rect 59632 62364 59684 62416
rect 59684 62364 59686 62416
rect 59630 62362 59686 62364
rect 59630 62300 59632 62338
rect 59632 62300 59684 62338
rect 59684 62300 59686 62338
rect 59630 62288 59686 62300
rect 59630 62282 59632 62288
rect 59632 62282 59684 62288
rect 59684 62282 59686 62288
rect 59630 62236 59632 62258
rect 59632 62236 59684 62258
rect 59684 62236 59686 62258
rect 59630 62224 59686 62236
rect 59630 62202 59632 62224
rect 59632 62202 59684 62224
rect 59684 62202 59686 62224
rect 59630 62172 59632 62178
rect 59632 62172 59684 62178
rect 59684 62172 59686 62178
rect 59630 62160 59686 62172
rect 59630 62122 59632 62160
rect 59632 62122 59684 62160
rect 59684 62122 59686 62160
rect 38221 62070 38277 62080
rect 38221 62024 38223 62070
rect 38223 62024 38275 62070
rect 38275 62024 38277 62070
rect 59094 62031 59150 62087
rect 59630 62096 59686 62098
rect 59630 62044 59632 62096
rect 59632 62044 59684 62096
rect 59684 62044 59686 62096
rect 59630 62042 59686 62044
rect 38221 61954 38223 62000
rect 38223 61954 38275 62000
rect 38275 61954 38277 62000
rect 38221 61944 38277 61954
rect 38221 61890 38223 61920
rect 38223 61890 38275 61920
rect 38275 61890 38277 61920
rect 38221 61878 38277 61890
rect 38221 61864 38223 61878
rect 38223 61864 38275 61878
rect 38275 61864 38277 61878
rect 38221 61826 38223 61840
rect 38223 61826 38275 61840
rect 38275 61826 38277 61840
rect 38221 61814 38277 61826
rect 38221 61784 38223 61814
rect 38223 61784 38275 61814
rect 38275 61784 38277 61814
rect 38221 61750 38277 61760
rect 38221 61704 38223 61750
rect 38223 61704 38275 61750
rect 38275 61704 38277 61750
rect 38221 61634 38223 61680
rect 38223 61634 38275 61680
rect 38275 61634 38277 61680
rect 38221 61624 38277 61634
rect 38221 61570 38223 61600
rect 38223 61570 38275 61600
rect 38275 61570 38277 61600
rect 38221 61558 38277 61570
rect 38221 61544 38223 61558
rect 38223 61544 38275 61558
rect 38275 61544 38277 61558
rect 38221 61506 38223 61520
rect 38223 61506 38275 61520
rect 38275 61506 38277 61520
rect 38221 61494 38277 61506
rect 38221 61464 38223 61494
rect 38223 61464 38275 61494
rect 38275 61464 38277 61494
rect 27468 61339 27524 61341
rect 27548 61339 27604 61341
rect 27628 61339 27684 61341
rect 27708 61339 27764 61341
rect 27788 61339 27844 61341
rect 27868 61339 27924 61341
rect 27468 61287 27498 61339
rect 27498 61287 27510 61339
rect 27510 61287 27524 61339
rect 27548 61287 27562 61339
rect 27562 61287 27574 61339
rect 27574 61287 27604 61339
rect 27628 61287 27638 61339
rect 27638 61287 27684 61339
rect 27708 61287 27754 61339
rect 27754 61287 27764 61339
rect 27788 61287 27818 61339
rect 27818 61287 27830 61339
rect 27830 61287 27844 61339
rect 27868 61287 27882 61339
rect 27882 61287 27894 61339
rect 27894 61287 27924 61339
rect 27468 61285 27524 61287
rect 27548 61285 27604 61287
rect 27628 61285 27684 61287
rect 27708 61285 27764 61287
rect 27788 61285 27844 61287
rect 27868 61285 27924 61287
rect 30029 61321 30031 61359
rect 30031 61321 30083 61359
rect 30083 61321 30085 61359
rect 30029 61309 30085 61321
rect 30029 61303 30031 61309
rect 30031 61303 30083 61309
rect 30083 61303 30085 61309
rect 30029 61257 30031 61279
rect 30031 61257 30083 61279
rect 30083 61257 30085 61279
rect 30029 61245 30085 61257
rect 30029 61223 30031 61245
rect 30031 61223 30083 61245
rect 30083 61223 30085 61245
rect 30029 61193 30031 61199
rect 30031 61193 30083 61199
rect 30083 61193 30085 61199
rect 30029 61181 30085 61193
rect 30029 61143 30031 61181
rect 30031 61143 30083 61181
rect 30083 61143 30085 61181
rect 30029 61117 30085 61119
rect 30029 61065 30031 61117
rect 30031 61065 30083 61117
rect 30083 61065 30085 61117
rect 30029 61063 30085 61065
rect 30029 61001 30031 61039
rect 30031 61001 30083 61039
rect 30083 61001 30085 61039
rect 30029 60989 30085 61001
rect 30029 60983 30031 60989
rect 30031 60983 30083 60989
rect 30083 60983 30085 60989
rect 30029 60937 30031 60959
rect 30031 60937 30083 60959
rect 30083 60937 30085 60959
rect 30029 60925 30085 60937
rect 30029 60903 30031 60925
rect 30031 60903 30083 60925
rect 30083 60903 30085 60925
rect 30029 60873 30031 60879
rect 30031 60873 30083 60879
rect 30083 60873 30085 60879
rect 30029 60861 30085 60873
rect 30029 60823 30031 60861
rect 30031 60823 30083 60861
rect 30083 60823 30085 60861
rect 30029 60797 30085 60799
rect 30029 60745 30031 60797
rect 30031 60745 30083 60797
rect 30083 60745 30085 60797
rect 30029 60743 30085 60745
rect 30029 60681 30031 60719
rect 30031 60681 30083 60719
rect 30083 60681 30085 60719
rect 30029 60669 30085 60681
rect 30029 60663 30031 60669
rect 30031 60663 30083 60669
rect 30083 60663 30085 60669
rect 30029 60617 30031 60639
rect 30031 60617 30083 60639
rect 30083 60617 30085 60639
rect 30029 60605 30085 60617
rect 30029 60583 30031 60605
rect 30031 60583 30083 60605
rect 30083 60583 30085 60605
rect 30029 60553 30031 60559
rect 30031 60553 30083 60559
rect 30083 60553 30085 60559
rect 30029 60541 30085 60553
rect 30029 60503 30031 60541
rect 30031 60503 30083 60541
rect 30083 60503 30085 60541
rect 38221 61430 38277 61440
rect 38221 61384 38223 61430
rect 38223 61384 38275 61430
rect 38275 61384 38277 61430
rect 38221 61314 38223 61360
rect 38223 61314 38275 61360
rect 38275 61314 38277 61360
rect 38221 61304 38277 61314
rect 38221 61250 38223 61280
rect 38223 61250 38275 61280
rect 38275 61250 38277 61280
rect 38221 61238 38277 61250
rect 38221 61224 38223 61238
rect 38223 61224 38275 61238
rect 38275 61224 38277 61238
rect 38221 61186 38223 61200
rect 38223 61186 38275 61200
rect 38275 61186 38277 61200
rect 38221 61174 38277 61186
rect 38221 61144 38223 61174
rect 38223 61144 38275 61174
rect 38275 61144 38277 61174
rect 38221 61110 38277 61120
rect 38221 61064 38223 61110
rect 38223 61064 38275 61110
rect 38275 61064 38277 61110
rect 58571 61091 58627 61147
rect 59266 61115 59268 61153
rect 59268 61115 59320 61153
rect 59320 61115 59322 61153
rect 59266 61103 59322 61115
rect 59266 61097 59268 61103
rect 59268 61097 59320 61103
rect 59320 61097 59322 61103
rect 38221 60994 38223 61040
rect 38223 60994 38275 61040
rect 38275 60994 38277 61040
rect 38221 60984 38277 60994
rect 38221 60930 38223 60960
rect 38223 60930 38275 60960
rect 38275 60930 38277 60960
rect 38221 60918 38277 60930
rect 38221 60904 38223 60918
rect 38223 60904 38275 60918
rect 38275 60904 38277 60918
rect 59266 61051 59268 61073
rect 59268 61051 59320 61073
rect 59320 61051 59322 61073
rect 59266 61039 59322 61051
rect 59266 61017 59268 61039
rect 59268 61017 59320 61039
rect 59320 61017 59322 61039
rect 59266 60987 59268 60993
rect 59268 60987 59320 60993
rect 59320 60987 59322 60993
rect 59266 60975 59322 60987
rect 59266 60937 59268 60975
rect 59268 60937 59320 60975
rect 59320 60937 59322 60975
rect 38221 60866 38223 60880
rect 38223 60866 38275 60880
rect 38275 60866 38277 60880
rect 38221 60854 38277 60866
rect 38221 60824 38223 60854
rect 38223 60824 38275 60854
rect 38275 60824 38277 60854
rect 38221 60790 38277 60800
rect 38221 60744 38223 60790
rect 38223 60744 38275 60790
rect 38275 60744 38277 60790
rect 38221 60674 38223 60720
rect 38223 60674 38275 60720
rect 38275 60674 38277 60720
rect 38221 60664 38277 60674
rect 38221 60610 38223 60640
rect 38223 60610 38275 60640
rect 38275 60610 38277 60640
rect 38221 60598 38277 60610
rect 38221 60584 38223 60598
rect 38223 60584 38275 60598
rect 38275 60584 38277 60598
rect 38221 60546 38223 60560
rect 38223 60546 38275 60560
rect 38275 60546 38277 60560
rect 38221 60534 38277 60546
rect 38221 60504 38223 60534
rect 38223 60504 38275 60534
rect 38275 60504 38277 60534
rect 38221 60470 38277 60480
rect 38221 60424 38223 60470
rect 38223 60424 38275 60470
rect 38275 60424 38277 60470
rect 38221 60354 38223 60400
rect 38223 60354 38275 60400
rect 38275 60354 38277 60400
rect 38221 60344 38277 60354
rect 59267 60667 59323 60669
rect 59267 60615 59269 60667
rect 59269 60615 59321 60667
rect 59321 60615 59323 60667
rect 59267 60613 59323 60615
rect 59267 60551 59269 60589
rect 59269 60551 59321 60589
rect 59321 60551 59323 60589
rect 59267 60539 59323 60551
rect 59267 60533 59269 60539
rect 59269 60533 59321 60539
rect 59321 60533 59323 60539
rect 59267 60487 59269 60509
rect 59269 60487 59321 60509
rect 59321 60487 59323 60509
rect 59267 60475 59323 60487
rect 59267 60453 59269 60475
rect 59269 60453 59321 60475
rect 59321 60453 59323 60475
rect 59267 60423 59269 60429
rect 59269 60423 59321 60429
rect 59321 60423 59323 60429
rect 59267 60411 59323 60423
rect 59267 60373 59269 60411
rect 59269 60373 59321 60411
rect 59321 60373 59323 60411
rect 38221 60290 38223 60320
rect 38223 60290 38275 60320
rect 38275 60290 38277 60320
rect 38221 60278 38277 60290
rect 38221 60264 38223 60278
rect 38223 60264 38275 60278
rect 38275 60264 38277 60278
rect 59094 60281 59150 60337
rect 59267 60347 59323 60349
rect 59267 60295 59269 60347
rect 59269 60295 59321 60347
rect 59321 60295 59323 60347
rect 59267 60293 59323 60295
rect 30029 60112 30031 60142
rect 30031 60112 30083 60142
rect 30083 60112 30085 60142
rect 30029 60100 30085 60112
rect 30029 60086 30031 60100
rect 30031 60086 30083 60100
rect 30083 60086 30085 60100
rect 38221 60226 38223 60240
rect 38223 60226 38275 60240
rect 38275 60226 38277 60240
rect 38221 60214 38277 60226
rect 38221 60184 38223 60214
rect 38223 60184 38275 60214
rect 38275 60184 38277 60214
rect 30029 60048 30031 60062
rect 30031 60048 30083 60062
rect 30083 60048 30085 60062
rect 30029 60036 30085 60048
rect 30029 60006 30031 60036
rect 30031 60006 30083 60036
rect 30083 60006 30085 60036
rect 60046 60107 60102 60109
rect 60126 60107 60182 60109
rect 60206 60107 60262 60109
rect 60286 60107 60342 60109
rect 60366 60107 60422 60109
rect 60046 60055 60048 60107
rect 60048 60055 60100 60107
rect 60100 60055 60102 60107
rect 60126 60055 60164 60107
rect 60164 60055 60176 60107
rect 60176 60055 60182 60107
rect 60206 60055 60228 60107
rect 60228 60055 60240 60107
rect 60240 60055 60262 60107
rect 60286 60055 60292 60107
rect 60292 60055 60304 60107
rect 60304 60055 60342 60107
rect 60366 60055 60368 60107
rect 60368 60055 60420 60107
rect 60420 60055 60422 60107
rect 60046 60053 60102 60055
rect 60126 60053 60182 60055
rect 60206 60053 60262 60055
rect 60286 60053 60342 60055
rect 60366 60053 60422 60055
rect 60682 60110 60738 60112
rect 60762 60110 60818 60112
rect 60842 60110 60898 60112
rect 60682 60058 60700 60110
rect 60700 60058 60738 60110
rect 60762 60058 60764 60110
rect 60764 60058 60816 60110
rect 60816 60058 60818 60110
rect 60842 60058 60880 60110
rect 60880 60058 60898 60110
rect 60682 60056 60738 60058
rect 60762 60056 60818 60058
rect 60842 60056 60898 60058
rect 30029 59972 30085 59982
rect 30029 59926 30031 59972
rect 30031 59926 30083 59972
rect 30083 59926 30085 59972
rect 30029 59856 30031 59902
rect 30031 59856 30083 59902
rect 30083 59856 30085 59902
rect 30029 59846 30085 59856
rect 63443 60559 63499 60615
rect 62149 60109 62205 60111
rect 62229 60109 62285 60111
rect 62309 60109 62365 60111
rect 62389 60109 62445 60111
rect 62149 60057 62175 60109
rect 62175 60057 62205 60109
rect 62229 60057 62239 60109
rect 62239 60057 62285 60109
rect 62309 60057 62355 60109
rect 62355 60057 62365 60109
rect 62389 60057 62419 60109
rect 62419 60057 62445 60109
rect 62149 60055 62205 60057
rect 62229 60055 62285 60057
rect 62309 60055 62365 60057
rect 62389 60055 62445 60057
rect 62673 60110 62729 60112
rect 62753 60110 62809 60112
rect 62833 60110 62889 60112
rect 62673 60058 62691 60110
rect 62691 60058 62729 60110
rect 62753 60058 62755 60110
rect 62755 60058 62807 60110
rect 62807 60058 62809 60110
rect 62833 60058 62871 60110
rect 62871 60058 62889 60110
rect 62673 60056 62729 60058
rect 62753 60056 62809 60058
rect 62833 60056 62889 60058
rect 63443 60215 63499 60271
rect 64032 60102 64088 60104
rect 64112 60102 64168 60104
rect 64192 60102 64248 60104
rect 64032 60050 64050 60102
rect 64050 60050 64088 60102
rect 64112 60050 64114 60102
rect 64114 60050 64166 60102
rect 64166 60050 64168 60102
rect 64192 60050 64230 60102
rect 64230 60050 64248 60102
rect 64032 60048 64088 60050
rect 64112 60048 64168 60050
rect 64192 60048 64248 60050
rect 64478 60109 64534 60111
rect 64558 60109 64614 60111
rect 64638 60109 64694 60111
rect 64718 60109 64774 60111
rect 64478 60057 64504 60109
rect 64504 60057 64534 60109
rect 64558 60057 64568 60109
rect 64568 60057 64614 60109
rect 64638 60057 64684 60109
rect 64684 60057 64694 60109
rect 64718 60057 64748 60109
rect 64748 60057 64774 60109
rect 64478 60055 64534 60057
rect 64558 60055 64614 60057
rect 64638 60055 64694 60057
rect 64718 60055 64774 60057
rect 66040 60108 66096 60110
rect 66120 60108 66176 60110
rect 66200 60108 66256 60110
rect 66280 60108 66336 60110
rect 66360 60108 66416 60110
rect 66040 60056 66042 60108
rect 66042 60056 66094 60108
rect 66094 60056 66096 60108
rect 66120 60056 66158 60108
rect 66158 60056 66170 60108
rect 66170 60056 66176 60108
rect 66200 60056 66222 60108
rect 66222 60056 66234 60108
rect 66234 60056 66256 60108
rect 66280 60056 66286 60108
rect 66286 60056 66298 60108
rect 66298 60056 66336 60108
rect 66360 60056 66362 60108
rect 66362 60056 66414 60108
rect 66414 60056 66416 60108
rect 66040 60054 66096 60056
rect 66120 60054 66176 60056
rect 66200 60054 66256 60056
rect 66280 60054 66336 60056
rect 66360 60054 66416 60056
rect 66674 60105 66730 60107
rect 66754 60105 66810 60107
rect 66834 60105 66890 60107
rect 66674 60053 66692 60105
rect 66692 60053 66730 60105
rect 66754 60053 66756 60105
rect 66756 60053 66808 60105
rect 66808 60053 66810 60105
rect 66834 60053 66872 60105
rect 66872 60053 66890 60105
rect 66674 60051 66730 60053
rect 66754 60051 66810 60053
rect 66834 60051 66890 60053
rect 30029 59792 30031 59822
rect 30031 59792 30083 59822
rect 30083 59792 30085 59822
rect 30029 59780 30085 59792
rect 30029 59766 30031 59780
rect 30031 59766 30083 59780
rect 30083 59766 30085 59780
rect 30029 59728 30031 59742
rect 30031 59728 30083 59742
rect 30083 59728 30085 59742
rect 30029 59716 30085 59728
rect 30029 59686 30031 59716
rect 30031 59686 30083 59716
rect 30083 59686 30085 59716
rect 30029 59652 30085 59662
rect 30029 59606 30031 59652
rect 30031 59606 30083 59652
rect 30083 59606 30085 59652
rect 30029 59536 30031 59582
rect 30031 59536 30083 59582
rect 30083 59536 30085 59582
rect 30029 59526 30085 59536
rect 30029 59472 30031 59502
rect 30031 59472 30083 59502
rect 30083 59472 30085 59502
rect 30029 59460 30085 59472
rect 30029 59446 30031 59460
rect 30031 59446 30083 59460
rect 30083 59446 30085 59460
rect 30029 59408 30031 59422
rect 30031 59408 30083 59422
rect 30083 59408 30085 59422
rect 30029 59396 30085 59408
rect 30029 59366 30031 59396
rect 30031 59366 30083 59396
rect 30083 59366 30085 59396
rect 30029 59332 30085 59342
rect 30029 59286 30031 59332
rect 30031 59286 30083 59332
rect 30083 59286 30085 59332
rect 30029 59216 30031 59262
rect 30031 59216 30083 59262
rect 30083 59216 30085 59262
rect 30029 59206 30085 59216
rect 30029 59152 30031 59182
rect 30031 59152 30083 59182
rect 30083 59152 30085 59182
rect 30029 59140 30085 59152
rect 30029 59126 30031 59140
rect 30031 59126 30083 59140
rect 30083 59126 30085 59140
rect 30029 59088 30031 59102
rect 30031 59088 30083 59102
rect 30083 59088 30085 59102
rect 30029 59076 30085 59088
rect 30029 59046 30031 59076
rect 30031 59046 30083 59076
rect 30083 59046 30085 59076
rect 30026 58686 30082 58704
rect 30026 58648 30028 58686
rect 30028 58648 30080 58686
rect 30080 58648 30082 58686
rect 47729 58692 47785 58694
rect 47729 58640 47731 58692
rect 47731 58640 47783 58692
rect 47783 58640 47785 58692
rect 47729 58638 47785 58640
rect 30026 58622 30082 58624
rect 30026 58570 30028 58622
rect 30028 58570 30080 58622
rect 30080 58570 30082 58622
rect 30026 58568 30082 58570
rect 30026 58506 30028 58544
rect 30028 58506 30080 58544
rect 30080 58506 30082 58544
rect 30026 58494 30082 58506
rect 30026 58488 30028 58494
rect 30028 58488 30080 58494
rect 30080 58488 30082 58494
rect 30026 58442 30028 58464
rect 30028 58442 30080 58464
rect 30080 58442 30082 58464
rect 30026 58430 30082 58442
rect 30026 58408 30028 58430
rect 30028 58408 30080 58430
rect 30080 58408 30082 58430
rect 30026 58378 30028 58384
rect 30028 58378 30080 58384
rect 30080 58378 30082 58384
rect 30026 58366 30082 58378
rect 30026 58328 30028 58366
rect 30028 58328 30080 58366
rect 30080 58328 30082 58366
rect 30026 58302 30082 58304
rect 30026 58250 30028 58302
rect 30028 58250 30080 58302
rect 30080 58250 30082 58302
rect 30026 58248 30082 58250
rect 30026 58186 30028 58224
rect 30028 58186 30080 58224
rect 30080 58186 30082 58224
rect 30026 58174 30082 58186
rect 30026 58168 30028 58174
rect 30028 58168 30080 58174
rect 30080 58168 30082 58174
rect 63030 58157 63086 58213
rect 30026 58122 30028 58144
rect 30028 58122 30080 58144
rect 30080 58122 30082 58144
rect 30026 58110 30082 58122
rect 30026 58088 30028 58110
rect 30028 58088 30080 58110
rect 30080 58088 30082 58110
rect 30026 58058 30028 58064
rect 30028 58058 30080 58064
rect 30080 58058 30082 58064
rect 30026 58046 30082 58058
rect 30026 58008 30028 58046
rect 30028 58008 30080 58046
rect 30080 58008 30082 58046
rect 30026 57982 30082 57984
rect 30026 57930 30028 57982
rect 30028 57930 30080 57982
rect 30080 57930 30082 57982
rect 30026 57928 30082 57930
rect 30026 57866 30028 57904
rect 30028 57866 30080 57904
rect 30080 57866 30082 57904
rect 30026 57854 30082 57866
rect 30026 57848 30028 57854
rect 30028 57848 30080 57854
rect 30080 57848 30082 57854
rect 30026 57802 30028 57824
rect 30028 57802 30080 57824
rect 30080 57802 30082 57824
rect 30026 57790 30082 57802
rect 30026 57768 30028 57790
rect 30028 57768 30080 57790
rect 30080 57768 30082 57790
rect 63836 57812 63892 57868
rect 30026 57738 30028 57744
rect 30028 57738 30080 57744
rect 30080 57738 30082 57744
rect 30026 57726 30082 57738
rect 30026 57688 30028 57726
rect 30028 57688 30080 57726
rect 30080 57688 30082 57726
rect 30026 57662 30082 57664
rect 30026 57610 30028 57662
rect 30028 57610 30080 57662
rect 30080 57610 30082 57662
rect 30026 57608 30082 57610
rect 30026 57546 30028 57584
rect 30028 57546 30080 57584
rect 30080 57546 30082 57584
rect 30026 57528 30082 57546
rect 35580 57513 35636 57569
rect 50150 57195 50206 57197
rect 50150 57143 50152 57195
rect 50152 57143 50204 57195
rect 50204 57143 50206 57195
rect 50150 57141 50206 57143
rect 30021 56852 30023 56882
rect 30023 56852 30075 56882
rect 30075 56852 30077 56882
rect 30021 56840 30077 56852
rect 30021 56826 30023 56840
rect 30023 56826 30075 56840
rect 30075 56826 30077 56840
rect 30021 56788 30023 56802
rect 30023 56788 30075 56802
rect 30075 56788 30077 56802
rect 30021 56776 30077 56788
rect 30021 56746 30023 56776
rect 30023 56746 30075 56776
rect 30075 56746 30077 56776
rect 30021 56712 30077 56722
rect 30021 56666 30023 56712
rect 30023 56666 30075 56712
rect 30075 56666 30077 56712
rect 30021 56596 30023 56642
rect 30023 56596 30075 56642
rect 30075 56596 30077 56642
rect 30021 56586 30077 56596
rect 30021 56532 30023 56562
rect 30023 56532 30075 56562
rect 30075 56532 30077 56562
rect 30021 56520 30077 56532
rect 30021 56506 30023 56520
rect 30023 56506 30075 56520
rect 30075 56506 30077 56520
rect 30021 56468 30023 56482
rect 30023 56468 30075 56482
rect 30075 56468 30077 56482
rect 30021 56456 30077 56468
rect 30021 56426 30023 56456
rect 30023 56426 30075 56456
rect 30075 56426 30077 56456
rect 62415 56307 62471 56363
rect 64462 56314 64518 56370
rect 65063 55773 65119 55829
rect 61452 54448 61508 54450
rect 61452 54396 61454 54448
rect 61454 54396 61506 54448
rect 61506 54396 61508 54448
rect 61452 54394 61508 54396
rect 65426 54453 65482 54455
rect 65426 54401 65428 54453
rect 65428 54401 65480 54453
rect 65480 54401 65482 54453
rect 65426 54399 65482 54401
rect 60424 54267 60480 54323
rect 44405 53768 44461 53770
rect 44405 53716 44407 53768
rect 44407 53716 44459 53768
rect 44459 53716 44461 53768
rect 44405 53714 44461 53716
rect 59011 53714 59067 53770
rect 73819 53714 73875 53770
rect 43629 53345 43685 53347
rect 43629 53293 43631 53345
rect 43631 53293 43683 53345
rect 43683 53293 43685 53345
rect 43629 53291 43685 53293
rect 59011 53291 59067 53347
rect 74510 53291 74566 53347
rect 18943 50610 18999 50612
rect 19023 50610 19079 50612
rect 19103 50610 19159 50612
rect 19183 50610 19239 50612
rect 19263 50610 19319 50612
rect 19343 50610 19399 50612
rect 19423 50610 19479 50612
rect 19503 50610 19559 50612
rect 19583 50610 19639 50612
rect 19663 50610 19719 50612
rect 19743 50610 19799 50612
rect 19823 50610 19879 50612
rect 19903 50610 19959 50612
rect 19983 50610 20039 50612
rect 20063 50610 20119 50612
rect 20143 50610 20199 50612
rect 20223 50610 20279 50612
rect 20303 50610 20359 50612
rect 20383 50610 20439 50612
rect 20463 50610 20519 50612
rect 20543 50610 20599 50612
rect 20623 50610 20679 50612
rect 20703 50610 20759 50612
rect 20783 50610 20839 50612
rect 20863 50610 20919 50612
rect 20943 50610 20999 50612
rect 21023 50610 21079 50612
rect 21103 50610 21159 50612
rect 21183 50610 21239 50612
rect 21263 50610 21319 50612
rect 21343 50610 21399 50612
rect 21423 50610 21479 50612
rect 21503 50610 21559 50612
rect 21583 50610 21639 50612
rect 21663 50610 21719 50612
rect 21743 50610 21799 50612
rect 21823 50610 21879 50612
rect 21903 50610 21959 50612
rect 21983 50610 22039 50612
rect 22063 50610 22119 50612
rect 22143 50610 22199 50612
rect 18943 50558 18965 50610
rect 18965 50558 18977 50610
rect 18977 50558 18999 50610
rect 19023 50558 19029 50610
rect 19029 50558 19041 50610
rect 19041 50558 19079 50610
rect 19103 50558 19105 50610
rect 19105 50558 19157 50610
rect 19157 50558 19159 50610
rect 19183 50558 19221 50610
rect 19221 50558 19233 50610
rect 19233 50558 19239 50610
rect 19263 50558 19285 50610
rect 19285 50558 19297 50610
rect 19297 50558 19319 50610
rect 19343 50558 19349 50610
rect 19349 50558 19361 50610
rect 19361 50558 19399 50610
rect 19423 50558 19425 50610
rect 19425 50558 19477 50610
rect 19477 50558 19479 50610
rect 19503 50558 19541 50610
rect 19541 50558 19553 50610
rect 19553 50558 19559 50610
rect 19583 50558 19605 50610
rect 19605 50558 19617 50610
rect 19617 50558 19639 50610
rect 19663 50558 19669 50610
rect 19669 50558 19681 50610
rect 19681 50558 19719 50610
rect 19743 50558 19745 50610
rect 19745 50558 19797 50610
rect 19797 50558 19799 50610
rect 19823 50558 19861 50610
rect 19861 50558 19873 50610
rect 19873 50558 19879 50610
rect 19903 50558 19925 50610
rect 19925 50558 19937 50610
rect 19937 50558 19959 50610
rect 19983 50558 19989 50610
rect 19989 50558 20001 50610
rect 20001 50558 20039 50610
rect 20063 50558 20065 50610
rect 20065 50558 20117 50610
rect 20117 50558 20119 50610
rect 20143 50558 20181 50610
rect 20181 50558 20193 50610
rect 20193 50558 20199 50610
rect 20223 50558 20245 50610
rect 20245 50558 20257 50610
rect 20257 50558 20279 50610
rect 20303 50558 20309 50610
rect 20309 50558 20321 50610
rect 20321 50558 20359 50610
rect 20383 50558 20385 50610
rect 20385 50558 20437 50610
rect 20437 50558 20439 50610
rect 20463 50558 20501 50610
rect 20501 50558 20513 50610
rect 20513 50558 20519 50610
rect 20543 50558 20565 50610
rect 20565 50558 20577 50610
rect 20577 50558 20599 50610
rect 20623 50558 20629 50610
rect 20629 50558 20641 50610
rect 20641 50558 20679 50610
rect 20703 50558 20705 50610
rect 20705 50558 20757 50610
rect 20757 50558 20759 50610
rect 20783 50558 20821 50610
rect 20821 50558 20833 50610
rect 20833 50558 20839 50610
rect 20863 50558 20885 50610
rect 20885 50558 20897 50610
rect 20897 50558 20919 50610
rect 20943 50558 20949 50610
rect 20949 50558 20961 50610
rect 20961 50558 20999 50610
rect 21023 50558 21025 50610
rect 21025 50558 21077 50610
rect 21077 50558 21079 50610
rect 21103 50558 21141 50610
rect 21141 50558 21153 50610
rect 21153 50558 21159 50610
rect 21183 50558 21205 50610
rect 21205 50558 21217 50610
rect 21217 50558 21239 50610
rect 21263 50558 21269 50610
rect 21269 50558 21281 50610
rect 21281 50558 21319 50610
rect 21343 50558 21345 50610
rect 21345 50558 21397 50610
rect 21397 50558 21399 50610
rect 21423 50558 21461 50610
rect 21461 50558 21473 50610
rect 21473 50558 21479 50610
rect 21503 50558 21525 50610
rect 21525 50558 21537 50610
rect 21537 50558 21559 50610
rect 21583 50558 21589 50610
rect 21589 50558 21601 50610
rect 21601 50558 21639 50610
rect 21663 50558 21665 50610
rect 21665 50558 21717 50610
rect 21717 50558 21719 50610
rect 21743 50558 21781 50610
rect 21781 50558 21793 50610
rect 21793 50558 21799 50610
rect 21823 50558 21845 50610
rect 21845 50558 21857 50610
rect 21857 50558 21879 50610
rect 21903 50558 21909 50610
rect 21909 50558 21921 50610
rect 21921 50558 21959 50610
rect 21983 50558 21985 50610
rect 21985 50558 22037 50610
rect 22037 50558 22039 50610
rect 22063 50558 22101 50610
rect 22101 50558 22113 50610
rect 22113 50558 22119 50610
rect 22143 50558 22165 50610
rect 22165 50558 22177 50610
rect 22177 50558 22199 50610
rect 18943 50556 18999 50558
rect 19023 50556 19079 50558
rect 19103 50556 19159 50558
rect 19183 50556 19239 50558
rect 19263 50556 19319 50558
rect 19343 50556 19399 50558
rect 19423 50556 19479 50558
rect 19503 50556 19559 50558
rect 19583 50556 19639 50558
rect 19663 50556 19719 50558
rect 19743 50556 19799 50558
rect 19823 50556 19879 50558
rect 19903 50556 19959 50558
rect 19983 50556 20039 50558
rect 20063 50556 20119 50558
rect 20143 50556 20199 50558
rect 20223 50556 20279 50558
rect 20303 50556 20359 50558
rect 20383 50556 20439 50558
rect 20463 50556 20519 50558
rect 20543 50556 20599 50558
rect 20623 50556 20679 50558
rect 20703 50556 20759 50558
rect 20783 50556 20839 50558
rect 20863 50556 20919 50558
rect 20943 50556 20999 50558
rect 21023 50556 21079 50558
rect 21103 50556 21159 50558
rect 21183 50556 21239 50558
rect 21263 50556 21319 50558
rect 21343 50556 21399 50558
rect 21423 50556 21479 50558
rect 21503 50556 21559 50558
rect 21583 50556 21639 50558
rect 21663 50556 21719 50558
rect 21743 50556 21799 50558
rect 21823 50556 21879 50558
rect 21903 50556 21959 50558
rect 21983 50556 22039 50558
rect 22063 50556 22119 50558
rect 22143 50556 22199 50558
rect 61799 52770 61855 52826
rect 65058 52862 65114 52864
rect 65058 52810 65060 52862
rect 65060 52810 65112 52862
rect 65112 52810 65114 52862
rect 65058 52808 65114 52810
rect 41403 52059 41405 52081
rect 41405 52059 41457 52081
rect 41457 52059 41459 52081
rect 41403 52047 41459 52059
rect 41403 52025 41405 52047
rect 41405 52025 41457 52047
rect 41457 52025 41459 52047
rect 41403 51995 41405 52001
rect 41405 51995 41457 52001
rect 41457 51995 41459 52001
rect 41403 51983 41459 51995
rect 41403 51945 41405 51983
rect 41405 51945 41457 51983
rect 41457 51945 41459 51983
rect 41403 51919 41459 51921
rect 41403 51867 41405 51919
rect 41405 51867 41457 51919
rect 41457 51867 41459 51919
rect 41403 51865 41459 51867
rect 41403 51803 41405 51841
rect 41405 51803 41457 51841
rect 41457 51803 41459 51841
rect 41403 51791 41459 51803
rect 41403 51785 41405 51791
rect 41405 51785 41457 51791
rect 41457 51785 41459 51791
rect 41403 51739 41405 51761
rect 41405 51739 41457 51761
rect 41457 51739 41459 51761
rect 41403 51727 41459 51739
rect 41403 51705 41405 51727
rect 41405 51705 41457 51727
rect 41457 51705 41459 51727
rect 39495 51574 39551 51630
rect 39495 50345 39551 50401
rect 41385 50274 41441 50292
rect 41385 50236 41387 50274
rect 41387 50236 41439 50274
rect 41439 50236 41441 50274
rect 41385 50210 41441 50212
rect 41385 50158 41387 50210
rect 41387 50158 41439 50210
rect 41439 50158 41441 50210
rect 41385 50156 41441 50158
rect 41385 50094 41387 50132
rect 41387 50094 41439 50132
rect 41439 50094 41441 50132
rect 41385 50076 41441 50094
rect 44713 52081 44769 52083
rect 44713 52029 44715 52081
rect 44715 52029 44767 52081
rect 44767 52029 44769 52081
rect 44713 52027 44769 52029
rect 44713 51965 44715 52003
rect 44715 51965 44767 52003
rect 44767 51965 44769 52003
rect 44713 51953 44769 51965
rect 44713 51947 44715 51953
rect 44715 51947 44767 51953
rect 44767 51947 44769 51953
rect 44713 51901 44715 51923
rect 44715 51901 44767 51923
rect 44767 51901 44769 51923
rect 44713 51889 44769 51901
rect 44713 51867 44715 51889
rect 44715 51867 44767 51889
rect 44767 51867 44769 51889
rect 44713 51837 44715 51843
rect 44715 51837 44767 51843
rect 44767 51837 44769 51843
rect 44713 51825 44769 51837
rect 44713 51787 44715 51825
rect 44715 51787 44767 51825
rect 44767 51787 44769 51825
rect 44713 51761 44769 51763
rect 44713 51709 44715 51761
rect 44715 51709 44767 51761
rect 44767 51709 44769 51761
rect 44713 51707 44769 51709
rect 44720 51424 44776 51442
rect 44720 51386 44722 51424
rect 44722 51386 44774 51424
rect 44774 51386 44776 51424
rect 44720 51360 44776 51362
rect 44720 51308 44722 51360
rect 44722 51308 44774 51360
rect 44774 51308 44776 51360
rect 44720 51306 44776 51308
rect 44720 51244 44722 51282
rect 44722 51244 44774 51282
rect 44774 51244 44776 51282
rect 44720 51226 44776 51244
rect 44717 50479 44773 50481
rect 44717 50427 44719 50479
rect 44719 50427 44771 50479
rect 44771 50427 44773 50479
rect 44717 50425 44773 50427
rect 44717 50363 44719 50401
rect 44719 50363 44771 50401
rect 44771 50363 44773 50401
rect 44717 50351 44773 50363
rect 44717 50345 44719 50351
rect 44719 50345 44771 50351
rect 44771 50345 44773 50351
rect 44717 50299 44719 50321
rect 44719 50299 44771 50321
rect 44771 50299 44773 50321
rect 44717 50287 44773 50299
rect 44717 50265 44719 50287
rect 44719 50265 44771 50287
rect 44771 50265 44773 50287
rect 44717 50235 44719 50241
rect 44719 50235 44771 50241
rect 44771 50235 44773 50241
rect 44717 50223 44773 50235
rect 44717 50185 44719 50223
rect 44719 50185 44771 50223
rect 44771 50185 44773 50223
rect 44717 50159 44773 50161
rect 44717 50107 44719 50159
rect 44719 50107 44771 50159
rect 44771 50107 44773 50159
rect 44717 50105 44773 50107
rect 44713 49825 44769 49843
rect 44713 49787 44715 49825
rect 44715 49787 44767 49825
rect 44767 49787 44769 49825
rect 44713 49761 44769 49763
rect 44713 49709 44715 49761
rect 44715 49709 44767 49761
rect 44767 49709 44769 49761
rect 44713 49707 44769 49709
rect 31657 49472 31713 49498
rect 31657 49442 31659 49472
rect 31659 49442 31711 49472
rect 31711 49442 31713 49472
rect 31657 49408 31713 49418
rect 31657 49362 31659 49408
rect 31659 49362 31711 49408
rect 31711 49362 31713 49408
rect 31657 49292 31659 49338
rect 31659 49292 31711 49338
rect 31711 49292 31713 49338
rect 31657 49282 31713 49292
rect 31657 49228 31659 49258
rect 31659 49228 31711 49258
rect 31711 49228 31713 49258
rect 31657 49202 31713 49228
rect 16511 49165 16727 49183
rect 16511 48985 16529 49165
rect 16529 48985 16709 49165
rect 16709 48985 16727 49165
rect 16511 48967 16727 48985
rect 18949 47602 19005 47604
rect 19029 47602 19085 47604
rect 19109 47602 19165 47604
rect 19189 47602 19245 47604
rect 19269 47602 19325 47604
rect 19349 47602 19405 47604
rect 19429 47602 19485 47604
rect 19509 47602 19565 47604
rect 19589 47602 19645 47604
rect 19669 47602 19725 47604
rect 19749 47602 19805 47604
rect 19829 47602 19885 47604
rect 19909 47602 19965 47604
rect 19989 47602 20045 47604
rect 20069 47602 20125 47604
rect 20149 47602 20205 47604
rect 20229 47602 20285 47604
rect 20309 47602 20365 47604
rect 20389 47602 20445 47604
rect 20469 47602 20525 47604
rect 20549 47602 20605 47604
rect 20629 47602 20685 47604
rect 20709 47602 20765 47604
rect 20789 47602 20845 47604
rect 20869 47602 20925 47604
rect 20949 47602 21005 47604
rect 21029 47602 21085 47604
rect 21109 47602 21165 47604
rect 21189 47602 21245 47604
rect 21269 47602 21325 47604
rect 21349 47602 21405 47604
rect 21429 47602 21485 47604
rect 21509 47602 21565 47604
rect 21589 47602 21645 47604
rect 21669 47602 21725 47604
rect 21749 47602 21805 47604
rect 21829 47602 21885 47604
rect 21909 47602 21965 47604
rect 21989 47602 22045 47604
rect 22069 47602 22125 47604
rect 22149 47602 22205 47604
rect 18949 47550 18971 47602
rect 18971 47550 18983 47602
rect 18983 47550 19005 47602
rect 19029 47550 19035 47602
rect 19035 47550 19047 47602
rect 19047 47550 19085 47602
rect 19109 47550 19111 47602
rect 19111 47550 19163 47602
rect 19163 47550 19165 47602
rect 19189 47550 19227 47602
rect 19227 47550 19239 47602
rect 19239 47550 19245 47602
rect 19269 47550 19291 47602
rect 19291 47550 19303 47602
rect 19303 47550 19325 47602
rect 19349 47550 19355 47602
rect 19355 47550 19367 47602
rect 19367 47550 19405 47602
rect 19429 47550 19431 47602
rect 19431 47550 19483 47602
rect 19483 47550 19485 47602
rect 19509 47550 19547 47602
rect 19547 47550 19559 47602
rect 19559 47550 19565 47602
rect 19589 47550 19611 47602
rect 19611 47550 19623 47602
rect 19623 47550 19645 47602
rect 19669 47550 19675 47602
rect 19675 47550 19687 47602
rect 19687 47550 19725 47602
rect 19749 47550 19751 47602
rect 19751 47550 19803 47602
rect 19803 47550 19805 47602
rect 19829 47550 19867 47602
rect 19867 47550 19879 47602
rect 19879 47550 19885 47602
rect 19909 47550 19931 47602
rect 19931 47550 19943 47602
rect 19943 47550 19965 47602
rect 19989 47550 19995 47602
rect 19995 47550 20007 47602
rect 20007 47550 20045 47602
rect 20069 47550 20071 47602
rect 20071 47550 20123 47602
rect 20123 47550 20125 47602
rect 20149 47550 20187 47602
rect 20187 47550 20199 47602
rect 20199 47550 20205 47602
rect 20229 47550 20251 47602
rect 20251 47550 20263 47602
rect 20263 47550 20285 47602
rect 20309 47550 20315 47602
rect 20315 47550 20327 47602
rect 20327 47550 20365 47602
rect 20389 47550 20391 47602
rect 20391 47550 20443 47602
rect 20443 47550 20445 47602
rect 20469 47550 20507 47602
rect 20507 47550 20519 47602
rect 20519 47550 20525 47602
rect 20549 47550 20571 47602
rect 20571 47550 20583 47602
rect 20583 47550 20605 47602
rect 20629 47550 20635 47602
rect 20635 47550 20647 47602
rect 20647 47550 20685 47602
rect 20709 47550 20711 47602
rect 20711 47550 20763 47602
rect 20763 47550 20765 47602
rect 20789 47550 20827 47602
rect 20827 47550 20839 47602
rect 20839 47550 20845 47602
rect 20869 47550 20891 47602
rect 20891 47550 20903 47602
rect 20903 47550 20925 47602
rect 20949 47550 20955 47602
rect 20955 47550 20967 47602
rect 20967 47550 21005 47602
rect 21029 47550 21031 47602
rect 21031 47550 21083 47602
rect 21083 47550 21085 47602
rect 21109 47550 21147 47602
rect 21147 47550 21159 47602
rect 21159 47550 21165 47602
rect 21189 47550 21211 47602
rect 21211 47550 21223 47602
rect 21223 47550 21245 47602
rect 21269 47550 21275 47602
rect 21275 47550 21287 47602
rect 21287 47550 21325 47602
rect 21349 47550 21351 47602
rect 21351 47550 21403 47602
rect 21403 47550 21405 47602
rect 21429 47550 21467 47602
rect 21467 47550 21479 47602
rect 21479 47550 21485 47602
rect 21509 47550 21531 47602
rect 21531 47550 21543 47602
rect 21543 47550 21565 47602
rect 21589 47550 21595 47602
rect 21595 47550 21607 47602
rect 21607 47550 21645 47602
rect 21669 47550 21671 47602
rect 21671 47550 21723 47602
rect 21723 47550 21725 47602
rect 21749 47550 21787 47602
rect 21787 47550 21799 47602
rect 21799 47550 21805 47602
rect 21829 47550 21851 47602
rect 21851 47550 21863 47602
rect 21863 47550 21885 47602
rect 21909 47550 21915 47602
rect 21915 47550 21927 47602
rect 21927 47550 21965 47602
rect 21989 47550 21991 47602
rect 21991 47550 22043 47602
rect 22043 47550 22045 47602
rect 22069 47550 22107 47602
rect 22107 47550 22119 47602
rect 22119 47550 22125 47602
rect 22149 47550 22171 47602
rect 22171 47550 22183 47602
rect 22183 47550 22205 47602
rect 18949 47548 19005 47550
rect 19029 47548 19085 47550
rect 19109 47548 19165 47550
rect 19189 47548 19245 47550
rect 19269 47548 19325 47550
rect 19349 47548 19405 47550
rect 19429 47548 19485 47550
rect 19509 47548 19565 47550
rect 19589 47548 19645 47550
rect 19669 47548 19725 47550
rect 19749 47548 19805 47550
rect 19829 47548 19885 47550
rect 19909 47548 19965 47550
rect 19989 47548 20045 47550
rect 20069 47548 20125 47550
rect 20149 47548 20205 47550
rect 20229 47548 20285 47550
rect 20309 47548 20365 47550
rect 20389 47548 20445 47550
rect 20469 47548 20525 47550
rect 20549 47548 20605 47550
rect 20629 47548 20685 47550
rect 20709 47548 20765 47550
rect 20789 47548 20845 47550
rect 20869 47548 20925 47550
rect 20949 47548 21005 47550
rect 21029 47548 21085 47550
rect 21109 47548 21165 47550
rect 21189 47548 21245 47550
rect 21269 47548 21325 47550
rect 21349 47548 21405 47550
rect 21429 47548 21485 47550
rect 21509 47548 21565 47550
rect 21589 47548 21645 47550
rect 21669 47548 21725 47550
rect 21749 47548 21805 47550
rect 21829 47548 21885 47550
rect 21909 47548 21965 47550
rect 21989 47548 22045 47550
rect 22069 47548 22125 47550
rect 22149 47548 22205 47550
rect 18951 43074 19007 43076
rect 19031 43074 19087 43076
rect 19111 43074 19167 43076
rect 19191 43074 19247 43076
rect 19271 43074 19327 43076
rect 19351 43074 19407 43076
rect 19431 43074 19487 43076
rect 19511 43074 19567 43076
rect 19591 43074 19647 43076
rect 19671 43074 19727 43076
rect 19751 43074 19807 43076
rect 19831 43074 19887 43076
rect 19911 43074 19967 43076
rect 19991 43074 20047 43076
rect 20071 43074 20127 43076
rect 20151 43074 20207 43076
rect 20231 43074 20287 43076
rect 20311 43074 20367 43076
rect 20391 43074 20447 43076
rect 20471 43074 20527 43076
rect 20551 43074 20607 43076
rect 20631 43074 20687 43076
rect 20711 43074 20767 43076
rect 20791 43074 20847 43076
rect 20871 43074 20927 43076
rect 20951 43074 21007 43076
rect 21031 43074 21087 43076
rect 21111 43074 21167 43076
rect 21191 43074 21247 43076
rect 21271 43074 21327 43076
rect 21351 43074 21407 43076
rect 21431 43074 21487 43076
rect 21511 43074 21567 43076
rect 21591 43074 21647 43076
rect 21671 43074 21727 43076
rect 21751 43074 21807 43076
rect 21831 43074 21887 43076
rect 21911 43074 21967 43076
rect 21991 43074 22047 43076
rect 22071 43074 22127 43076
rect 22151 43074 22207 43076
rect 18951 43022 18953 43074
rect 18953 43022 19005 43074
rect 19005 43022 19007 43074
rect 19031 43022 19069 43074
rect 19069 43022 19081 43074
rect 19081 43022 19087 43074
rect 19111 43022 19133 43074
rect 19133 43022 19145 43074
rect 19145 43022 19167 43074
rect 19191 43022 19197 43074
rect 19197 43022 19209 43074
rect 19209 43022 19247 43074
rect 19271 43022 19273 43074
rect 19273 43022 19325 43074
rect 19325 43022 19327 43074
rect 19351 43022 19389 43074
rect 19389 43022 19401 43074
rect 19401 43022 19407 43074
rect 19431 43022 19453 43074
rect 19453 43022 19465 43074
rect 19465 43022 19487 43074
rect 19511 43022 19517 43074
rect 19517 43022 19529 43074
rect 19529 43022 19567 43074
rect 19591 43022 19593 43074
rect 19593 43022 19645 43074
rect 19645 43022 19647 43074
rect 19671 43022 19709 43074
rect 19709 43022 19721 43074
rect 19721 43022 19727 43074
rect 19751 43022 19773 43074
rect 19773 43022 19785 43074
rect 19785 43022 19807 43074
rect 19831 43022 19837 43074
rect 19837 43022 19849 43074
rect 19849 43022 19887 43074
rect 19911 43022 19913 43074
rect 19913 43022 19965 43074
rect 19965 43022 19967 43074
rect 19991 43022 20029 43074
rect 20029 43022 20041 43074
rect 20041 43022 20047 43074
rect 20071 43022 20093 43074
rect 20093 43022 20105 43074
rect 20105 43022 20127 43074
rect 20151 43022 20157 43074
rect 20157 43022 20169 43074
rect 20169 43022 20207 43074
rect 20231 43022 20233 43074
rect 20233 43022 20285 43074
rect 20285 43022 20287 43074
rect 20311 43022 20349 43074
rect 20349 43022 20361 43074
rect 20361 43022 20367 43074
rect 20391 43022 20413 43074
rect 20413 43022 20425 43074
rect 20425 43022 20447 43074
rect 20471 43022 20477 43074
rect 20477 43022 20489 43074
rect 20489 43022 20527 43074
rect 20551 43022 20553 43074
rect 20553 43022 20605 43074
rect 20605 43022 20607 43074
rect 20631 43022 20669 43074
rect 20669 43022 20681 43074
rect 20681 43022 20687 43074
rect 20711 43022 20733 43074
rect 20733 43022 20745 43074
rect 20745 43022 20767 43074
rect 20791 43022 20797 43074
rect 20797 43022 20809 43074
rect 20809 43022 20847 43074
rect 20871 43022 20873 43074
rect 20873 43022 20925 43074
rect 20925 43022 20927 43074
rect 20951 43022 20989 43074
rect 20989 43022 21001 43074
rect 21001 43022 21007 43074
rect 21031 43022 21053 43074
rect 21053 43022 21065 43074
rect 21065 43022 21087 43074
rect 21111 43022 21117 43074
rect 21117 43022 21129 43074
rect 21129 43022 21167 43074
rect 21191 43022 21193 43074
rect 21193 43022 21245 43074
rect 21245 43022 21247 43074
rect 21271 43022 21309 43074
rect 21309 43022 21321 43074
rect 21321 43022 21327 43074
rect 21351 43022 21373 43074
rect 21373 43022 21385 43074
rect 21385 43022 21407 43074
rect 21431 43022 21437 43074
rect 21437 43022 21449 43074
rect 21449 43022 21487 43074
rect 21511 43022 21513 43074
rect 21513 43022 21565 43074
rect 21565 43022 21567 43074
rect 21591 43022 21629 43074
rect 21629 43022 21641 43074
rect 21641 43022 21647 43074
rect 21671 43022 21693 43074
rect 21693 43022 21705 43074
rect 21705 43022 21727 43074
rect 21751 43022 21757 43074
rect 21757 43022 21769 43074
rect 21769 43022 21807 43074
rect 21831 43022 21833 43074
rect 21833 43022 21885 43074
rect 21885 43022 21887 43074
rect 21911 43022 21949 43074
rect 21949 43022 21961 43074
rect 21961 43022 21967 43074
rect 21991 43022 22013 43074
rect 22013 43022 22025 43074
rect 22025 43022 22047 43074
rect 22071 43022 22077 43074
rect 22077 43022 22089 43074
rect 22089 43022 22127 43074
rect 22151 43022 22153 43074
rect 22153 43022 22205 43074
rect 22205 43022 22207 43074
rect 18951 43020 19007 43022
rect 19031 43020 19087 43022
rect 19111 43020 19167 43022
rect 19191 43020 19247 43022
rect 19271 43020 19327 43022
rect 19351 43020 19407 43022
rect 19431 43020 19487 43022
rect 19511 43020 19567 43022
rect 19591 43020 19647 43022
rect 19671 43020 19727 43022
rect 19751 43020 19807 43022
rect 19831 43020 19887 43022
rect 19911 43020 19967 43022
rect 19991 43020 20047 43022
rect 20071 43020 20127 43022
rect 20151 43020 20207 43022
rect 20231 43020 20287 43022
rect 20311 43020 20367 43022
rect 20391 43020 20447 43022
rect 20471 43020 20527 43022
rect 20551 43020 20607 43022
rect 20631 43020 20687 43022
rect 20711 43020 20767 43022
rect 20791 43020 20847 43022
rect 20871 43020 20927 43022
rect 20951 43020 21007 43022
rect 21031 43020 21087 43022
rect 21111 43020 21167 43022
rect 21191 43020 21247 43022
rect 21271 43020 21327 43022
rect 21351 43020 21407 43022
rect 21431 43020 21487 43022
rect 21511 43020 21567 43022
rect 21591 43020 21647 43022
rect 21671 43020 21727 43022
rect 21751 43020 21807 43022
rect 21831 43020 21887 43022
rect 21911 43020 21967 43022
rect 21991 43020 22047 43022
rect 22071 43020 22127 43022
rect 22151 43020 22207 43022
rect 16508 41624 16724 41642
rect 16508 41444 16526 41624
rect 16526 41444 16706 41624
rect 16706 41444 16724 41624
rect 16508 41426 16724 41444
rect 18953 40079 19009 40081
rect 19033 40079 19089 40081
rect 19113 40079 19169 40081
rect 19193 40079 19249 40081
rect 19273 40079 19329 40081
rect 19353 40079 19409 40081
rect 19433 40079 19489 40081
rect 19513 40079 19569 40081
rect 19593 40079 19649 40081
rect 19673 40079 19729 40081
rect 19753 40079 19809 40081
rect 19833 40079 19889 40081
rect 19913 40079 19969 40081
rect 19993 40079 20049 40081
rect 20073 40079 20129 40081
rect 20153 40079 20209 40081
rect 20233 40079 20289 40081
rect 20313 40079 20369 40081
rect 20393 40079 20449 40081
rect 20473 40079 20529 40081
rect 20553 40079 20609 40081
rect 20633 40079 20689 40081
rect 20713 40079 20769 40081
rect 20793 40079 20849 40081
rect 20873 40079 20929 40081
rect 20953 40079 21009 40081
rect 21033 40079 21089 40081
rect 21113 40079 21169 40081
rect 21193 40079 21249 40081
rect 21273 40079 21329 40081
rect 21353 40079 21409 40081
rect 21433 40079 21489 40081
rect 21513 40079 21569 40081
rect 21593 40079 21649 40081
rect 21673 40079 21729 40081
rect 21753 40079 21809 40081
rect 21833 40079 21889 40081
rect 21913 40079 21969 40081
rect 21993 40079 22049 40081
rect 22073 40079 22129 40081
rect 22153 40079 22209 40081
rect 18953 40027 18975 40079
rect 18975 40027 18987 40079
rect 18987 40027 19009 40079
rect 19033 40027 19039 40079
rect 19039 40027 19051 40079
rect 19051 40027 19089 40079
rect 19113 40027 19115 40079
rect 19115 40027 19167 40079
rect 19167 40027 19169 40079
rect 19193 40027 19231 40079
rect 19231 40027 19243 40079
rect 19243 40027 19249 40079
rect 19273 40027 19295 40079
rect 19295 40027 19307 40079
rect 19307 40027 19329 40079
rect 19353 40027 19359 40079
rect 19359 40027 19371 40079
rect 19371 40027 19409 40079
rect 19433 40027 19435 40079
rect 19435 40027 19487 40079
rect 19487 40027 19489 40079
rect 19513 40027 19551 40079
rect 19551 40027 19563 40079
rect 19563 40027 19569 40079
rect 19593 40027 19615 40079
rect 19615 40027 19627 40079
rect 19627 40027 19649 40079
rect 19673 40027 19679 40079
rect 19679 40027 19691 40079
rect 19691 40027 19729 40079
rect 19753 40027 19755 40079
rect 19755 40027 19807 40079
rect 19807 40027 19809 40079
rect 19833 40027 19871 40079
rect 19871 40027 19883 40079
rect 19883 40027 19889 40079
rect 19913 40027 19935 40079
rect 19935 40027 19947 40079
rect 19947 40027 19969 40079
rect 19993 40027 19999 40079
rect 19999 40027 20011 40079
rect 20011 40027 20049 40079
rect 20073 40027 20075 40079
rect 20075 40027 20127 40079
rect 20127 40027 20129 40079
rect 20153 40027 20191 40079
rect 20191 40027 20203 40079
rect 20203 40027 20209 40079
rect 20233 40027 20255 40079
rect 20255 40027 20267 40079
rect 20267 40027 20289 40079
rect 20313 40027 20319 40079
rect 20319 40027 20331 40079
rect 20331 40027 20369 40079
rect 20393 40027 20395 40079
rect 20395 40027 20447 40079
rect 20447 40027 20449 40079
rect 20473 40027 20511 40079
rect 20511 40027 20523 40079
rect 20523 40027 20529 40079
rect 20553 40027 20575 40079
rect 20575 40027 20587 40079
rect 20587 40027 20609 40079
rect 20633 40027 20639 40079
rect 20639 40027 20651 40079
rect 20651 40027 20689 40079
rect 20713 40027 20715 40079
rect 20715 40027 20767 40079
rect 20767 40027 20769 40079
rect 20793 40027 20831 40079
rect 20831 40027 20843 40079
rect 20843 40027 20849 40079
rect 20873 40027 20895 40079
rect 20895 40027 20907 40079
rect 20907 40027 20929 40079
rect 20953 40027 20959 40079
rect 20959 40027 20971 40079
rect 20971 40027 21009 40079
rect 21033 40027 21035 40079
rect 21035 40027 21087 40079
rect 21087 40027 21089 40079
rect 21113 40027 21151 40079
rect 21151 40027 21163 40079
rect 21163 40027 21169 40079
rect 21193 40027 21215 40079
rect 21215 40027 21227 40079
rect 21227 40027 21249 40079
rect 21273 40027 21279 40079
rect 21279 40027 21291 40079
rect 21291 40027 21329 40079
rect 21353 40027 21355 40079
rect 21355 40027 21407 40079
rect 21407 40027 21409 40079
rect 21433 40027 21471 40079
rect 21471 40027 21483 40079
rect 21483 40027 21489 40079
rect 21513 40027 21535 40079
rect 21535 40027 21547 40079
rect 21547 40027 21569 40079
rect 21593 40027 21599 40079
rect 21599 40027 21611 40079
rect 21611 40027 21649 40079
rect 21673 40027 21675 40079
rect 21675 40027 21727 40079
rect 21727 40027 21729 40079
rect 21753 40027 21791 40079
rect 21791 40027 21803 40079
rect 21803 40027 21809 40079
rect 21833 40027 21855 40079
rect 21855 40027 21867 40079
rect 21867 40027 21889 40079
rect 21913 40027 21919 40079
rect 21919 40027 21931 40079
rect 21931 40027 21969 40079
rect 21993 40027 21995 40079
rect 21995 40027 22047 40079
rect 22047 40027 22049 40079
rect 22073 40027 22111 40079
rect 22111 40027 22123 40079
rect 22123 40027 22129 40079
rect 22153 40027 22175 40079
rect 22175 40027 22187 40079
rect 22187 40027 22209 40079
rect 18953 40025 19009 40027
rect 19033 40025 19089 40027
rect 19113 40025 19169 40027
rect 19193 40025 19249 40027
rect 19273 40025 19329 40027
rect 19353 40025 19409 40027
rect 19433 40025 19489 40027
rect 19513 40025 19569 40027
rect 19593 40025 19649 40027
rect 19673 40025 19729 40027
rect 19753 40025 19809 40027
rect 19833 40025 19889 40027
rect 19913 40025 19969 40027
rect 19993 40025 20049 40027
rect 20073 40025 20129 40027
rect 20153 40025 20209 40027
rect 20233 40025 20289 40027
rect 20313 40025 20369 40027
rect 20393 40025 20449 40027
rect 20473 40025 20529 40027
rect 20553 40025 20609 40027
rect 20633 40025 20689 40027
rect 20713 40025 20769 40027
rect 20793 40025 20849 40027
rect 20873 40025 20929 40027
rect 20953 40025 21009 40027
rect 21033 40025 21089 40027
rect 21113 40025 21169 40027
rect 21193 40025 21249 40027
rect 21273 40025 21329 40027
rect 21353 40025 21409 40027
rect 21433 40025 21489 40027
rect 21513 40025 21569 40027
rect 21593 40025 21649 40027
rect 21673 40025 21729 40027
rect 21753 40025 21809 40027
rect 21833 40025 21889 40027
rect 21913 40025 21969 40027
rect 21993 40025 22049 40027
rect 22073 40025 22129 40027
rect 22153 40025 22209 40027
rect 31657 48941 31713 48959
rect 31657 48903 31659 48941
rect 31659 48903 31711 48941
rect 31711 48903 31713 48941
rect 31657 48877 31713 48879
rect 31657 48825 31659 48877
rect 31659 48825 31711 48877
rect 31711 48825 31713 48877
rect 31657 48823 31713 48825
rect 31657 48761 31659 48799
rect 31659 48761 31711 48799
rect 31711 48761 31713 48799
rect 31657 48743 31713 48761
rect 41386 49440 41442 49442
rect 41386 49388 41388 49440
rect 41388 49388 41440 49440
rect 41440 49388 41442 49440
rect 41386 49386 41442 49388
rect 41386 49324 41388 49362
rect 41388 49324 41440 49362
rect 41440 49324 41442 49362
rect 41386 49312 41442 49324
rect 41386 49306 41388 49312
rect 41388 49306 41440 49312
rect 41440 49306 41442 49312
rect 41386 49260 41388 49282
rect 41388 49260 41440 49282
rect 41440 49260 41442 49282
rect 41386 49248 41442 49260
rect 41386 49226 41388 49248
rect 41388 49226 41440 49248
rect 41440 49226 41442 49248
rect 41386 49196 41388 49202
rect 41388 49196 41440 49202
rect 41440 49196 41442 49202
rect 41386 49184 41442 49196
rect 41386 49146 41388 49184
rect 41388 49146 41440 49184
rect 41440 49146 41442 49184
rect 41386 49120 41442 49122
rect 41386 49068 41388 49120
rect 41388 49068 41440 49120
rect 41440 49068 41442 49120
rect 41386 49066 41442 49068
rect 39495 48932 39551 48988
rect 43109 49626 43165 49682
rect 44713 49645 44715 49683
rect 44715 49645 44767 49683
rect 44767 49645 44769 49683
rect 44713 49627 44769 49645
rect 42688 48834 42744 48890
rect 39495 47703 39551 47759
rect 41374 47633 41430 47651
rect 41374 47595 41376 47633
rect 41376 47595 41428 47633
rect 41428 47595 41430 47633
rect 41374 47569 41430 47571
rect 41374 47517 41376 47569
rect 41376 47517 41428 47569
rect 41428 47517 41430 47569
rect 41374 47515 41430 47517
rect 41374 47453 41376 47491
rect 41376 47453 41428 47491
rect 41428 47453 41430 47491
rect 41374 47435 41430 47453
rect 44705 48677 44707 48715
rect 44707 48677 44759 48715
rect 44759 48677 44761 48715
rect 44705 48665 44761 48677
rect 44705 48659 44707 48665
rect 44707 48659 44759 48665
rect 44759 48659 44761 48665
rect 44705 48613 44707 48635
rect 44707 48613 44759 48635
rect 44759 48613 44761 48635
rect 44705 48601 44761 48613
rect 44705 48579 44707 48601
rect 44707 48579 44759 48601
rect 44759 48579 44761 48601
rect 44705 48549 44707 48555
rect 44707 48549 44759 48555
rect 44759 48549 44761 48555
rect 44705 48537 44761 48549
rect 44705 48499 44707 48537
rect 44707 48499 44759 48537
rect 44759 48499 44761 48537
rect 44709 48233 44765 48251
rect 44709 48195 44711 48233
rect 44711 48195 44763 48233
rect 44763 48195 44765 48233
rect 44709 48169 44765 48171
rect 44709 48117 44711 48169
rect 44711 48117 44763 48169
rect 44763 48117 44765 48169
rect 44709 48115 44765 48117
rect 44709 48053 44711 48091
rect 44711 48053 44763 48091
rect 44763 48053 44765 48091
rect 44709 48035 44765 48053
rect 44712 47275 44768 47277
rect 44712 47223 44714 47275
rect 44714 47223 44766 47275
rect 44766 47223 44768 47275
rect 44712 47221 44768 47223
rect 44712 47159 44714 47197
rect 44714 47159 44766 47197
rect 44766 47159 44768 47197
rect 44712 47147 44768 47159
rect 44712 47141 44714 47147
rect 44714 47141 44766 47147
rect 44766 47141 44768 47147
rect 44712 47095 44714 47117
rect 44714 47095 44766 47117
rect 44766 47095 44768 47117
rect 44712 47083 44768 47095
rect 44712 47061 44714 47083
rect 44714 47061 44766 47083
rect 44766 47061 44768 47083
rect 44712 47031 44714 47037
rect 44714 47031 44766 47037
rect 44766 47031 44768 47037
rect 44712 47019 44768 47031
rect 44712 46981 44714 47019
rect 44714 46981 44766 47019
rect 44766 46981 44768 47019
rect 44712 46955 44768 46957
rect 44712 46903 44714 46955
rect 44714 46903 44766 46955
rect 44766 46903 44768 46955
rect 44712 46901 44768 46903
rect 44709 46623 44765 46641
rect 44709 46585 44711 46623
rect 44711 46585 44763 46623
rect 44763 46585 44765 46623
rect 44709 46559 44765 46561
rect 44709 46507 44711 46559
rect 44711 46507 44763 46559
rect 44763 46507 44765 46559
rect 44709 46505 44765 46507
rect 44709 46443 44711 46481
rect 44711 46443 44763 46481
rect 44763 46443 44765 46481
rect 44709 46425 44765 46443
rect 31646 41866 31648 41904
rect 31648 41866 31700 41904
rect 31700 41866 31702 41904
rect 31646 41854 31702 41866
rect 31646 41848 31648 41854
rect 31648 41848 31700 41854
rect 31700 41848 31702 41854
rect 31646 41802 31648 41824
rect 31648 41802 31700 41824
rect 31700 41802 31702 41824
rect 31646 41790 31702 41802
rect 31646 41768 31648 41790
rect 31648 41768 31700 41790
rect 31700 41768 31702 41790
rect 31646 41738 31648 41744
rect 31648 41738 31700 41744
rect 31700 41738 31702 41744
rect 31646 41726 31702 41738
rect 31646 41688 31648 41726
rect 31648 41688 31700 41726
rect 31700 41688 31702 41726
rect 31652 41398 31708 41416
rect 31652 41360 31654 41398
rect 31654 41360 31706 41398
rect 31706 41360 31708 41398
rect 31652 41334 31708 41336
rect 31652 41282 31654 41334
rect 31654 41282 31706 41334
rect 31706 41282 31708 41334
rect 31652 41280 31708 41282
rect 31652 41218 31654 41256
rect 31654 41218 31706 41256
rect 31706 41218 31708 41256
rect 31652 41200 31708 41218
rect 32928 40211 32984 40267
rect 29178 39403 29234 39459
rect 31585 38393 31587 38431
rect 31587 38393 31639 38431
rect 31639 38393 31641 38431
rect 31585 38381 31641 38393
rect 31585 38375 31587 38381
rect 31587 38375 31639 38381
rect 31639 38375 31641 38381
rect 31585 38329 31587 38351
rect 31587 38329 31639 38351
rect 31639 38329 31641 38351
rect 31585 38317 31641 38329
rect 31585 38295 31587 38317
rect 31587 38295 31639 38317
rect 31639 38295 31641 38317
rect 31585 38265 31587 38271
rect 31587 38265 31639 38271
rect 31639 38265 31641 38271
rect 31585 38253 31641 38265
rect 31585 38215 31587 38253
rect 31587 38215 31639 38253
rect 31639 38215 31641 38253
rect 31584 37919 31640 37937
rect 31584 37881 31586 37919
rect 31586 37881 31638 37919
rect 31638 37881 31640 37919
rect 31584 37855 31640 37857
rect 31584 37803 31586 37855
rect 31586 37803 31638 37855
rect 31638 37803 31640 37855
rect 31584 37801 31640 37803
rect 31584 37739 31586 37777
rect 31586 37739 31638 37777
rect 31638 37739 31640 37777
rect 31584 37721 31640 37739
rect 38875 38089 38931 38091
rect 38875 38037 38877 38089
rect 38877 38037 38929 38089
rect 38929 38037 38931 38089
rect 38875 38035 38931 38037
rect 61426 52557 61482 52613
rect 65436 52554 65492 52610
rect 51819 51494 51875 51550
rect 53180 50817 53236 50873
rect 76969 49971 77025 50027
rect 76971 49560 77027 49616
rect 62815 48598 62871 48600
rect 62815 48546 62817 48598
rect 62817 48546 62869 48598
rect 62869 48546 62871 48598
rect 62815 48544 62871 48546
rect 64166 48554 64222 48610
rect 62815 48482 62817 48520
rect 62817 48482 62869 48520
rect 62869 48482 62871 48520
rect 62815 48470 62871 48482
rect 62815 48464 62817 48470
rect 62817 48464 62869 48470
rect 62869 48464 62871 48470
rect 62815 48418 62817 48440
rect 62817 48418 62869 48440
rect 62869 48418 62871 48440
rect 62815 48406 62871 48418
rect 62815 48384 62817 48406
rect 62817 48384 62869 48406
rect 62869 48384 62871 48406
rect 62815 48354 62817 48360
rect 62817 48354 62869 48360
rect 62869 48354 62871 48360
rect 62815 48342 62871 48354
rect 62815 48304 62817 48342
rect 62817 48304 62869 48342
rect 62869 48304 62871 48342
rect 62815 48278 62871 48280
rect 62815 48226 62817 48278
rect 62817 48226 62869 48278
rect 62869 48226 62871 48278
rect 62815 48224 62871 48226
rect 99989 48167 100045 48169
rect 100069 48167 100125 48169
rect 100149 48167 100205 48169
rect 100229 48167 100285 48169
rect 100309 48167 100365 48169
rect 100389 48167 100445 48169
rect 100469 48167 100525 48169
rect 100549 48167 100605 48169
rect 100629 48167 100685 48169
rect 100709 48167 100765 48169
rect 100789 48167 100845 48169
rect 100869 48167 100925 48169
rect 100949 48167 101005 48169
rect 101029 48167 101085 48169
rect 101109 48167 101165 48169
rect 101189 48167 101245 48169
rect 101269 48167 101325 48169
rect 101349 48167 101405 48169
rect 101429 48167 101485 48169
rect 101509 48167 101565 48169
rect 101589 48167 101645 48169
rect 101669 48167 101725 48169
rect 101749 48167 101805 48169
rect 101829 48167 101885 48169
rect 101909 48167 101965 48169
rect 101989 48167 102045 48169
rect 102069 48167 102125 48169
rect 102149 48167 102205 48169
rect 102229 48167 102285 48169
rect 102309 48167 102365 48169
rect 102389 48167 102445 48169
rect 102469 48167 102525 48169
rect 102549 48167 102605 48169
rect 102629 48167 102685 48169
rect 102709 48167 102765 48169
rect 102789 48167 102845 48169
rect 102869 48167 102925 48169
rect 102949 48167 103005 48169
rect 103029 48167 103085 48169
rect 103109 48167 103165 48169
rect 103189 48167 103245 48169
rect 99989 48115 100011 48167
rect 100011 48115 100023 48167
rect 100023 48115 100045 48167
rect 100069 48115 100075 48167
rect 100075 48115 100087 48167
rect 100087 48115 100125 48167
rect 100149 48115 100151 48167
rect 100151 48115 100203 48167
rect 100203 48115 100205 48167
rect 100229 48115 100267 48167
rect 100267 48115 100279 48167
rect 100279 48115 100285 48167
rect 100309 48115 100331 48167
rect 100331 48115 100343 48167
rect 100343 48115 100365 48167
rect 100389 48115 100395 48167
rect 100395 48115 100407 48167
rect 100407 48115 100445 48167
rect 100469 48115 100471 48167
rect 100471 48115 100523 48167
rect 100523 48115 100525 48167
rect 100549 48115 100587 48167
rect 100587 48115 100599 48167
rect 100599 48115 100605 48167
rect 100629 48115 100651 48167
rect 100651 48115 100663 48167
rect 100663 48115 100685 48167
rect 100709 48115 100715 48167
rect 100715 48115 100727 48167
rect 100727 48115 100765 48167
rect 100789 48115 100791 48167
rect 100791 48115 100843 48167
rect 100843 48115 100845 48167
rect 100869 48115 100907 48167
rect 100907 48115 100919 48167
rect 100919 48115 100925 48167
rect 100949 48115 100971 48167
rect 100971 48115 100983 48167
rect 100983 48115 101005 48167
rect 101029 48115 101035 48167
rect 101035 48115 101047 48167
rect 101047 48115 101085 48167
rect 101109 48115 101111 48167
rect 101111 48115 101163 48167
rect 101163 48115 101165 48167
rect 101189 48115 101227 48167
rect 101227 48115 101239 48167
rect 101239 48115 101245 48167
rect 101269 48115 101291 48167
rect 101291 48115 101303 48167
rect 101303 48115 101325 48167
rect 101349 48115 101355 48167
rect 101355 48115 101367 48167
rect 101367 48115 101405 48167
rect 101429 48115 101431 48167
rect 101431 48115 101483 48167
rect 101483 48115 101485 48167
rect 101509 48115 101547 48167
rect 101547 48115 101559 48167
rect 101559 48115 101565 48167
rect 101589 48115 101611 48167
rect 101611 48115 101623 48167
rect 101623 48115 101645 48167
rect 101669 48115 101675 48167
rect 101675 48115 101687 48167
rect 101687 48115 101725 48167
rect 101749 48115 101751 48167
rect 101751 48115 101803 48167
rect 101803 48115 101805 48167
rect 101829 48115 101867 48167
rect 101867 48115 101879 48167
rect 101879 48115 101885 48167
rect 101909 48115 101931 48167
rect 101931 48115 101943 48167
rect 101943 48115 101965 48167
rect 101989 48115 101995 48167
rect 101995 48115 102007 48167
rect 102007 48115 102045 48167
rect 102069 48115 102071 48167
rect 102071 48115 102123 48167
rect 102123 48115 102125 48167
rect 102149 48115 102187 48167
rect 102187 48115 102199 48167
rect 102199 48115 102205 48167
rect 102229 48115 102251 48167
rect 102251 48115 102263 48167
rect 102263 48115 102285 48167
rect 102309 48115 102315 48167
rect 102315 48115 102327 48167
rect 102327 48115 102365 48167
rect 102389 48115 102391 48167
rect 102391 48115 102443 48167
rect 102443 48115 102445 48167
rect 102469 48115 102507 48167
rect 102507 48115 102519 48167
rect 102519 48115 102525 48167
rect 102549 48115 102571 48167
rect 102571 48115 102583 48167
rect 102583 48115 102605 48167
rect 102629 48115 102635 48167
rect 102635 48115 102647 48167
rect 102647 48115 102685 48167
rect 102709 48115 102711 48167
rect 102711 48115 102763 48167
rect 102763 48115 102765 48167
rect 102789 48115 102827 48167
rect 102827 48115 102839 48167
rect 102839 48115 102845 48167
rect 102869 48115 102891 48167
rect 102891 48115 102903 48167
rect 102903 48115 102925 48167
rect 102949 48115 102955 48167
rect 102955 48115 102967 48167
rect 102967 48115 103005 48167
rect 103029 48115 103031 48167
rect 103031 48115 103083 48167
rect 103083 48115 103085 48167
rect 103109 48115 103147 48167
rect 103147 48115 103159 48167
rect 103159 48115 103165 48167
rect 103189 48115 103211 48167
rect 103211 48115 103223 48167
rect 103223 48115 103245 48167
rect 99989 48113 100045 48115
rect 100069 48113 100125 48115
rect 100149 48113 100205 48115
rect 100229 48113 100285 48115
rect 100309 48113 100365 48115
rect 100389 48113 100445 48115
rect 100469 48113 100525 48115
rect 100549 48113 100605 48115
rect 100629 48113 100685 48115
rect 100709 48113 100765 48115
rect 100789 48113 100845 48115
rect 100869 48113 100925 48115
rect 100949 48113 101005 48115
rect 101029 48113 101085 48115
rect 101109 48113 101165 48115
rect 101189 48113 101245 48115
rect 101269 48113 101325 48115
rect 101349 48113 101405 48115
rect 101429 48113 101485 48115
rect 101509 48113 101565 48115
rect 101589 48113 101645 48115
rect 101669 48113 101725 48115
rect 101749 48113 101805 48115
rect 101829 48113 101885 48115
rect 101909 48113 101965 48115
rect 101989 48113 102045 48115
rect 102069 48113 102125 48115
rect 102149 48113 102205 48115
rect 102229 48113 102285 48115
rect 102309 48113 102365 48115
rect 102389 48113 102445 48115
rect 102469 48113 102525 48115
rect 102549 48113 102605 48115
rect 102629 48113 102685 48115
rect 102709 48113 102765 48115
rect 102789 48113 102845 48115
rect 102869 48113 102925 48115
rect 102949 48113 103005 48115
rect 103029 48113 103085 48115
rect 103109 48113 103165 48115
rect 103189 48113 103245 48115
rect 93164 47980 93220 48036
rect 92250 47882 92306 47884
rect 92250 47830 92252 47882
rect 92252 47830 92304 47882
rect 92304 47830 92306 47882
rect 92250 47828 92306 47830
rect 64189 47614 64245 47670
rect 96449 47715 96505 47733
rect 96449 47677 96451 47715
rect 96451 47677 96503 47715
rect 96503 47677 96505 47715
rect 94921 47579 94923 47601
rect 94923 47579 94975 47601
rect 94975 47579 94977 47601
rect 94921 47567 94977 47579
rect 94921 47545 94923 47567
rect 94923 47545 94975 47567
rect 94975 47545 94977 47567
rect 96449 47651 96505 47653
rect 96449 47599 96451 47651
rect 96451 47599 96503 47651
rect 96503 47599 96505 47651
rect 96449 47597 96505 47599
rect 96449 47535 96451 47573
rect 96451 47535 96503 47573
rect 96503 47535 96505 47573
rect 96449 47517 96505 47535
rect 65891 47349 65947 47351
rect 65971 47349 66027 47351
rect 65891 47297 65901 47349
rect 65901 47297 65947 47349
rect 65971 47297 66017 47349
rect 66017 47297 66027 47349
rect 65891 47295 65947 47297
rect 65971 47295 66027 47297
rect 94928 47162 94930 47200
rect 94930 47162 94982 47200
rect 94982 47162 94984 47200
rect 94928 47150 94984 47162
rect 94928 47144 94930 47150
rect 94930 47144 94982 47150
rect 94982 47144 94984 47150
rect 59648 47079 59704 47081
rect 59648 47027 59650 47079
rect 59650 47027 59702 47079
rect 59702 47027 59704 47079
rect 59648 47025 59704 47027
rect 67300 47079 67356 47081
rect 67300 47027 67302 47079
rect 67302 47027 67354 47079
rect 67354 47027 67356 47079
rect 67300 47025 67356 47027
rect 94928 47098 94930 47120
rect 94930 47098 94982 47120
rect 94982 47098 94984 47120
rect 94928 47086 94984 47098
rect 94928 47064 94930 47086
rect 94930 47064 94982 47086
rect 94982 47064 94984 47086
rect 94928 47034 94930 47040
rect 94930 47034 94982 47040
rect 94982 47034 94984 47040
rect 94928 47022 94984 47034
rect 94928 46984 94930 47022
rect 94930 46984 94982 47022
rect 94982 46984 94984 47022
rect 96444 47168 96446 47206
rect 96446 47168 96498 47206
rect 96498 47168 96500 47206
rect 96444 47156 96500 47168
rect 96444 47150 96446 47156
rect 96446 47150 96498 47156
rect 96498 47150 96500 47156
rect 96444 47104 96446 47126
rect 96446 47104 96498 47126
rect 96498 47104 96500 47126
rect 96444 47092 96500 47104
rect 96444 47070 96446 47092
rect 96446 47070 96498 47092
rect 96498 47070 96500 47092
rect 96444 47040 96446 47046
rect 96446 47040 96498 47046
rect 96498 47040 96500 47046
rect 96444 47028 96500 47040
rect 96444 46990 96446 47028
rect 96446 46990 96498 47028
rect 96498 46990 96500 47028
rect 92216 46654 92352 46790
rect 92876 46747 92932 46749
rect 92956 46747 93012 46749
rect 93036 46747 93092 46749
rect 92876 46695 92914 46747
rect 92914 46695 92926 46747
rect 92926 46695 92932 46747
rect 92956 46695 92978 46747
rect 92978 46695 92990 46747
rect 92990 46695 93012 46747
rect 93036 46695 93042 46747
rect 93042 46695 93054 46747
rect 93054 46695 93092 46747
rect 92876 46693 92932 46695
rect 92956 46693 93012 46695
rect 93036 46693 93092 46695
rect 104660 46728 104876 46746
rect 104660 46548 104678 46728
rect 104678 46548 104858 46728
rect 104858 46548 104876 46728
rect 104660 46530 104876 46548
rect 96449 46389 96505 46407
rect 96449 46351 96451 46389
rect 96451 46351 96503 46389
rect 96503 46351 96505 46389
rect 94927 46243 94929 46265
rect 94929 46243 94981 46265
rect 94981 46243 94983 46265
rect 94927 46231 94983 46243
rect 94927 46209 94929 46231
rect 94929 46209 94981 46231
rect 94981 46209 94983 46231
rect 96449 46325 96505 46327
rect 96449 46273 96451 46325
rect 96451 46273 96503 46325
rect 96503 46273 96505 46325
rect 96449 46271 96505 46273
rect 96449 46209 96451 46247
rect 96451 46209 96503 46247
rect 96503 46209 96505 46247
rect 96449 46191 96505 46209
rect 56127 45587 56183 45643
rect 63405 45587 63461 45643
rect 94922 45782 94924 45812
rect 94924 45782 94976 45812
rect 94976 45782 94978 45812
rect 94922 45770 94978 45782
rect 94922 45756 94924 45770
rect 94924 45756 94976 45770
rect 94976 45756 94978 45770
rect 94922 45718 94924 45732
rect 94924 45718 94976 45732
rect 94976 45718 94978 45732
rect 94922 45706 94978 45718
rect 94922 45676 94924 45706
rect 94924 45676 94976 45706
rect 94976 45676 94978 45706
rect 96450 45802 96452 45840
rect 96452 45802 96504 45840
rect 96504 45802 96506 45840
rect 96450 45790 96506 45802
rect 96450 45784 96452 45790
rect 96452 45784 96504 45790
rect 96504 45784 96506 45790
rect 96450 45738 96452 45760
rect 96452 45738 96504 45760
rect 96504 45738 96506 45760
rect 96450 45726 96506 45738
rect 96450 45704 96452 45726
rect 96452 45704 96504 45726
rect 96504 45704 96506 45726
rect 96450 45674 96452 45680
rect 96452 45674 96504 45680
rect 96504 45674 96506 45680
rect 96450 45662 96506 45674
rect 96450 45624 96452 45662
rect 96452 45624 96504 45662
rect 96504 45624 96506 45662
rect 92250 45601 92306 45603
rect 92250 45549 92252 45601
rect 92252 45549 92304 45601
rect 92304 45549 92306 45601
rect 92250 45547 92306 45549
rect 92575 45341 92631 45397
rect 99987 45171 100043 45173
rect 100067 45171 100123 45173
rect 100147 45171 100203 45173
rect 100227 45171 100283 45173
rect 100307 45171 100363 45173
rect 100387 45171 100443 45173
rect 100467 45171 100523 45173
rect 100547 45171 100603 45173
rect 100627 45171 100683 45173
rect 100707 45171 100763 45173
rect 100787 45171 100843 45173
rect 100867 45171 100923 45173
rect 100947 45171 101003 45173
rect 101027 45171 101083 45173
rect 101107 45171 101163 45173
rect 101187 45171 101243 45173
rect 101267 45171 101323 45173
rect 101347 45171 101403 45173
rect 101427 45171 101483 45173
rect 101507 45171 101563 45173
rect 101587 45171 101643 45173
rect 101667 45171 101723 45173
rect 101747 45171 101803 45173
rect 101827 45171 101883 45173
rect 101907 45171 101963 45173
rect 101987 45171 102043 45173
rect 102067 45171 102123 45173
rect 102147 45171 102203 45173
rect 102227 45171 102283 45173
rect 102307 45171 102363 45173
rect 102387 45171 102443 45173
rect 102467 45171 102523 45173
rect 102547 45171 102603 45173
rect 102627 45171 102683 45173
rect 102707 45171 102763 45173
rect 102787 45171 102843 45173
rect 102867 45171 102923 45173
rect 102947 45171 103003 45173
rect 103027 45171 103083 45173
rect 103107 45171 103163 45173
rect 103187 45171 103243 45173
rect 99987 45119 100009 45171
rect 100009 45119 100021 45171
rect 100021 45119 100043 45171
rect 100067 45119 100073 45171
rect 100073 45119 100085 45171
rect 100085 45119 100123 45171
rect 100147 45119 100149 45171
rect 100149 45119 100201 45171
rect 100201 45119 100203 45171
rect 100227 45119 100265 45171
rect 100265 45119 100277 45171
rect 100277 45119 100283 45171
rect 100307 45119 100329 45171
rect 100329 45119 100341 45171
rect 100341 45119 100363 45171
rect 100387 45119 100393 45171
rect 100393 45119 100405 45171
rect 100405 45119 100443 45171
rect 100467 45119 100469 45171
rect 100469 45119 100521 45171
rect 100521 45119 100523 45171
rect 100547 45119 100585 45171
rect 100585 45119 100597 45171
rect 100597 45119 100603 45171
rect 100627 45119 100649 45171
rect 100649 45119 100661 45171
rect 100661 45119 100683 45171
rect 100707 45119 100713 45171
rect 100713 45119 100725 45171
rect 100725 45119 100763 45171
rect 100787 45119 100789 45171
rect 100789 45119 100841 45171
rect 100841 45119 100843 45171
rect 100867 45119 100905 45171
rect 100905 45119 100917 45171
rect 100917 45119 100923 45171
rect 100947 45119 100969 45171
rect 100969 45119 100981 45171
rect 100981 45119 101003 45171
rect 101027 45119 101033 45171
rect 101033 45119 101045 45171
rect 101045 45119 101083 45171
rect 101107 45119 101109 45171
rect 101109 45119 101161 45171
rect 101161 45119 101163 45171
rect 101187 45119 101225 45171
rect 101225 45119 101237 45171
rect 101237 45119 101243 45171
rect 101267 45119 101289 45171
rect 101289 45119 101301 45171
rect 101301 45119 101323 45171
rect 101347 45119 101353 45171
rect 101353 45119 101365 45171
rect 101365 45119 101403 45171
rect 101427 45119 101429 45171
rect 101429 45119 101481 45171
rect 101481 45119 101483 45171
rect 101507 45119 101545 45171
rect 101545 45119 101557 45171
rect 101557 45119 101563 45171
rect 101587 45119 101609 45171
rect 101609 45119 101621 45171
rect 101621 45119 101643 45171
rect 101667 45119 101673 45171
rect 101673 45119 101685 45171
rect 101685 45119 101723 45171
rect 101747 45119 101749 45171
rect 101749 45119 101801 45171
rect 101801 45119 101803 45171
rect 101827 45119 101865 45171
rect 101865 45119 101877 45171
rect 101877 45119 101883 45171
rect 101907 45119 101929 45171
rect 101929 45119 101941 45171
rect 101941 45119 101963 45171
rect 101987 45119 101993 45171
rect 101993 45119 102005 45171
rect 102005 45119 102043 45171
rect 102067 45119 102069 45171
rect 102069 45119 102121 45171
rect 102121 45119 102123 45171
rect 102147 45119 102185 45171
rect 102185 45119 102197 45171
rect 102197 45119 102203 45171
rect 102227 45119 102249 45171
rect 102249 45119 102261 45171
rect 102261 45119 102283 45171
rect 102307 45119 102313 45171
rect 102313 45119 102325 45171
rect 102325 45119 102363 45171
rect 102387 45119 102389 45171
rect 102389 45119 102441 45171
rect 102441 45119 102443 45171
rect 102467 45119 102505 45171
rect 102505 45119 102517 45171
rect 102517 45119 102523 45171
rect 102547 45119 102569 45171
rect 102569 45119 102581 45171
rect 102581 45119 102603 45171
rect 102627 45119 102633 45171
rect 102633 45119 102645 45171
rect 102645 45119 102683 45171
rect 102707 45119 102709 45171
rect 102709 45119 102761 45171
rect 102761 45119 102763 45171
rect 102787 45119 102825 45171
rect 102825 45119 102837 45171
rect 102837 45119 102843 45171
rect 102867 45119 102889 45171
rect 102889 45119 102901 45171
rect 102901 45119 102923 45171
rect 102947 45119 102953 45171
rect 102953 45119 102965 45171
rect 102965 45119 103003 45171
rect 103027 45119 103029 45171
rect 103029 45119 103081 45171
rect 103081 45119 103083 45171
rect 103107 45119 103145 45171
rect 103145 45119 103157 45171
rect 103157 45119 103163 45171
rect 103187 45119 103209 45171
rect 103209 45119 103221 45171
rect 103221 45119 103243 45171
rect 99987 45117 100043 45119
rect 100067 45117 100123 45119
rect 100147 45117 100203 45119
rect 100227 45117 100283 45119
rect 100307 45117 100363 45119
rect 100387 45117 100443 45119
rect 100467 45117 100523 45119
rect 100547 45117 100603 45119
rect 100627 45117 100683 45119
rect 100707 45117 100763 45119
rect 100787 45117 100843 45119
rect 100867 45117 100923 45119
rect 100947 45117 101003 45119
rect 101027 45117 101083 45119
rect 101107 45117 101163 45119
rect 101187 45117 101243 45119
rect 101267 45117 101323 45119
rect 101347 45117 101403 45119
rect 101427 45117 101483 45119
rect 101507 45117 101563 45119
rect 101587 45117 101643 45119
rect 101667 45117 101723 45119
rect 101747 45117 101803 45119
rect 101827 45117 101883 45119
rect 101907 45117 101963 45119
rect 101987 45117 102043 45119
rect 102067 45117 102123 45119
rect 102147 45117 102203 45119
rect 102227 45117 102283 45119
rect 102307 45117 102363 45119
rect 102387 45117 102443 45119
rect 102467 45117 102523 45119
rect 102547 45117 102603 45119
rect 102627 45117 102683 45119
rect 102707 45117 102763 45119
rect 102787 45117 102843 45119
rect 102867 45117 102923 45119
rect 102947 45117 103003 45119
rect 103027 45117 103083 45119
rect 103107 45117 103163 45119
rect 103187 45117 103243 45119
rect 71786 45043 71842 45045
rect 71786 44991 71788 45043
rect 71788 44991 71840 45043
rect 71840 44991 71842 45043
rect 71786 44989 71842 44991
rect 63408 44919 63464 44975
rect 56127 44677 56183 44733
rect 42946 39332 43002 39388
rect 44034 38157 44090 38159
rect 44034 38105 44036 38157
rect 44036 38105 44088 38157
rect 44088 38105 44090 38157
rect 44034 38103 44090 38105
rect 57149 43475 57205 43531
rect 56342 43174 56398 43230
rect 71785 43289 71841 43345
rect 61971 43180 62267 43190
rect 60159 43122 60215 43124
rect 60159 43070 60161 43122
rect 60161 43070 60213 43122
rect 60213 43070 60215 43122
rect 60159 43068 60215 43070
rect 61971 43064 62267 43180
rect 61971 43054 62267 43064
rect 64183 43122 64239 43124
rect 64183 43070 64185 43122
rect 64185 43070 64237 43122
rect 64237 43070 64239 43122
rect 64183 43068 64239 43070
rect 66079 43122 66135 43124
rect 66079 43070 66081 43122
rect 66081 43070 66133 43122
rect 66133 43070 66135 43122
rect 66079 43068 66135 43070
rect 67330 43074 67386 43076
rect 67330 43022 67332 43074
rect 67332 43022 67384 43074
rect 67384 43022 67386 43074
rect 67330 43020 67386 43022
rect 80787 43398 80843 43400
rect 80787 43346 80789 43398
rect 80789 43346 80841 43398
rect 80841 43346 80843 43398
rect 80787 43344 80843 43346
rect 78069 43024 78125 43080
rect 62805 42872 62861 42928
rect 64804 42872 64860 42928
rect 61997 42613 62053 42669
rect 63995 42613 64051 42669
rect 65378 42734 65434 42736
rect 65378 42682 65380 42734
rect 65380 42682 65432 42734
rect 65432 42682 65434 42734
rect 65378 42680 65434 42682
rect 70672 42704 70728 42706
rect 70672 42652 70674 42704
rect 70674 42652 70726 42704
rect 70726 42652 70728 42704
rect 70672 42650 70728 42652
rect 60805 42274 60861 42330
rect 66804 42274 66860 42330
rect 59996 41993 60052 42049
rect 65997 41993 66053 42049
rect 57331 41788 57387 41790
rect 57331 41736 57333 41788
rect 57333 41736 57385 41788
rect 57385 41736 57387 41788
rect 57331 41734 57387 41736
rect 56277 41541 56333 41543
rect 56277 41489 56279 41541
rect 56279 41489 56331 41541
rect 56331 41489 56333 41541
rect 56277 41487 56333 41489
rect 71787 41504 71843 41560
rect 80787 41568 80843 41570
rect 80787 41516 80789 41568
rect 80789 41516 80841 41568
rect 80841 41516 80843 41568
rect 80787 41514 80843 41516
rect 61393 41305 61449 41307
rect 61393 41253 61395 41305
rect 61395 41253 61447 41305
rect 61447 41253 61449 41305
rect 61393 41251 61449 41253
rect 63325 41305 63381 41307
rect 63325 41253 63327 41305
rect 63327 41253 63379 41305
rect 63379 41253 63381 41305
rect 63325 41251 63381 41253
rect 46682 41119 46738 41175
rect 70701 41045 70757 41101
rect 46683 40250 46739 40306
rect 57361 40296 68217 40432
rect 51312 39724 51368 39726
rect 51312 39672 51314 39724
rect 51314 39672 51366 39724
rect 51366 39672 51368 39724
rect 51312 39670 51368 39672
rect 54090 39416 54146 39472
rect 52199 38401 52201 38431
rect 52201 38401 52253 38431
rect 52253 38401 52255 38431
rect 52199 38389 52255 38401
rect 52199 38375 52201 38389
rect 52201 38375 52253 38389
rect 52253 38375 52255 38389
rect 52199 38337 52201 38351
rect 52201 38337 52253 38351
rect 52253 38337 52255 38351
rect 52199 38325 52255 38337
rect 52199 38295 52201 38325
rect 52201 38295 52253 38325
rect 52253 38295 52255 38325
rect 52191 37944 52193 37982
rect 52193 37944 52245 37982
rect 52245 37944 52247 37982
rect 52191 37932 52247 37944
rect 52191 37926 52193 37932
rect 52193 37926 52245 37932
rect 52245 37926 52247 37932
rect 52191 37880 52193 37902
rect 52193 37880 52245 37902
rect 52245 37880 52247 37902
rect 52191 37868 52247 37880
rect 52191 37846 52193 37868
rect 52193 37846 52245 37868
rect 52245 37846 52247 37868
rect 52191 37816 52193 37822
rect 52193 37816 52245 37822
rect 52245 37816 52247 37822
rect 52191 37804 52247 37816
rect 52191 37766 52193 37804
rect 52193 37766 52245 37804
rect 52245 37766 52247 37804
rect 50936 34843 50992 34845
rect 51016 34843 51072 34845
rect 51096 34843 51152 34845
rect 50936 34791 50954 34843
rect 50954 34791 50992 34843
rect 51016 34791 51018 34843
rect 51018 34791 51070 34843
rect 51070 34791 51072 34843
rect 51096 34791 51134 34843
rect 51134 34791 51152 34843
rect 50936 34789 50992 34791
rect 51016 34789 51072 34791
rect 51096 34789 51152 34791
rect 46128 34185 46184 34241
rect 51392 34842 51448 34844
rect 51472 34842 51528 34844
rect 51552 34842 51608 34844
rect 51632 34842 51688 34844
rect 51392 34790 51418 34842
rect 51418 34790 51448 34842
rect 51472 34790 51482 34842
rect 51482 34790 51528 34842
rect 51552 34790 51598 34842
rect 51598 34790 51608 34842
rect 51632 34790 51662 34842
rect 51662 34790 51688 34842
rect 51392 34788 51448 34790
rect 51472 34788 51528 34790
rect 51552 34788 51608 34790
rect 51632 34788 51688 34790
rect 50942 34166 50998 34222
rect 50938 33600 50994 33602
rect 51018 33600 51074 33602
rect 51098 33600 51154 33602
rect 50938 33548 50956 33600
rect 50956 33548 50994 33600
rect 51018 33548 51020 33600
rect 51020 33548 51072 33600
rect 51072 33548 51074 33600
rect 51098 33548 51136 33600
rect 51136 33548 51154 33600
rect 50938 33546 50994 33548
rect 51018 33546 51074 33548
rect 51098 33546 51154 33548
rect 53963 38950 53965 38988
rect 53965 38950 54017 38988
rect 54017 38950 54019 38988
rect 53963 38938 54019 38950
rect 53963 38932 53965 38938
rect 53965 38932 54017 38938
rect 54017 38932 54019 38938
rect 53963 38886 53965 38908
rect 53965 38886 54017 38908
rect 54017 38886 54019 38908
rect 53963 38874 54019 38886
rect 53963 38852 53965 38874
rect 53965 38852 54017 38874
rect 54017 38852 54019 38874
rect 53963 38822 53965 38828
rect 53965 38822 54017 38828
rect 54017 38822 54019 38828
rect 53963 38810 54019 38822
rect 53963 38772 53965 38810
rect 53965 38772 54017 38810
rect 54017 38772 54019 38810
rect 54075 38606 54131 38662
rect 54500 37099 54556 37155
rect 55299 37137 55355 37139
rect 55299 37085 55301 37137
rect 55301 37085 55353 37137
rect 55353 37085 55355 37137
rect 55299 37083 55355 37085
rect 55299 37021 55301 37059
rect 55301 37021 55353 37059
rect 55353 37021 55355 37059
rect 55299 37009 55355 37021
rect 55299 37003 55301 37009
rect 55301 37003 55353 37009
rect 55353 37003 55355 37009
rect 55299 36957 55301 36979
rect 55301 36957 55353 36979
rect 55353 36957 55355 36979
rect 55299 36945 55355 36957
rect 55299 36923 55301 36945
rect 55301 36923 55353 36945
rect 55353 36923 55355 36945
rect 55299 36893 55301 36899
rect 55301 36893 55353 36899
rect 55353 36893 55355 36899
rect 55299 36881 55355 36893
rect 55299 36843 55301 36881
rect 55301 36843 55353 36881
rect 55353 36843 55355 36881
rect 55299 36817 55355 36819
rect 55299 36765 55301 36817
rect 55301 36765 55353 36817
rect 55353 36765 55355 36817
rect 55299 36763 55355 36765
rect 51737 34166 51793 34222
rect 52309 34195 52365 34251
rect 52650 34195 52706 34251
rect 51392 33600 51448 33602
rect 51472 33600 51528 33602
rect 51552 33600 51608 33602
rect 51632 33600 51688 33602
rect 51392 33548 51438 33600
rect 51438 33548 51448 33600
rect 51472 33548 51502 33600
rect 51502 33548 51514 33600
rect 51514 33548 51528 33600
rect 51552 33548 51566 33600
rect 51566 33548 51578 33600
rect 51578 33548 51608 33600
rect 51632 33548 51642 33600
rect 51642 33548 51688 33600
rect 51392 33546 51448 33548
rect 51472 33546 51528 33548
rect 51552 33546 51608 33548
rect 51632 33546 51688 33548
rect 40349 31569 40405 31625
rect 49883 31235 50339 31253
rect 49883 31055 49893 31235
rect 49893 31055 50329 31235
rect 50329 31055 50339 31235
rect 49883 31037 50339 31055
rect 31582 30630 31584 30668
rect 31584 30630 31636 30668
rect 31636 30630 31638 30668
rect 31582 30618 31638 30630
rect 31582 30612 31584 30618
rect 31584 30612 31636 30618
rect 31636 30612 31638 30618
rect 31582 30566 31584 30588
rect 31584 30566 31636 30588
rect 31636 30566 31638 30588
rect 31582 30554 31638 30566
rect 31582 30532 31584 30554
rect 31584 30532 31636 30554
rect 31636 30532 31638 30554
rect 31582 30502 31584 30508
rect 31584 30502 31636 30508
rect 31636 30502 31638 30508
rect 31582 30490 31638 30502
rect 31582 30452 31584 30490
rect 31584 30452 31636 30490
rect 31636 30452 31638 30490
rect 38847 30319 38903 30321
rect 38847 30267 38849 30319
rect 38849 30267 38901 30319
rect 38901 30267 38903 30319
rect 38847 30265 38903 30267
rect 44023 30329 44079 30331
rect 44023 30277 44025 30329
rect 44025 30277 44077 30329
rect 44077 30277 44079 30329
rect 44023 30275 44079 30277
rect 52189 30687 52245 30713
rect 52189 30657 52191 30687
rect 52191 30657 52243 30687
rect 52243 30657 52245 30687
rect 52189 30623 52245 30633
rect 52189 30577 52191 30623
rect 52191 30577 52243 30623
rect 52243 30577 52245 30623
rect 52189 30507 52191 30553
rect 52191 30507 52243 30553
rect 52243 30507 52245 30553
rect 52189 30497 52245 30507
rect 52189 30443 52191 30473
rect 52191 30443 52243 30473
rect 52243 30443 52245 30473
rect 52189 30417 52245 30443
rect 31581 30143 31583 30181
rect 31583 30143 31635 30181
rect 31635 30143 31637 30181
rect 31581 30131 31637 30143
rect 31581 30125 31583 30131
rect 31583 30125 31635 30131
rect 31635 30125 31637 30131
rect 31581 30079 31583 30101
rect 31583 30079 31635 30101
rect 31635 30079 31637 30101
rect 31581 30067 31637 30079
rect 31581 30045 31583 30067
rect 31583 30045 31635 30067
rect 31635 30045 31637 30067
rect 31581 30015 31583 30021
rect 31583 30015 31635 30021
rect 31635 30015 31637 30021
rect 31581 30003 31637 30015
rect 31581 29965 31583 30003
rect 31583 29965 31635 30003
rect 31635 29965 31637 30003
rect 52192 30116 52194 30146
rect 52194 30116 52246 30146
rect 52246 30116 52248 30146
rect 52192 30104 52248 30116
rect 52192 30090 52194 30104
rect 52194 30090 52246 30104
rect 52246 30090 52248 30104
rect 52192 30052 52194 30066
rect 52194 30052 52246 30066
rect 52246 30052 52248 30066
rect 52192 30040 52248 30052
rect 52192 30010 52194 30040
rect 52194 30010 52246 30040
rect 52246 30010 52248 30040
rect 55600 36425 55656 36427
rect 55600 36373 55602 36425
rect 55602 36373 55654 36425
rect 55654 36373 55656 36425
rect 55600 36371 55656 36373
rect 54213 36290 54269 36346
rect 55172 35497 55228 35553
rect 55340 35542 55396 35544
rect 55340 35490 55342 35542
rect 55342 35490 55394 35542
rect 55394 35490 55396 35542
rect 55340 35488 55396 35490
rect 55340 35426 55342 35464
rect 55342 35426 55394 35464
rect 55394 35426 55396 35464
rect 55340 35414 55396 35426
rect 55340 35408 55342 35414
rect 55342 35408 55394 35414
rect 55394 35408 55396 35414
rect 55340 35362 55342 35384
rect 55342 35362 55394 35384
rect 55394 35362 55396 35384
rect 55340 35350 55396 35362
rect 55340 35328 55342 35350
rect 55342 35328 55394 35350
rect 55394 35328 55396 35350
rect 55340 35298 55342 35304
rect 55342 35298 55394 35304
rect 55394 35298 55396 35304
rect 55340 35286 55396 35298
rect 55340 35248 55342 35286
rect 55342 35248 55394 35286
rect 55394 35248 55396 35286
rect 55340 35222 55396 35224
rect 55340 35170 55342 35222
rect 55342 35170 55394 35222
rect 55394 35170 55396 35222
rect 55340 35168 55396 35170
rect 54886 34691 54942 34747
rect 55600 34799 55656 34801
rect 55600 34747 55602 34799
rect 55602 34747 55654 34799
rect 55654 34747 55656 34799
rect 55600 34745 55656 34747
rect 55172 33899 55228 33955
rect 55339 33939 55395 33941
rect 55339 33887 55341 33939
rect 55341 33887 55393 33939
rect 55393 33887 55395 33939
rect 55339 33885 55395 33887
rect 55339 33823 55341 33861
rect 55341 33823 55393 33861
rect 55393 33823 55395 33861
rect 55339 33811 55395 33823
rect 55339 33805 55341 33811
rect 55341 33805 55393 33811
rect 55393 33805 55395 33811
rect 55339 33759 55341 33781
rect 55341 33759 55393 33781
rect 55393 33759 55395 33781
rect 55339 33747 55395 33759
rect 55339 33725 55341 33747
rect 55341 33725 55393 33747
rect 55393 33725 55395 33747
rect 55339 33695 55341 33701
rect 55341 33695 55393 33701
rect 55393 33695 55395 33701
rect 55339 33683 55395 33695
rect 55339 33645 55341 33683
rect 55341 33645 55393 33683
rect 55393 33645 55395 33683
rect 55339 33619 55395 33621
rect 55339 33567 55341 33619
rect 55341 33567 55393 33619
rect 55393 33567 55395 33619
rect 55339 33565 55395 33567
rect 54886 33091 54942 33147
rect 55600 33141 55656 33143
rect 55600 33089 55602 33141
rect 55602 33089 55654 33141
rect 55654 33089 55656 33141
rect 55600 33087 55656 33089
rect 54500 32297 54556 32353
rect 55342 32338 55398 32340
rect 55342 32286 55344 32338
rect 55344 32286 55396 32338
rect 55396 32286 55398 32338
rect 55342 32284 55398 32286
rect 55342 32222 55344 32260
rect 55344 32222 55396 32260
rect 55396 32222 55398 32260
rect 55342 32210 55398 32222
rect 55342 32204 55344 32210
rect 55344 32204 55396 32210
rect 55396 32204 55398 32210
rect 55342 32158 55344 32180
rect 55344 32158 55396 32180
rect 55396 32158 55398 32180
rect 55342 32146 55398 32158
rect 55342 32124 55344 32146
rect 55344 32124 55396 32146
rect 55396 32124 55398 32146
rect 55342 32094 55344 32100
rect 55344 32094 55396 32100
rect 55396 32094 55398 32100
rect 55342 32082 55398 32094
rect 55342 32044 55344 32082
rect 55344 32044 55396 32082
rect 55396 32044 55398 32082
rect 55342 32018 55398 32020
rect 55342 31966 55344 32018
rect 55344 31966 55396 32018
rect 55396 31966 55398 32018
rect 55342 31964 55398 31966
rect 54213 31489 54269 31545
rect 55600 31602 55656 31604
rect 55600 31550 55602 31602
rect 55602 31550 55654 31602
rect 55654 31550 55656 31602
rect 55600 31548 55656 31550
rect 55600 31208 55602 31246
rect 55602 31208 55654 31246
rect 55654 31208 55656 31246
rect 55600 31196 55656 31208
rect 55600 31190 55602 31196
rect 55602 31190 55654 31196
rect 55654 31190 55656 31196
rect 55600 31144 55602 31166
rect 55602 31144 55654 31166
rect 55654 31144 55656 31166
rect 55600 31132 55656 31144
rect 55600 31110 55602 31132
rect 55602 31110 55654 31132
rect 55654 31110 55656 31132
rect 55600 31080 55602 31086
rect 55602 31080 55654 31086
rect 55654 31080 55656 31086
rect 55600 31068 55656 31080
rect 55600 31030 55602 31068
rect 55602 31030 55654 31068
rect 55654 31030 55656 31068
rect 55600 30467 55656 30469
rect 55600 30415 55602 30467
rect 55602 30415 55654 30467
rect 55654 30415 55656 30467
rect 55600 30413 55656 30415
rect 54048 30004 54104 30060
rect 53914 29528 53916 29566
rect 53916 29528 53968 29566
rect 53968 29528 53970 29566
rect 53914 29516 53970 29528
rect 53914 29510 53916 29516
rect 53916 29510 53968 29516
rect 53968 29510 53970 29516
rect 53914 29464 53916 29486
rect 53916 29464 53968 29486
rect 53968 29464 53970 29486
rect 53914 29452 53970 29464
rect 53914 29430 53916 29452
rect 53916 29430 53968 29452
rect 53968 29430 53970 29452
rect 53914 29400 53916 29406
rect 53916 29400 53968 29406
rect 53968 29400 53970 29406
rect 53914 29388 53970 29400
rect 53914 29350 53916 29388
rect 53916 29350 53968 29388
rect 53968 29350 53970 29388
rect 54070 29195 54126 29251
rect 46332 29009 46388 29065
rect 57133 40182 57269 40184
rect 57133 34690 57143 40182
rect 57143 34690 57259 40182
rect 57259 34690 57269 40182
rect 57133 34688 57269 34690
rect 68345 40185 68481 40195
rect 68345 38469 68355 40185
rect 68355 38469 68471 40185
rect 68471 38469 68481 40185
rect 68345 38459 68481 38469
rect 80784 39804 80840 39806
rect 80784 39752 80786 39804
rect 80786 39752 80838 39804
rect 80838 39752 80840 39804
rect 80784 39750 80840 39752
rect 71784 39673 71840 39729
rect 78026 39512 78082 39514
rect 78026 39460 78028 39512
rect 78028 39460 78080 39512
rect 78080 39460 78082 39512
rect 78026 39458 78082 39460
rect 71788 39244 71844 39246
rect 71788 39192 71790 39244
rect 71790 39192 71842 39244
rect 71842 39192 71844 39244
rect 71788 39190 71844 39192
rect 68386 37906 68442 37962
rect 68386 37826 68442 37882
rect 68386 37746 68442 37802
rect 68386 37666 68442 37722
rect 68386 37586 68442 37642
rect 68386 37506 68442 37562
rect 68386 37426 68442 37482
rect 68386 37346 68442 37402
rect 68386 37266 68442 37322
rect 68386 37186 68442 37242
rect 68386 37106 68442 37162
rect 68386 37026 68442 37082
rect 71783 37981 71839 37983
rect 71783 37929 71785 37981
rect 71785 37929 71837 37981
rect 71837 37929 71839 37981
rect 71783 37927 71839 37929
rect 80784 38013 80840 38015
rect 80784 37961 80786 38013
rect 80786 37961 80838 38013
rect 80838 37961 80840 38013
rect 80784 37959 80840 37961
rect 70734 37490 70790 37546
rect 68346 36122 68482 36132
rect 68346 35366 68356 36122
rect 68356 35366 68472 36122
rect 68472 35366 68482 36122
rect 68346 35356 68482 35366
rect 71800 36196 71856 36198
rect 71800 36144 71802 36196
rect 71802 36144 71854 36196
rect 71854 36144 71856 36196
rect 71800 36142 71856 36144
rect 80789 36206 80845 36208
rect 80789 36154 80791 36206
rect 80791 36154 80843 36206
rect 80843 36154 80845 36206
rect 80789 36152 80845 36154
rect 78083 35868 78139 35924
rect 70797 35638 70853 35694
rect 63596 34400 68292 34536
rect 71789 34399 71845 34401
rect 71789 34347 71791 34399
rect 71791 34347 71843 34399
rect 71843 34347 71845 34399
rect 71789 34345 71845 34347
rect 80789 34396 80845 34398
rect 80789 34344 80791 34396
rect 80791 34344 80843 34396
rect 80843 34344 80845 34396
rect 80789 34342 80845 34344
rect 92587 32493 92643 32549
rect 93164 33116 93220 33172
rect 93729 32431 93785 32487
rect 92122 32299 92178 32301
rect 92122 32247 92124 32299
rect 92124 32247 92176 32299
rect 92176 32247 92178 32299
rect 92122 32245 92178 32247
rect 95676 32045 95732 32055
rect 95676 31999 95678 32045
rect 95678 31999 95730 32045
rect 95730 31999 95732 32045
rect 95676 31929 95678 31975
rect 95678 31929 95730 31975
rect 95730 31929 95732 31975
rect 95676 31919 95732 31929
rect 97206 32087 97208 32117
rect 97208 32087 97260 32117
rect 97260 32087 97262 32117
rect 97206 32075 97262 32087
rect 97206 32061 97208 32075
rect 97208 32061 97260 32075
rect 97260 32061 97262 32075
rect 97206 32023 97208 32037
rect 97208 32023 97260 32037
rect 97260 32023 97262 32037
rect 97206 32011 97262 32023
rect 97206 31981 97208 32011
rect 97208 31981 97260 32011
rect 97260 31981 97262 32011
rect 93402 31895 93458 31897
rect 93482 31895 93538 31897
rect 93562 31895 93618 31897
rect 93402 31843 93420 31895
rect 93420 31843 93458 31895
rect 93482 31843 93484 31895
rect 93484 31843 93536 31895
rect 93536 31843 93538 31895
rect 93562 31843 93600 31895
rect 93600 31843 93618 31895
rect 93402 31841 93458 31843
rect 93482 31841 93538 31843
rect 93562 31841 93618 31843
rect 95674 31529 95676 31559
rect 95676 31529 95728 31559
rect 95728 31529 95730 31559
rect 95674 31517 95730 31529
rect 95674 31503 95676 31517
rect 95676 31503 95728 31517
rect 95728 31503 95730 31517
rect 95674 31465 95676 31479
rect 95676 31465 95728 31479
rect 95728 31465 95730 31479
rect 95674 31453 95730 31465
rect 95674 31423 95676 31453
rect 95676 31423 95728 31453
rect 95728 31423 95730 31453
rect 97193 31542 97195 31572
rect 97195 31542 97247 31572
rect 97247 31542 97249 31572
rect 97193 31530 97249 31542
rect 97193 31516 97195 31530
rect 97195 31516 97247 31530
rect 97247 31516 97249 31530
rect 97193 31478 97195 31492
rect 97195 31478 97247 31492
rect 97247 31478 97249 31492
rect 97193 31466 97249 31478
rect 97193 31436 97195 31466
rect 97195 31436 97247 31466
rect 97247 31436 97249 31466
rect 93472 31354 93528 31356
rect 93552 31354 93608 31356
rect 93472 31302 93482 31354
rect 93482 31302 93528 31354
rect 93552 31302 93598 31354
rect 93598 31302 93608 31354
rect 93472 31300 93528 31302
rect 93552 31300 93608 31302
rect 92126 31239 92182 31241
rect 92126 31187 92128 31239
rect 92128 31187 92180 31239
rect 92180 31187 92182 31239
rect 92126 31185 92182 31187
rect 99728 31235 99784 31237
rect 99808 31235 99864 31237
rect 99888 31235 99944 31237
rect 99968 31235 100024 31237
rect 100048 31235 100104 31237
rect 100128 31235 100184 31237
rect 100208 31235 100264 31237
rect 100288 31235 100344 31237
rect 100368 31235 100424 31237
rect 100448 31235 100504 31237
rect 100528 31235 100584 31237
rect 100608 31235 100664 31237
rect 100688 31235 100744 31237
rect 100768 31235 100824 31237
rect 100848 31235 100904 31237
rect 100928 31235 100984 31237
rect 101008 31235 101064 31237
rect 101088 31235 101144 31237
rect 101168 31235 101224 31237
rect 101248 31235 101304 31237
rect 101328 31235 101384 31237
rect 101408 31235 101464 31237
rect 101488 31235 101544 31237
rect 101568 31235 101624 31237
rect 101648 31235 101704 31237
rect 101728 31235 101784 31237
rect 101808 31235 101864 31237
rect 101888 31235 101944 31237
rect 101968 31235 102024 31237
rect 102048 31235 102104 31237
rect 102128 31235 102184 31237
rect 102208 31235 102264 31237
rect 102288 31235 102344 31237
rect 102368 31235 102424 31237
rect 102448 31235 102504 31237
rect 102528 31235 102584 31237
rect 102608 31235 102664 31237
rect 102688 31235 102744 31237
rect 102768 31235 102824 31237
rect 102848 31235 102904 31237
rect 102928 31235 102984 31237
rect 99728 31183 99750 31235
rect 99750 31183 99762 31235
rect 99762 31183 99784 31235
rect 99808 31183 99814 31235
rect 99814 31183 99826 31235
rect 99826 31183 99864 31235
rect 99888 31183 99890 31235
rect 99890 31183 99942 31235
rect 99942 31183 99944 31235
rect 99968 31183 100006 31235
rect 100006 31183 100018 31235
rect 100018 31183 100024 31235
rect 100048 31183 100070 31235
rect 100070 31183 100082 31235
rect 100082 31183 100104 31235
rect 100128 31183 100134 31235
rect 100134 31183 100146 31235
rect 100146 31183 100184 31235
rect 100208 31183 100210 31235
rect 100210 31183 100262 31235
rect 100262 31183 100264 31235
rect 100288 31183 100326 31235
rect 100326 31183 100338 31235
rect 100338 31183 100344 31235
rect 100368 31183 100390 31235
rect 100390 31183 100402 31235
rect 100402 31183 100424 31235
rect 100448 31183 100454 31235
rect 100454 31183 100466 31235
rect 100466 31183 100504 31235
rect 100528 31183 100530 31235
rect 100530 31183 100582 31235
rect 100582 31183 100584 31235
rect 100608 31183 100646 31235
rect 100646 31183 100658 31235
rect 100658 31183 100664 31235
rect 100688 31183 100710 31235
rect 100710 31183 100722 31235
rect 100722 31183 100744 31235
rect 100768 31183 100774 31235
rect 100774 31183 100786 31235
rect 100786 31183 100824 31235
rect 100848 31183 100850 31235
rect 100850 31183 100902 31235
rect 100902 31183 100904 31235
rect 100928 31183 100966 31235
rect 100966 31183 100978 31235
rect 100978 31183 100984 31235
rect 101008 31183 101030 31235
rect 101030 31183 101042 31235
rect 101042 31183 101064 31235
rect 101088 31183 101094 31235
rect 101094 31183 101106 31235
rect 101106 31183 101144 31235
rect 101168 31183 101170 31235
rect 101170 31183 101222 31235
rect 101222 31183 101224 31235
rect 101248 31183 101286 31235
rect 101286 31183 101298 31235
rect 101298 31183 101304 31235
rect 101328 31183 101350 31235
rect 101350 31183 101362 31235
rect 101362 31183 101384 31235
rect 101408 31183 101414 31235
rect 101414 31183 101426 31235
rect 101426 31183 101464 31235
rect 101488 31183 101490 31235
rect 101490 31183 101542 31235
rect 101542 31183 101544 31235
rect 101568 31183 101606 31235
rect 101606 31183 101618 31235
rect 101618 31183 101624 31235
rect 101648 31183 101670 31235
rect 101670 31183 101682 31235
rect 101682 31183 101704 31235
rect 101728 31183 101734 31235
rect 101734 31183 101746 31235
rect 101746 31183 101784 31235
rect 101808 31183 101810 31235
rect 101810 31183 101862 31235
rect 101862 31183 101864 31235
rect 101888 31183 101926 31235
rect 101926 31183 101938 31235
rect 101938 31183 101944 31235
rect 101968 31183 101990 31235
rect 101990 31183 102002 31235
rect 102002 31183 102024 31235
rect 102048 31183 102054 31235
rect 102054 31183 102066 31235
rect 102066 31183 102104 31235
rect 102128 31183 102130 31235
rect 102130 31183 102182 31235
rect 102182 31183 102184 31235
rect 102208 31183 102246 31235
rect 102246 31183 102258 31235
rect 102258 31183 102264 31235
rect 102288 31183 102310 31235
rect 102310 31183 102322 31235
rect 102322 31183 102344 31235
rect 102368 31183 102374 31235
rect 102374 31183 102386 31235
rect 102386 31183 102424 31235
rect 102448 31183 102450 31235
rect 102450 31183 102502 31235
rect 102502 31183 102504 31235
rect 102528 31183 102566 31235
rect 102566 31183 102578 31235
rect 102578 31183 102584 31235
rect 102608 31183 102630 31235
rect 102630 31183 102642 31235
rect 102642 31183 102664 31235
rect 102688 31183 102694 31235
rect 102694 31183 102706 31235
rect 102706 31183 102744 31235
rect 102768 31183 102770 31235
rect 102770 31183 102822 31235
rect 102822 31183 102824 31235
rect 102848 31183 102886 31235
rect 102886 31183 102898 31235
rect 102898 31183 102904 31235
rect 102928 31183 102950 31235
rect 102950 31183 102962 31235
rect 102962 31183 102984 31235
rect 99728 31181 99784 31183
rect 99808 31181 99864 31183
rect 99888 31181 99944 31183
rect 99968 31181 100024 31183
rect 100048 31181 100104 31183
rect 100128 31181 100184 31183
rect 100208 31181 100264 31183
rect 100288 31181 100344 31183
rect 100368 31181 100424 31183
rect 100448 31181 100504 31183
rect 100528 31181 100584 31183
rect 100608 31181 100664 31183
rect 100688 31181 100744 31183
rect 100768 31181 100824 31183
rect 100848 31181 100904 31183
rect 100928 31181 100984 31183
rect 101008 31181 101064 31183
rect 101088 31181 101144 31183
rect 101168 31181 101224 31183
rect 101248 31181 101304 31183
rect 101328 31181 101384 31183
rect 101408 31181 101464 31183
rect 101488 31181 101544 31183
rect 101568 31181 101624 31183
rect 101648 31181 101704 31183
rect 101728 31181 101784 31183
rect 101808 31181 101864 31183
rect 101888 31181 101944 31183
rect 101968 31181 102024 31183
rect 102048 31181 102104 31183
rect 102128 31181 102184 31183
rect 102208 31181 102264 31183
rect 102288 31181 102344 31183
rect 102368 31181 102424 31183
rect 102448 31181 102504 31183
rect 102528 31181 102584 31183
rect 102608 31181 102664 31183
rect 102688 31181 102744 31183
rect 102768 31181 102824 31183
rect 102848 31181 102904 31183
rect 102928 31181 102984 31183
rect 92125 30970 92181 30972
rect 92125 30918 92127 30970
rect 92127 30918 92179 30970
rect 92179 30918 92181 30970
rect 92125 30916 92181 30918
rect 93460 30806 93516 30808
rect 93460 30754 93462 30806
rect 93462 30754 93514 30806
rect 93514 30754 93516 30806
rect 93460 30752 93516 30754
rect 95676 30672 95678 30694
rect 95678 30672 95730 30694
rect 95730 30672 95732 30694
rect 95676 30660 95732 30672
rect 95676 30638 95678 30660
rect 95678 30638 95730 30660
rect 95730 30638 95732 30660
rect 97198 30751 97200 30781
rect 97200 30751 97252 30781
rect 97252 30751 97254 30781
rect 97198 30739 97254 30751
rect 97198 30725 97200 30739
rect 97200 30725 97252 30739
rect 97252 30725 97254 30739
rect 97198 30687 97200 30701
rect 97200 30687 97252 30701
rect 97252 30687 97254 30701
rect 97198 30675 97254 30687
rect 97198 30645 97200 30675
rect 97200 30645 97252 30675
rect 97252 30645 97254 30675
rect 94085 30265 94141 30267
rect 94085 30213 94087 30265
rect 94087 30213 94139 30265
rect 94139 30213 94141 30265
rect 94085 30211 94141 30213
rect 95669 30198 95671 30228
rect 95671 30198 95723 30228
rect 95723 30198 95725 30228
rect 95669 30186 95725 30198
rect 95669 30172 95671 30186
rect 95671 30172 95723 30186
rect 95723 30172 95725 30186
rect 95669 30134 95671 30148
rect 95671 30134 95723 30148
rect 95723 30134 95725 30148
rect 95669 30122 95725 30134
rect 95669 30092 95671 30122
rect 95671 30092 95723 30122
rect 95723 30092 95725 30122
rect 97198 30195 97200 30225
rect 97200 30195 97252 30225
rect 97252 30195 97254 30225
rect 97198 30183 97254 30195
rect 97198 30169 97200 30183
rect 97200 30169 97252 30183
rect 97252 30169 97254 30183
rect 97198 30131 97200 30145
rect 97200 30131 97252 30145
rect 97252 30131 97254 30145
rect 97198 30119 97254 30131
rect 97198 30089 97200 30119
rect 97200 30089 97252 30119
rect 97252 30089 97254 30119
rect 92125 29901 92181 29903
rect 92125 29849 92127 29901
rect 92127 29849 92179 29901
rect 92179 29849 92181 29901
rect 92125 29847 92181 29849
rect 93085 29723 93141 29725
rect 93165 29723 93221 29725
rect 93085 29671 93095 29723
rect 93095 29671 93141 29723
rect 93165 29671 93211 29723
rect 93211 29671 93221 29723
rect 93085 29669 93141 29671
rect 93165 29669 93221 29671
rect 104577 29794 104793 29812
rect 104577 29614 104595 29794
rect 104595 29614 104775 29794
rect 104775 29614 104793 29794
rect 104577 29596 104793 29614
rect 92122 29578 92178 29580
rect 92122 29526 92124 29578
rect 92124 29526 92176 29578
rect 92176 29526 92178 29578
rect 92122 29524 92178 29526
rect 95677 29282 95679 29304
rect 95679 29282 95731 29304
rect 95731 29282 95733 29304
rect 95677 29270 95733 29282
rect 95677 29248 95679 29270
rect 95679 29248 95731 29270
rect 95731 29248 95733 29270
rect 97215 29371 97217 29401
rect 97217 29371 97269 29401
rect 97269 29371 97271 29401
rect 97215 29359 97271 29371
rect 97215 29345 97217 29359
rect 97217 29345 97269 29359
rect 97269 29345 97271 29359
rect 97215 29307 97217 29321
rect 97217 29307 97269 29321
rect 97269 29307 97271 29321
rect 97215 29295 97271 29307
rect 97215 29265 97217 29295
rect 97217 29265 97269 29295
rect 97269 29265 97271 29295
rect 93610 29175 93666 29177
rect 93690 29175 93746 29177
rect 93770 29175 93826 29177
rect 93610 29123 93628 29175
rect 93628 29123 93666 29175
rect 93690 29123 93692 29175
rect 93692 29123 93744 29175
rect 93744 29123 93746 29175
rect 93770 29123 93808 29175
rect 93808 29123 93826 29175
rect 93610 29121 93666 29123
rect 93690 29121 93746 29123
rect 93770 29121 93826 29123
rect 95668 28845 95670 28875
rect 95670 28845 95722 28875
rect 95722 28845 95724 28875
rect 95668 28833 95724 28845
rect 95668 28819 95670 28833
rect 95670 28819 95722 28833
rect 95722 28819 95724 28833
rect 95668 28781 95670 28795
rect 95670 28781 95722 28795
rect 95722 28781 95724 28795
rect 95668 28769 95724 28781
rect 95668 28739 95670 28769
rect 95670 28739 95722 28769
rect 95722 28739 95724 28769
rect 97198 28823 97200 28853
rect 97200 28823 97252 28853
rect 97252 28823 97254 28853
rect 97198 28811 97254 28823
rect 97198 28797 97200 28811
rect 97200 28797 97252 28811
rect 97252 28797 97254 28811
rect 97198 28759 97200 28773
rect 97200 28759 97252 28773
rect 97252 28759 97254 28773
rect 97198 28747 97254 28759
rect 97198 28717 97200 28747
rect 97200 28717 97252 28747
rect 97252 28717 97254 28747
rect 93462 28632 93518 28634
rect 93542 28632 93598 28634
rect 93462 28580 93472 28632
rect 93472 28580 93518 28632
rect 93542 28580 93588 28632
rect 93588 28580 93598 28632
rect 93462 28578 93518 28580
rect 93542 28578 93598 28580
rect 92133 28508 92189 28510
rect 92133 28456 92135 28508
rect 92135 28456 92187 28508
rect 92187 28456 92189 28508
rect 92133 28454 92189 28456
rect 92122 28203 92178 28205
rect 92122 28151 92124 28203
rect 92124 28151 92176 28203
rect 92176 28151 92178 28203
rect 92122 28149 92178 28151
rect 99705 28236 99761 28238
rect 99785 28236 99841 28238
rect 99865 28236 99921 28238
rect 99945 28236 100001 28238
rect 100025 28236 100081 28238
rect 100105 28236 100161 28238
rect 100185 28236 100241 28238
rect 100265 28236 100321 28238
rect 100345 28236 100401 28238
rect 100425 28236 100481 28238
rect 100505 28236 100561 28238
rect 100585 28236 100641 28238
rect 100665 28236 100721 28238
rect 100745 28236 100801 28238
rect 100825 28236 100881 28238
rect 100905 28236 100961 28238
rect 100985 28236 101041 28238
rect 101065 28236 101121 28238
rect 101145 28236 101201 28238
rect 101225 28236 101281 28238
rect 101305 28236 101361 28238
rect 101385 28236 101441 28238
rect 101465 28236 101521 28238
rect 101545 28236 101601 28238
rect 101625 28236 101681 28238
rect 101705 28236 101761 28238
rect 101785 28236 101841 28238
rect 101865 28236 101921 28238
rect 101945 28236 102001 28238
rect 102025 28236 102081 28238
rect 102105 28236 102161 28238
rect 102185 28236 102241 28238
rect 102265 28236 102321 28238
rect 102345 28236 102401 28238
rect 102425 28236 102481 28238
rect 102505 28236 102561 28238
rect 102585 28236 102641 28238
rect 102665 28236 102721 28238
rect 102745 28236 102801 28238
rect 102825 28236 102881 28238
rect 102905 28236 102961 28238
rect 102985 28236 103041 28238
rect 99705 28184 99715 28236
rect 99715 28184 99761 28236
rect 99785 28184 99831 28236
rect 99831 28184 99841 28236
rect 99865 28184 99895 28236
rect 99895 28184 99907 28236
rect 99907 28184 99921 28236
rect 99945 28184 99959 28236
rect 99959 28184 99971 28236
rect 99971 28184 100001 28236
rect 100025 28184 100035 28236
rect 100035 28184 100081 28236
rect 100105 28184 100151 28236
rect 100151 28184 100161 28236
rect 100185 28184 100215 28236
rect 100215 28184 100227 28236
rect 100227 28184 100241 28236
rect 100265 28184 100279 28236
rect 100279 28184 100291 28236
rect 100291 28184 100321 28236
rect 100345 28184 100355 28236
rect 100355 28184 100401 28236
rect 100425 28184 100471 28236
rect 100471 28184 100481 28236
rect 100505 28184 100535 28236
rect 100535 28184 100547 28236
rect 100547 28184 100561 28236
rect 100585 28184 100599 28236
rect 100599 28184 100611 28236
rect 100611 28184 100641 28236
rect 100665 28184 100675 28236
rect 100675 28184 100721 28236
rect 100745 28184 100791 28236
rect 100791 28184 100801 28236
rect 100825 28184 100855 28236
rect 100855 28184 100867 28236
rect 100867 28184 100881 28236
rect 100905 28184 100919 28236
rect 100919 28184 100931 28236
rect 100931 28184 100961 28236
rect 100985 28184 100995 28236
rect 100995 28184 101041 28236
rect 101065 28184 101111 28236
rect 101111 28184 101121 28236
rect 101145 28184 101175 28236
rect 101175 28184 101187 28236
rect 101187 28184 101201 28236
rect 101225 28184 101239 28236
rect 101239 28184 101251 28236
rect 101251 28184 101281 28236
rect 101305 28184 101315 28236
rect 101315 28184 101361 28236
rect 101385 28184 101431 28236
rect 101431 28184 101441 28236
rect 101465 28184 101495 28236
rect 101495 28184 101507 28236
rect 101507 28184 101521 28236
rect 101545 28184 101559 28236
rect 101559 28184 101571 28236
rect 101571 28184 101601 28236
rect 101625 28184 101635 28236
rect 101635 28184 101681 28236
rect 101705 28184 101751 28236
rect 101751 28184 101761 28236
rect 101785 28184 101815 28236
rect 101815 28184 101827 28236
rect 101827 28184 101841 28236
rect 101865 28184 101879 28236
rect 101879 28184 101891 28236
rect 101891 28184 101921 28236
rect 101945 28184 101955 28236
rect 101955 28184 102001 28236
rect 102025 28184 102071 28236
rect 102071 28184 102081 28236
rect 102105 28184 102135 28236
rect 102135 28184 102147 28236
rect 102147 28184 102161 28236
rect 102185 28184 102199 28236
rect 102199 28184 102211 28236
rect 102211 28184 102241 28236
rect 102265 28184 102275 28236
rect 102275 28184 102321 28236
rect 102345 28184 102391 28236
rect 102391 28184 102401 28236
rect 102425 28184 102455 28236
rect 102455 28184 102467 28236
rect 102467 28184 102481 28236
rect 102505 28184 102519 28236
rect 102519 28184 102531 28236
rect 102531 28184 102561 28236
rect 102585 28184 102595 28236
rect 102595 28184 102641 28236
rect 102665 28184 102711 28236
rect 102711 28184 102721 28236
rect 102745 28184 102775 28236
rect 102775 28184 102787 28236
rect 102787 28184 102801 28236
rect 102825 28184 102839 28236
rect 102839 28184 102851 28236
rect 102851 28184 102881 28236
rect 102905 28184 102915 28236
rect 102915 28184 102961 28236
rect 102985 28184 103031 28236
rect 103031 28184 103041 28236
rect 99705 28182 99761 28184
rect 99785 28182 99841 28184
rect 99865 28182 99921 28184
rect 99945 28182 100001 28184
rect 100025 28182 100081 28184
rect 100105 28182 100161 28184
rect 100185 28182 100241 28184
rect 100265 28182 100321 28184
rect 100345 28182 100401 28184
rect 100425 28182 100481 28184
rect 100505 28182 100561 28184
rect 100585 28182 100641 28184
rect 100665 28182 100721 28184
rect 100745 28182 100801 28184
rect 100825 28182 100881 28184
rect 100905 28182 100961 28184
rect 100985 28182 101041 28184
rect 101065 28182 101121 28184
rect 101145 28182 101201 28184
rect 101225 28182 101281 28184
rect 101305 28182 101361 28184
rect 101385 28182 101441 28184
rect 101465 28182 101521 28184
rect 101545 28182 101601 28184
rect 101625 28182 101681 28184
rect 101705 28182 101761 28184
rect 101785 28182 101841 28184
rect 101865 28182 101921 28184
rect 101945 28182 102001 28184
rect 102025 28182 102081 28184
rect 102105 28182 102161 28184
rect 102185 28182 102241 28184
rect 102265 28182 102321 28184
rect 102345 28182 102401 28184
rect 102425 28182 102481 28184
rect 102505 28182 102561 28184
rect 102585 28182 102641 28184
rect 102665 28182 102721 28184
rect 102745 28182 102801 28184
rect 102825 28182 102881 28184
rect 102905 28182 102961 28184
rect 102985 28182 103041 28184
rect 94086 28089 94142 28091
rect 94086 28037 94088 28089
rect 94088 28037 94140 28089
rect 94140 28037 94142 28089
rect 94086 28035 94142 28037
rect 97205 27992 97207 28022
rect 97207 27992 97259 28022
rect 97259 27992 97261 28022
rect 97205 27980 97261 27992
rect 97205 27966 97207 27980
rect 97207 27966 97259 27980
rect 97259 27966 97261 27980
rect 95677 27937 95733 27947
rect 95677 27891 95679 27937
rect 95679 27891 95731 27937
rect 95731 27891 95733 27937
rect 95677 27821 95679 27867
rect 95679 27821 95731 27867
rect 95731 27821 95733 27867
rect 95677 27811 95733 27821
rect 97205 27928 97207 27942
rect 97207 27928 97259 27942
rect 97259 27928 97261 27942
rect 97205 27916 97261 27928
rect 97205 27886 97207 27916
rect 97207 27886 97259 27916
rect 97259 27886 97261 27916
rect 93488 27543 93544 27545
rect 93488 27491 93510 27543
rect 93510 27491 93522 27543
rect 93522 27491 93544 27543
rect 93488 27489 93544 27491
rect 95671 27445 95673 27475
rect 95673 27445 95725 27475
rect 95725 27445 95727 27475
rect 95671 27433 95727 27445
rect 95671 27419 95673 27433
rect 95673 27419 95725 27433
rect 95725 27419 95727 27433
rect 95671 27381 95673 27395
rect 95673 27381 95725 27395
rect 95725 27381 95727 27395
rect 95671 27369 95727 27381
rect 95671 27339 95673 27369
rect 95673 27339 95725 27369
rect 95725 27339 95727 27369
rect 97195 27439 97197 27469
rect 97197 27439 97249 27469
rect 97249 27439 97251 27469
rect 97195 27427 97251 27439
rect 97195 27413 97197 27427
rect 97197 27413 97249 27427
rect 97249 27413 97251 27427
rect 97195 27375 97197 27389
rect 97197 27375 97249 27389
rect 97249 27375 97251 27389
rect 97195 27363 97251 27375
rect 97195 27333 97197 27363
rect 97197 27333 97249 27363
rect 97249 27333 97251 27363
rect 92129 27138 92185 27140
rect 92129 27086 92131 27138
rect 92131 27086 92183 27138
rect 92183 27086 92185 27138
rect 92129 27084 92185 27086
rect 92587 25553 92643 25609
rect 93164 26176 93220 26232
rect 93729 25491 93785 25547
rect 92122 25359 92178 25361
rect 92122 25307 92124 25359
rect 92124 25307 92176 25359
rect 92176 25307 92178 25359
rect 92122 25305 92178 25307
rect 95676 25105 95732 25115
rect 95676 25059 95678 25105
rect 95678 25059 95730 25105
rect 95730 25059 95732 25105
rect 95676 24989 95678 25035
rect 95678 24989 95730 25035
rect 95730 24989 95732 25035
rect 95676 24979 95732 24989
rect 97206 25147 97208 25177
rect 97208 25147 97260 25177
rect 97260 25147 97262 25177
rect 97206 25135 97262 25147
rect 97206 25121 97208 25135
rect 97208 25121 97260 25135
rect 97260 25121 97262 25135
rect 97206 25083 97208 25097
rect 97208 25083 97260 25097
rect 97260 25083 97262 25097
rect 97206 25071 97262 25083
rect 97206 25041 97208 25071
rect 97208 25041 97260 25071
rect 97260 25041 97262 25071
rect 93402 24955 93458 24957
rect 93482 24955 93538 24957
rect 93562 24955 93618 24957
rect 93402 24903 93420 24955
rect 93420 24903 93458 24955
rect 93482 24903 93484 24955
rect 93484 24903 93536 24955
rect 93536 24903 93538 24955
rect 93562 24903 93600 24955
rect 93600 24903 93618 24955
rect 93402 24901 93458 24903
rect 93482 24901 93538 24903
rect 93562 24901 93618 24903
rect 95674 24589 95676 24619
rect 95676 24589 95728 24619
rect 95728 24589 95730 24619
rect 95674 24577 95730 24589
rect 95674 24563 95676 24577
rect 95676 24563 95728 24577
rect 95728 24563 95730 24577
rect 95674 24525 95676 24539
rect 95676 24525 95728 24539
rect 95728 24525 95730 24539
rect 95674 24513 95730 24525
rect 95674 24483 95676 24513
rect 95676 24483 95728 24513
rect 95728 24483 95730 24513
rect 97193 24602 97195 24632
rect 97195 24602 97247 24632
rect 97247 24602 97249 24632
rect 97193 24590 97249 24602
rect 97193 24576 97195 24590
rect 97195 24576 97247 24590
rect 97247 24576 97249 24590
rect 97193 24538 97195 24552
rect 97195 24538 97247 24552
rect 97247 24538 97249 24552
rect 97193 24526 97249 24538
rect 97193 24496 97195 24526
rect 97195 24496 97247 24526
rect 97247 24496 97249 24526
rect 93472 24414 93528 24416
rect 93552 24414 93608 24416
rect 93472 24362 93482 24414
rect 93482 24362 93528 24414
rect 93552 24362 93598 24414
rect 93598 24362 93608 24414
rect 93472 24360 93528 24362
rect 93552 24360 93608 24362
rect 57420 24229 78196 24239
rect 57420 24113 57446 24229
rect 57446 24113 78170 24229
rect 78170 24113 78196 24229
rect 57420 24103 78196 24113
rect 92126 24299 92182 24301
rect 92126 24247 92128 24299
rect 92128 24247 92180 24299
rect 92180 24247 92182 24299
rect 92126 24245 92182 24247
rect 99730 24302 99786 24304
rect 99810 24302 99866 24304
rect 99890 24302 99946 24304
rect 99970 24302 100026 24304
rect 100050 24302 100106 24304
rect 100130 24302 100186 24304
rect 100210 24302 100266 24304
rect 100290 24302 100346 24304
rect 100370 24302 100426 24304
rect 100450 24302 100506 24304
rect 100530 24302 100586 24304
rect 100610 24302 100666 24304
rect 100690 24302 100746 24304
rect 100770 24302 100826 24304
rect 100850 24302 100906 24304
rect 100930 24302 100986 24304
rect 101010 24302 101066 24304
rect 101090 24302 101146 24304
rect 101170 24302 101226 24304
rect 101250 24302 101306 24304
rect 101330 24302 101386 24304
rect 101410 24302 101466 24304
rect 101490 24302 101546 24304
rect 101570 24302 101626 24304
rect 101650 24302 101706 24304
rect 101730 24302 101786 24304
rect 101810 24302 101866 24304
rect 101890 24302 101946 24304
rect 101970 24302 102026 24304
rect 102050 24302 102106 24304
rect 102130 24302 102186 24304
rect 102210 24302 102266 24304
rect 102290 24302 102346 24304
rect 102370 24302 102426 24304
rect 102450 24302 102506 24304
rect 102530 24302 102586 24304
rect 102610 24302 102666 24304
rect 102690 24302 102746 24304
rect 102770 24302 102826 24304
rect 102850 24302 102906 24304
rect 102930 24302 102986 24304
rect 99730 24250 99752 24302
rect 99752 24250 99764 24302
rect 99764 24250 99786 24302
rect 99810 24250 99816 24302
rect 99816 24250 99828 24302
rect 99828 24250 99866 24302
rect 99890 24250 99892 24302
rect 99892 24250 99944 24302
rect 99944 24250 99946 24302
rect 99970 24250 100008 24302
rect 100008 24250 100020 24302
rect 100020 24250 100026 24302
rect 100050 24250 100072 24302
rect 100072 24250 100084 24302
rect 100084 24250 100106 24302
rect 100130 24250 100136 24302
rect 100136 24250 100148 24302
rect 100148 24250 100186 24302
rect 100210 24250 100212 24302
rect 100212 24250 100264 24302
rect 100264 24250 100266 24302
rect 100290 24250 100328 24302
rect 100328 24250 100340 24302
rect 100340 24250 100346 24302
rect 100370 24250 100392 24302
rect 100392 24250 100404 24302
rect 100404 24250 100426 24302
rect 100450 24250 100456 24302
rect 100456 24250 100468 24302
rect 100468 24250 100506 24302
rect 100530 24250 100532 24302
rect 100532 24250 100584 24302
rect 100584 24250 100586 24302
rect 100610 24250 100648 24302
rect 100648 24250 100660 24302
rect 100660 24250 100666 24302
rect 100690 24250 100712 24302
rect 100712 24250 100724 24302
rect 100724 24250 100746 24302
rect 100770 24250 100776 24302
rect 100776 24250 100788 24302
rect 100788 24250 100826 24302
rect 100850 24250 100852 24302
rect 100852 24250 100904 24302
rect 100904 24250 100906 24302
rect 100930 24250 100968 24302
rect 100968 24250 100980 24302
rect 100980 24250 100986 24302
rect 101010 24250 101032 24302
rect 101032 24250 101044 24302
rect 101044 24250 101066 24302
rect 101090 24250 101096 24302
rect 101096 24250 101108 24302
rect 101108 24250 101146 24302
rect 101170 24250 101172 24302
rect 101172 24250 101224 24302
rect 101224 24250 101226 24302
rect 101250 24250 101288 24302
rect 101288 24250 101300 24302
rect 101300 24250 101306 24302
rect 101330 24250 101352 24302
rect 101352 24250 101364 24302
rect 101364 24250 101386 24302
rect 101410 24250 101416 24302
rect 101416 24250 101428 24302
rect 101428 24250 101466 24302
rect 101490 24250 101492 24302
rect 101492 24250 101544 24302
rect 101544 24250 101546 24302
rect 101570 24250 101608 24302
rect 101608 24250 101620 24302
rect 101620 24250 101626 24302
rect 101650 24250 101672 24302
rect 101672 24250 101684 24302
rect 101684 24250 101706 24302
rect 101730 24250 101736 24302
rect 101736 24250 101748 24302
rect 101748 24250 101786 24302
rect 101810 24250 101812 24302
rect 101812 24250 101864 24302
rect 101864 24250 101866 24302
rect 101890 24250 101928 24302
rect 101928 24250 101940 24302
rect 101940 24250 101946 24302
rect 101970 24250 101992 24302
rect 101992 24250 102004 24302
rect 102004 24250 102026 24302
rect 102050 24250 102056 24302
rect 102056 24250 102068 24302
rect 102068 24250 102106 24302
rect 102130 24250 102132 24302
rect 102132 24250 102184 24302
rect 102184 24250 102186 24302
rect 102210 24250 102248 24302
rect 102248 24250 102260 24302
rect 102260 24250 102266 24302
rect 102290 24250 102312 24302
rect 102312 24250 102324 24302
rect 102324 24250 102346 24302
rect 102370 24250 102376 24302
rect 102376 24250 102388 24302
rect 102388 24250 102426 24302
rect 102450 24250 102452 24302
rect 102452 24250 102504 24302
rect 102504 24250 102506 24302
rect 102530 24250 102568 24302
rect 102568 24250 102580 24302
rect 102580 24250 102586 24302
rect 102610 24250 102632 24302
rect 102632 24250 102644 24302
rect 102644 24250 102666 24302
rect 102690 24250 102696 24302
rect 102696 24250 102708 24302
rect 102708 24250 102746 24302
rect 102770 24250 102772 24302
rect 102772 24250 102824 24302
rect 102824 24250 102826 24302
rect 102850 24250 102888 24302
rect 102888 24250 102900 24302
rect 102900 24250 102906 24302
rect 102930 24250 102952 24302
rect 102952 24250 102964 24302
rect 102964 24250 102986 24302
rect 99730 24248 99786 24250
rect 99810 24248 99866 24250
rect 99890 24248 99946 24250
rect 99970 24248 100026 24250
rect 100050 24248 100106 24250
rect 100130 24248 100186 24250
rect 100210 24248 100266 24250
rect 100290 24248 100346 24250
rect 100370 24248 100426 24250
rect 100450 24248 100506 24250
rect 100530 24248 100586 24250
rect 100610 24248 100666 24250
rect 100690 24248 100746 24250
rect 100770 24248 100826 24250
rect 100850 24248 100906 24250
rect 100930 24248 100986 24250
rect 101010 24248 101066 24250
rect 101090 24248 101146 24250
rect 101170 24248 101226 24250
rect 101250 24248 101306 24250
rect 101330 24248 101386 24250
rect 101410 24248 101466 24250
rect 101490 24248 101546 24250
rect 101570 24248 101626 24250
rect 101650 24248 101706 24250
rect 101730 24248 101786 24250
rect 101810 24248 101866 24250
rect 101890 24248 101946 24250
rect 101970 24248 102026 24250
rect 102050 24248 102106 24250
rect 102130 24248 102186 24250
rect 102210 24248 102266 24250
rect 102290 24248 102346 24250
rect 102370 24248 102426 24250
rect 102450 24248 102506 24250
rect 102530 24248 102586 24250
rect 102610 24248 102666 24250
rect 102690 24248 102746 24250
rect 102770 24248 102826 24250
rect 102850 24248 102906 24250
rect 102930 24248 102986 24250
rect 92125 24030 92181 24032
rect 92125 23978 92127 24030
rect 92127 23978 92179 24030
rect 92179 23978 92181 24030
rect 92125 23976 92181 23978
rect 93460 23866 93516 23868
rect 93460 23814 93462 23866
rect 93462 23814 93514 23866
rect 93514 23814 93516 23866
rect 93460 23812 93516 23814
rect 95676 23732 95678 23754
rect 95678 23732 95730 23754
rect 95730 23732 95732 23754
rect 95676 23720 95732 23732
rect 95676 23698 95678 23720
rect 95678 23698 95730 23720
rect 95730 23698 95732 23720
rect 97198 23811 97200 23841
rect 97200 23811 97252 23841
rect 97252 23811 97254 23841
rect 97198 23799 97254 23811
rect 97198 23785 97200 23799
rect 97200 23785 97252 23799
rect 97252 23785 97254 23799
rect 97198 23747 97200 23761
rect 97200 23747 97252 23761
rect 97252 23747 97254 23761
rect 97198 23735 97254 23747
rect 97198 23705 97200 23735
rect 97200 23705 97252 23735
rect 97252 23705 97254 23735
rect 94085 23325 94141 23327
rect 94085 23273 94087 23325
rect 94087 23273 94139 23325
rect 94139 23273 94141 23325
rect 94085 23271 94141 23273
rect 95669 23258 95671 23288
rect 95671 23258 95723 23288
rect 95723 23258 95725 23288
rect 95669 23246 95725 23258
rect 95669 23232 95671 23246
rect 95671 23232 95723 23246
rect 95723 23232 95725 23246
rect 95669 23194 95671 23208
rect 95671 23194 95723 23208
rect 95723 23194 95725 23208
rect 95669 23182 95725 23194
rect 95669 23152 95671 23182
rect 95671 23152 95723 23182
rect 95723 23152 95725 23182
rect 97198 23255 97200 23285
rect 97200 23255 97252 23285
rect 97252 23255 97254 23285
rect 97198 23243 97254 23255
rect 97198 23229 97200 23243
rect 97200 23229 97252 23243
rect 97252 23229 97254 23243
rect 97198 23191 97200 23205
rect 97200 23191 97252 23205
rect 97252 23191 97254 23205
rect 97198 23179 97254 23191
rect 97198 23149 97200 23179
rect 97200 23149 97252 23179
rect 97252 23149 97254 23179
rect 92125 22961 92181 22963
rect 92125 22909 92127 22961
rect 92127 22909 92179 22961
rect 92179 22909 92181 22961
rect 92125 22907 92181 22909
rect 93085 22783 93141 22785
rect 93165 22783 93221 22785
rect 93085 22731 93095 22783
rect 93095 22731 93141 22783
rect 93165 22731 93211 22783
rect 93211 22731 93221 22783
rect 93085 22729 93141 22731
rect 93165 22729 93221 22731
rect 104593 22854 104809 22872
rect 104593 22674 104611 22854
rect 104611 22674 104791 22854
rect 104791 22674 104809 22854
rect 104593 22656 104809 22674
rect 92122 22638 92178 22640
rect 92122 22586 92124 22638
rect 92124 22586 92176 22638
rect 92176 22586 92178 22638
rect 92122 22584 92178 22586
rect 95677 22342 95679 22364
rect 95679 22342 95731 22364
rect 95731 22342 95733 22364
rect 95677 22330 95733 22342
rect 95677 22308 95679 22330
rect 95679 22308 95731 22330
rect 95731 22308 95733 22330
rect 97215 22431 97217 22461
rect 97217 22431 97269 22461
rect 97269 22431 97271 22461
rect 97215 22419 97271 22431
rect 97215 22405 97217 22419
rect 97217 22405 97269 22419
rect 97269 22405 97271 22419
rect 97215 22367 97217 22381
rect 97217 22367 97269 22381
rect 97269 22367 97271 22381
rect 97215 22355 97271 22367
rect 97215 22325 97217 22355
rect 97217 22325 97269 22355
rect 97269 22325 97271 22355
rect 93610 22235 93666 22237
rect 93690 22235 93746 22237
rect 93770 22235 93826 22237
rect 93610 22183 93628 22235
rect 93628 22183 93666 22235
rect 93690 22183 93692 22235
rect 93692 22183 93744 22235
rect 93744 22183 93746 22235
rect 93770 22183 93808 22235
rect 93808 22183 93826 22235
rect 93610 22181 93666 22183
rect 93690 22181 93746 22183
rect 93770 22181 93826 22183
rect 95668 21905 95670 21935
rect 95670 21905 95722 21935
rect 95722 21905 95724 21935
rect 95668 21893 95724 21905
rect 95668 21879 95670 21893
rect 95670 21879 95722 21893
rect 95722 21879 95724 21893
rect 95668 21841 95670 21855
rect 95670 21841 95722 21855
rect 95722 21841 95724 21855
rect 95668 21829 95724 21841
rect 95668 21799 95670 21829
rect 95670 21799 95722 21829
rect 95722 21799 95724 21829
rect 97198 21883 97200 21913
rect 97200 21883 97252 21913
rect 97252 21883 97254 21913
rect 97198 21871 97254 21883
rect 97198 21857 97200 21871
rect 97200 21857 97252 21871
rect 97252 21857 97254 21871
rect 97198 21819 97200 21833
rect 97200 21819 97252 21833
rect 97252 21819 97254 21833
rect 97198 21807 97254 21819
rect 97198 21777 97200 21807
rect 97200 21777 97252 21807
rect 97252 21777 97254 21807
rect 93462 21692 93518 21694
rect 93542 21692 93598 21694
rect 93462 21640 93472 21692
rect 93472 21640 93518 21692
rect 93542 21640 93588 21692
rect 93588 21640 93598 21692
rect 93462 21638 93518 21640
rect 93542 21638 93598 21640
rect 92133 21568 92189 21570
rect 92133 21516 92135 21568
rect 92135 21516 92187 21568
rect 92187 21516 92189 21568
rect 92133 21514 92189 21516
rect 92122 21263 92178 21265
rect 92122 21211 92124 21263
rect 92124 21211 92176 21263
rect 92176 21211 92178 21263
rect 92122 21209 92178 21211
rect 99686 21296 99742 21298
rect 99766 21296 99822 21298
rect 99846 21296 99902 21298
rect 99926 21296 99982 21298
rect 100006 21296 100062 21298
rect 100086 21296 100142 21298
rect 100166 21296 100222 21298
rect 100246 21296 100302 21298
rect 100326 21296 100382 21298
rect 100406 21296 100462 21298
rect 100486 21296 100542 21298
rect 100566 21296 100622 21298
rect 100646 21296 100702 21298
rect 100726 21296 100782 21298
rect 100806 21296 100862 21298
rect 100886 21296 100942 21298
rect 100966 21296 101022 21298
rect 101046 21296 101102 21298
rect 101126 21296 101182 21298
rect 101206 21296 101262 21298
rect 101286 21296 101342 21298
rect 101366 21296 101422 21298
rect 101446 21296 101502 21298
rect 101526 21296 101582 21298
rect 101606 21296 101662 21298
rect 101686 21296 101742 21298
rect 101766 21296 101822 21298
rect 101846 21296 101902 21298
rect 101926 21296 101982 21298
rect 102006 21296 102062 21298
rect 102086 21296 102142 21298
rect 102166 21296 102222 21298
rect 102246 21296 102302 21298
rect 102326 21296 102382 21298
rect 102406 21296 102462 21298
rect 102486 21296 102542 21298
rect 102566 21296 102622 21298
rect 102646 21296 102702 21298
rect 102726 21296 102782 21298
rect 102806 21296 102862 21298
rect 102886 21296 102942 21298
rect 102966 21296 103022 21298
rect 99686 21244 99696 21296
rect 99696 21244 99742 21296
rect 99766 21244 99812 21296
rect 99812 21244 99822 21296
rect 99846 21244 99876 21296
rect 99876 21244 99888 21296
rect 99888 21244 99902 21296
rect 99926 21244 99940 21296
rect 99940 21244 99952 21296
rect 99952 21244 99982 21296
rect 100006 21244 100016 21296
rect 100016 21244 100062 21296
rect 100086 21244 100132 21296
rect 100132 21244 100142 21296
rect 100166 21244 100196 21296
rect 100196 21244 100208 21296
rect 100208 21244 100222 21296
rect 100246 21244 100260 21296
rect 100260 21244 100272 21296
rect 100272 21244 100302 21296
rect 100326 21244 100336 21296
rect 100336 21244 100382 21296
rect 100406 21244 100452 21296
rect 100452 21244 100462 21296
rect 100486 21244 100516 21296
rect 100516 21244 100528 21296
rect 100528 21244 100542 21296
rect 100566 21244 100580 21296
rect 100580 21244 100592 21296
rect 100592 21244 100622 21296
rect 100646 21244 100656 21296
rect 100656 21244 100702 21296
rect 100726 21244 100772 21296
rect 100772 21244 100782 21296
rect 100806 21244 100836 21296
rect 100836 21244 100848 21296
rect 100848 21244 100862 21296
rect 100886 21244 100900 21296
rect 100900 21244 100912 21296
rect 100912 21244 100942 21296
rect 100966 21244 100976 21296
rect 100976 21244 101022 21296
rect 101046 21244 101092 21296
rect 101092 21244 101102 21296
rect 101126 21244 101156 21296
rect 101156 21244 101168 21296
rect 101168 21244 101182 21296
rect 101206 21244 101220 21296
rect 101220 21244 101232 21296
rect 101232 21244 101262 21296
rect 101286 21244 101296 21296
rect 101296 21244 101342 21296
rect 101366 21244 101412 21296
rect 101412 21244 101422 21296
rect 101446 21244 101476 21296
rect 101476 21244 101488 21296
rect 101488 21244 101502 21296
rect 101526 21244 101540 21296
rect 101540 21244 101552 21296
rect 101552 21244 101582 21296
rect 101606 21244 101616 21296
rect 101616 21244 101662 21296
rect 101686 21244 101732 21296
rect 101732 21244 101742 21296
rect 101766 21244 101796 21296
rect 101796 21244 101808 21296
rect 101808 21244 101822 21296
rect 101846 21244 101860 21296
rect 101860 21244 101872 21296
rect 101872 21244 101902 21296
rect 101926 21244 101936 21296
rect 101936 21244 101982 21296
rect 102006 21244 102052 21296
rect 102052 21244 102062 21296
rect 102086 21244 102116 21296
rect 102116 21244 102128 21296
rect 102128 21244 102142 21296
rect 102166 21244 102180 21296
rect 102180 21244 102192 21296
rect 102192 21244 102222 21296
rect 102246 21244 102256 21296
rect 102256 21244 102302 21296
rect 102326 21244 102372 21296
rect 102372 21244 102382 21296
rect 102406 21244 102436 21296
rect 102436 21244 102448 21296
rect 102448 21244 102462 21296
rect 102486 21244 102500 21296
rect 102500 21244 102512 21296
rect 102512 21244 102542 21296
rect 102566 21244 102576 21296
rect 102576 21244 102622 21296
rect 102646 21244 102692 21296
rect 102692 21244 102702 21296
rect 102726 21244 102756 21296
rect 102756 21244 102768 21296
rect 102768 21244 102782 21296
rect 102806 21244 102820 21296
rect 102820 21244 102832 21296
rect 102832 21244 102862 21296
rect 102886 21244 102896 21296
rect 102896 21244 102942 21296
rect 102966 21244 103012 21296
rect 103012 21244 103022 21296
rect 99686 21242 99742 21244
rect 99766 21242 99822 21244
rect 99846 21242 99902 21244
rect 99926 21242 99982 21244
rect 100006 21242 100062 21244
rect 100086 21242 100142 21244
rect 100166 21242 100222 21244
rect 100246 21242 100302 21244
rect 100326 21242 100382 21244
rect 100406 21242 100462 21244
rect 100486 21242 100542 21244
rect 100566 21242 100622 21244
rect 100646 21242 100702 21244
rect 100726 21242 100782 21244
rect 100806 21242 100862 21244
rect 100886 21242 100942 21244
rect 100966 21242 101022 21244
rect 101046 21242 101102 21244
rect 101126 21242 101182 21244
rect 101206 21242 101262 21244
rect 101286 21242 101342 21244
rect 101366 21242 101422 21244
rect 101446 21242 101502 21244
rect 101526 21242 101582 21244
rect 101606 21242 101662 21244
rect 101686 21242 101742 21244
rect 101766 21242 101822 21244
rect 101846 21242 101902 21244
rect 101926 21242 101982 21244
rect 102006 21242 102062 21244
rect 102086 21242 102142 21244
rect 102166 21242 102222 21244
rect 102246 21242 102302 21244
rect 102326 21242 102382 21244
rect 102406 21242 102462 21244
rect 102486 21242 102542 21244
rect 102566 21242 102622 21244
rect 102646 21242 102702 21244
rect 102726 21242 102782 21244
rect 102806 21242 102862 21244
rect 102886 21242 102942 21244
rect 102966 21242 103022 21244
rect 94086 21149 94142 21151
rect 94086 21097 94088 21149
rect 94088 21097 94140 21149
rect 94140 21097 94142 21149
rect 94086 21095 94142 21097
rect 97205 21052 97207 21082
rect 97207 21052 97259 21082
rect 97259 21052 97261 21082
rect 97205 21040 97261 21052
rect 97205 21026 97207 21040
rect 97207 21026 97259 21040
rect 97259 21026 97261 21040
rect 95677 20997 95733 21007
rect 95677 20951 95679 20997
rect 95679 20951 95731 20997
rect 95731 20951 95733 20997
rect 95677 20881 95679 20927
rect 95679 20881 95731 20927
rect 95731 20881 95733 20927
rect 95677 20871 95733 20881
rect 97205 20988 97207 21002
rect 97207 20988 97259 21002
rect 97259 20988 97261 21002
rect 97205 20976 97261 20988
rect 97205 20946 97207 20976
rect 97207 20946 97259 20976
rect 97259 20946 97261 20976
rect 93488 20603 93544 20605
rect 93488 20551 93510 20603
rect 93510 20551 93522 20603
rect 93522 20551 93544 20603
rect 93488 20549 93544 20551
rect 95671 20505 95673 20535
rect 95673 20505 95725 20535
rect 95725 20505 95727 20535
rect 95671 20493 95727 20505
rect 95671 20479 95673 20493
rect 95673 20479 95725 20493
rect 95725 20479 95727 20493
rect 95671 20441 95673 20455
rect 95673 20441 95725 20455
rect 95725 20441 95727 20455
rect 95671 20429 95727 20441
rect 95671 20399 95673 20429
rect 95673 20399 95725 20429
rect 95725 20399 95727 20429
rect 97195 20499 97197 20529
rect 97197 20499 97249 20529
rect 97249 20499 97251 20529
rect 97195 20487 97251 20499
rect 97195 20473 97197 20487
rect 97197 20473 97249 20487
rect 97249 20473 97251 20487
rect 97195 20435 97197 20449
rect 97197 20435 97249 20449
rect 97249 20435 97251 20449
rect 97195 20423 97251 20435
rect 97195 20393 97197 20423
rect 97197 20393 97249 20423
rect 97249 20393 97251 20423
rect 92129 20198 92185 20200
rect 92129 20146 92131 20198
rect 92131 20146 92183 20198
rect 92183 20146 92185 20198
rect 92129 20144 92185 20146
rect 53517 17172 53573 17174
rect 53517 17120 53519 17172
rect 53519 17120 53571 17172
rect 53571 17120 53573 17172
rect 53517 17118 53573 17120
rect 53517 17056 53519 17094
rect 53519 17056 53571 17094
rect 53571 17056 53573 17094
rect 53517 17044 53573 17056
rect 53517 17038 53519 17044
rect 53519 17038 53571 17044
rect 53571 17038 53573 17044
rect 53517 16992 53519 17014
rect 53519 16992 53571 17014
rect 53571 16992 53573 17014
rect 53517 16980 53573 16992
rect 53517 16958 53519 16980
rect 53519 16958 53571 16980
rect 53571 16958 53573 16980
rect 53517 16928 53519 16934
rect 53519 16928 53571 16934
rect 53571 16928 53573 16934
rect 53517 16916 53573 16928
rect 53517 16878 53519 16916
rect 53519 16878 53571 16916
rect 53571 16878 53573 16916
rect 53517 16852 53573 16854
rect 53517 16800 53519 16852
rect 53519 16800 53571 16852
rect 53571 16800 53573 16852
rect 53517 16798 53573 16800
rect 53517 16736 53519 16774
rect 53519 16736 53571 16774
rect 53571 16736 53573 16774
rect 53517 16724 53573 16736
rect 53517 16718 53519 16724
rect 53519 16718 53571 16724
rect 53571 16718 53573 16724
rect 53517 16672 53519 16694
rect 53519 16672 53571 16694
rect 53571 16672 53573 16694
rect 53517 16660 53573 16672
rect 53517 16638 53519 16660
rect 53519 16638 53571 16660
rect 53571 16638 53573 16660
rect 53517 16608 53519 16614
rect 53519 16608 53571 16614
rect 53571 16608 53573 16614
rect 53517 16596 53573 16608
rect 53517 16558 53519 16596
rect 53519 16558 53571 16596
rect 53571 16558 53573 16596
rect 53517 16532 53573 16534
rect 53517 16480 53519 16532
rect 53519 16480 53571 16532
rect 53571 16480 53573 16532
rect 53517 16478 53573 16480
rect 53517 16416 53519 16454
rect 53519 16416 53571 16454
rect 53571 16416 53573 16454
rect 53517 16404 53573 16416
rect 53517 16398 53519 16404
rect 53519 16398 53571 16404
rect 53571 16398 53573 16404
rect 53517 16352 53519 16374
rect 53519 16352 53571 16374
rect 53571 16352 53573 16374
rect 53517 16340 53573 16352
rect 53517 16318 53519 16340
rect 53519 16318 53571 16340
rect 53571 16318 53573 16340
rect 53517 16288 53519 16294
rect 53519 16288 53571 16294
rect 53571 16288 53573 16294
rect 53517 16276 53573 16288
rect 53517 16238 53519 16276
rect 53519 16238 53571 16276
rect 53571 16238 53573 16276
rect 53517 16212 53573 16214
rect 53517 16160 53519 16212
rect 53519 16160 53571 16212
rect 53571 16160 53573 16212
rect 53517 16158 53573 16160
rect 53517 16096 53519 16134
rect 53519 16096 53571 16134
rect 53571 16096 53573 16134
rect 53517 16084 53573 16096
rect 53517 16078 53519 16084
rect 53519 16078 53571 16084
rect 53571 16078 53573 16084
rect 53517 16032 53519 16054
rect 53519 16032 53571 16054
rect 53571 16032 53573 16054
rect 53517 16020 53573 16032
rect 53517 15998 53519 16020
rect 53519 15998 53571 16020
rect 53571 15998 53573 16020
rect 53517 15968 53519 15974
rect 53519 15968 53571 15974
rect 53571 15968 53573 15974
rect 53517 15956 53573 15968
rect 53517 15918 53519 15956
rect 53519 15918 53571 15956
rect 53571 15918 53573 15956
rect 53517 15892 53573 15894
rect 53517 15840 53519 15892
rect 53519 15840 53571 15892
rect 53571 15840 53573 15892
rect 53517 15838 53573 15840
rect 53517 15776 53519 15814
rect 53519 15776 53571 15814
rect 53571 15776 53573 15814
rect 53517 15764 53573 15776
rect 53517 15758 53519 15764
rect 53519 15758 53571 15764
rect 53571 15758 53573 15764
rect 53517 15712 53519 15734
rect 53519 15712 53571 15734
rect 53571 15712 53573 15734
rect 53517 15700 53573 15712
rect 53517 15678 53519 15700
rect 53519 15678 53571 15700
rect 53571 15678 53573 15700
rect 53517 15648 53519 15654
rect 53519 15648 53571 15654
rect 53571 15648 53573 15654
rect 53517 15636 53573 15648
rect 53517 15598 53519 15636
rect 53519 15598 53571 15636
rect 53571 15598 53573 15636
rect 53517 15572 53573 15574
rect 53517 15520 53519 15572
rect 53519 15520 53571 15572
rect 53571 15520 53573 15572
rect 53517 15518 53573 15520
rect 53517 15456 53519 15494
rect 53519 15456 53571 15494
rect 53571 15456 53573 15494
rect 53517 15444 53573 15456
rect 53517 15438 53519 15444
rect 53519 15438 53571 15444
rect 53571 15438 53573 15444
rect 53517 15392 53519 15414
rect 53519 15392 53571 15414
rect 53571 15392 53573 15414
rect 53517 15380 53573 15392
rect 53517 15358 53519 15380
rect 53519 15358 53571 15380
rect 53571 15358 53573 15380
rect 53517 15328 53519 15334
rect 53519 15328 53571 15334
rect 53571 15328 53573 15334
rect 53517 15316 53573 15328
rect 53517 15278 53519 15316
rect 53519 15278 53571 15316
rect 53571 15278 53573 15316
rect 53517 15252 53573 15254
rect 53517 15200 53519 15252
rect 53519 15200 53571 15252
rect 53571 15200 53573 15252
rect 53517 15198 53573 15200
rect 53517 15136 53519 15174
rect 53519 15136 53571 15174
rect 53571 15136 53573 15174
rect 53517 15124 53573 15136
rect 53517 15118 53519 15124
rect 53519 15118 53571 15124
rect 53571 15118 53573 15124
rect 53517 15072 53519 15094
rect 53519 15072 53571 15094
rect 53571 15072 53573 15094
rect 53517 15060 53573 15072
rect 53517 15038 53519 15060
rect 53519 15038 53571 15060
rect 53571 15038 53573 15060
rect 53517 15008 53519 15014
rect 53519 15008 53571 15014
rect 53571 15008 53573 15014
rect 53517 14996 53573 15008
rect 53517 14958 53519 14996
rect 53519 14958 53571 14996
rect 53571 14958 53573 14996
rect 53517 14932 53573 14934
rect 53517 14880 53519 14932
rect 53519 14880 53571 14932
rect 53571 14880 53573 14932
rect 53517 14878 53573 14880
rect 53517 14816 53519 14854
rect 53519 14816 53571 14854
rect 53571 14816 53573 14854
rect 53517 14804 53573 14816
rect 53517 14798 53519 14804
rect 53519 14798 53571 14804
rect 53571 14798 53573 14804
rect 53517 14752 53519 14774
rect 53519 14752 53571 14774
rect 53571 14752 53573 14774
rect 53517 14740 53573 14752
rect 53517 14718 53519 14740
rect 53519 14718 53571 14740
rect 53571 14718 53573 14740
rect 53517 14688 53519 14694
rect 53519 14688 53571 14694
rect 53571 14688 53573 14694
rect 53517 14676 53573 14688
rect 53517 14638 53519 14676
rect 53519 14638 53571 14676
rect 53571 14638 53573 14676
rect 53517 14612 53573 14614
rect 53517 14560 53519 14612
rect 53519 14560 53571 14612
rect 53571 14560 53573 14612
rect 53517 14558 53573 14560
rect 53517 14496 53519 14534
rect 53519 14496 53571 14534
rect 53571 14496 53573 14534
rect 53517 14484 53573 14496
rect 53517 14478 53519 14484
rect 53519 14478 53571 14484
rect 53571 14478 53573 14484
rect 53517 14432 53519 14454
rect 53519 14432 53571 14454
rect 53571 14432 53573 14454
rect 53517 14420 53573 14432
rect 53517 14398 53519 14420
rect 53519 14398 53571 14420
rect 53571 14398 53573 14420
rect 53517 14368 53519 14374
rect 53519 14368 53571 14374
rect 53571 14368 53573 14374
rect 53517 14356 53573 14368
rect 53517 14318 53519 14356
rect 53519 14318 53571 14356
rect 53571 14318 53573 14356
rect 53517 14292 53573 14294
rect 53517 14240 53519 14292
rect 53519 14240 53571 14292
rect 53571 14240 53573 14292
rect 53517 14238 53573 14240
rect 53517 14176 53519 14214
rect 53519 14176 53571 14214
rect 53571 14176 53573 14214
rect 53517 14164 53573 14176
rect 53517 14158 53519 14164
rect 53519 14158 53571 14164
rect 53571 14158 53573 14164
rect 53517 14112 53519 14134
rect 53519 14112 53571 14134
rect 53571 14112 53573 14134
rect 53517 14100 53573 14112
rect 53517 14078 53519 14100
rect 53519 14078 53571 14100
rect 53571 14078 53573 14100
rect 53517 14048 53519 14054
rect 53519 14048 53571 14054
rect 53571 14048 53573 14054
rect 53517 14036 53573 14048
rect 53517 13998 53519 14036
rect 53519 13998 53571 14036
rect 53571 13998 53573 14036
rect 53517 13972 53573 13974
rect 53517 13920 53519 13972
rect 53519 13920 53571 13972
rect 53571 13920 53573 13972
rect 53517 13918 53573 13920
rect 56523 17165 56579 17167
rect 56523 17113 56525 17165
rect 56525 17113 56577 17165
rect 56577 17113 56579 17165
rect 56523 17111 56579 17113
rect 56523 17049 56525 17087
rect 56525 17049 56577 17087
rect 56577 17049 56579 17087
rect 56523 17037 56579 17049
rect 56523 17031 56525 17037
rect 56525 17031 56577 17037
rect 56577 17031 56579 17037
rect 56523 16985 56525 17007
rect 56525 16985 56577 17007
rect 56577 16985 56579 17007
rect 56523 16973 56579 16985
rect 56523 16951 56525 16973
rect 56525 16951 56577 16973
rect 56577 16951 56579 16973
rect 56523 16921 56525 16927
rect 56525 16921 56577 16927
rect 56577 16921 56579 16927
rect 56523 16909 56579 16921
rect 56523 16871 56525 16909
rect 56525 16871 56577 16909
rect 56577 16871 56579 16909
rect 56523 16845 56579 16847
rect 56523 16793 56525 16845
rect 56525 16793 56577 16845
rect 56577 16793 56579 16845
rect 56523 16791 56579 16793
rect 56523 16729 56525 16767
rect 56525 16729 56577 16767
rect 56577 16729 56579 16767
rect 56523 16717 56579 16729
rect 56523 16711 56525 16717
rect 56525 16711 56577 16717
rect 56577 16711 56579 16717
rect 56523 16665 56525 16687
rect 56525 16665 56577 16687
rect 56577 16665 56579 16687
rect 56523 16653 56579 16665
rect 56523 16631 56525 16653
rect 56525 16631 56577 16653
rect 56577 16631 56579 16653
rect 56523 16601 56525 16607
rect 56525 16601 56577 16607
rect 56577 16601 56579 16607
rect 56523 16589 56579 16601
rect 56523 16551 56525 16589
rect 56525 16551 56577 16589
rect 56577 16551 56579 16589
rect 56523 16525 56579 16527
rect 56523 16473 56525 16525
rect 56525 16473 56577 16525
rect 56577 16473 56579 16525
rect 56523 16471 56579 16473
rect 56523 16409 56525 16447
rect 56525 16409 56577 16447
rect 56577 16409 56579 16447
rect 56523 16397 56579 16409
rect 56523 16391 56525 16397
rect 56525 16391 56577 16397
rect 56577 16391 56579 16397
rect 56523 16345 56525 16367
rect 56525 16345 56577 16367
rect 56577 16345 56579 16367
rect 56523 16333 56579 16345
rect 56523 16311 56525 16333
rect 56525 16311 56577 16333
rect 56577 16311 56579 16333
rect 56523 16281 56525 16287
rect 56525 16281 56577 16287
rect 56577 16281 56579 16287
rect 56523 16269 56579 16281
rect 56523 16231 56525 16269
rect 56525 16231 56577 16269
rect 56577 16231 56579 16269
rect 56523 16205 56579 16207
rect 56523 16153 56525 16205
rect 56525 16153 56577 16205
rect 56577 16153 56579 16205
rect 56523 16151 56579 16153
rect 56523 16089 56525 16127
rect 56525 16089 56577 16127
rect 56577 16089 56579 16127
rect 56523 16077 56579 16089
rect 56523 16071 56525 16077
rect 56525 16071 56577 16077
rect 56577 16071 56579 16077
rect 56523 16025 56525 16047
rect 56525 16025 56577 16047
rect 56577 16025 56579 16047
rect 56523 16013 56579 16025
rect 56523 15991 56525 16013
rect 56525 15991 56577 16013
rect 56577 15991 56579 16013
rect 56523 15961 56525 15967
rect 56525 15961 56577 15967
rect 56577 15961 56579 15967
rect 56523 15949 56579 15961
rect 56523 15911 56525 15949
rect 56525 15911 56577 15949
rect 56577 15911 56579 15949
rect 56523 15885 56579 15887
rect 56523 15833 56525 15885
rect 56525 15833 56577 15885
rect 56577 15833 56579 15885
rect 56523 15831 56579 15833
rect 56523 15769 56525 15807
rect 56525 15769 56577 15807
rect 56577 15769 56579 15807
rect 56523 15757 56579 15769
rect 56523 15751 56525 15757
rect 56525 15751 56577 15757
rect 56577 15751 56579 15757
rect 56523 15705 56525 15727
rect 56525 15705 56577 15727
rect 56577 15705 56579 15727
rect 56523 15693 56579 15705
rect 56523 15671 56525 15693
rect 56525 15671 56577 15693
rect 56577 15671 56579 15693
rect 56523 15641 56525 15647
rect 56525 15641 56577 15647
rect 56577 15641 56579 15647
rect 56523 15629 56579 15641
rect 56523 15591 56525 15629
rect 56525 15591 56577 15629
rect 56577 15591 56579 15629
rect 56523 15565 56579 15567
rect 56523 15513 56525 15565
rect 56525 15513 56577 15565
rect 56577 15513 56579 15565
rect 56523 15511 56579 15513
rect 56523 15449 56525 15487
rect 56525 15449 56577 15487
rect 56577 15449 56579 15487
rect 56523 15437 56579 15449
rect 56523 15431 56525 15437
rect 56525 15431 56577 15437
rect 56577 15431 56579 15437
rect 56523 15385 56525 15407
rect 56525 15385 56577 15407
rect 56577 15385 56579 15407
rect 56523 15373 56579 15385
rect 56523 15351 56525 15373
rect 56525 15351 56577 15373
rect 56577 15351 56579 15373
rect 56523 15321 56525 15327
rect 56525 15321 56577 15327
rect 56577 15321 56579 15327
rect 56523 15309 56579 15321
rect 56523 15271 56525 15309
rect 56525 15271 56577 15309
rect 56577 15271 56579 15309
rect 56523 15245 56579 15247
rect 56523 15193 56525 15245
rect 56525 15193 56577 15245
rect 56577 15193 56579 15245
rect 56523 15191 56579 15193
rect 56523 15129 56525 15167
rect 56525 15129 56577 15167
rect 56577 15129 56579 15167
rect 56523 15117 56579 15129
rect 56523 15111 56525 15117
rect 56525 15111 56577 15117
rect 56577 15111 56579 15117
rect 56523 15065 56525 15087
rect 56525 15065 56577 15087
rect 56577 15065 56579 15087
rect 56523 15053 56579 15065
rect 56523 15031 56525 15053
rect 56525 15031 56577 15053
rect 56577 15031 56579 15053
rect 56523 15001 56525 15007
rect 56525 15001 56577 15007
rect 56577 15001 56579 15007
rect 56523 14989 56579 15001
rect 56523 14951 56525 14989
rect 56525 14951 56577 14989
rect 56577 14951 56579 14989
rect 56523 14925 56579 14927
rect 56523 14873 56525 14925
rect 56525 14873 56577 14925
rect 56577 14873 56579 14925
rect 56523 14871 56579 14873
rect 56523 14809 56525 14847
rect 56525 14809 56577 14847
rect 56577 14809 56579 14847
rect 56523 14797 56579 14809
rect 56523 14791 56525 14797
rect 56525 14791 56577 14797
rect 56577 14791 56579 14797
rect 56523 14745 56525 14767
rect 56525 14745 56577 14767
rect 56577 14745 56579 14767
rect 56523 14733 56579 14745
rect 56523 14711 56525 14733
rect 56525 14711 56577 14733
rect 56577 14711 56579 14733
rect 56523 14681 56525 14687
rect 56525 14681 56577 14687
rect 56577 14681 56579 14687
rect 56523 14669 56579 14681
rect 56523 14631 56525 14669
rect 56525 14631 56577 14669
rect 56577 14631 56579 14669
rect 56523 14605 56579 14607
rect 56523 14553 56525 14605
rect 56525 14553 56577 14605
rect 56577 14553 56579 14605
rect 56523 14551 56579 14553
rect 56523 14489 56525 14527
rect 56525 14489 56577 14527
rect 56577 14489 56579 14527
rect 56523 14477 56579 14489
rect 56523 14471 56525 14477
rect 56525 14471 56577 14477
rect 56577 14471 56579 14477
rect 56523 14425 56525 14447
rect 56525 14425 56577 14447
rect 56577 14425 56579 14447
rect 56523 14413 56579 14425
rect 56523 14391 56525 14413
rect 56525 14391 56577 14413
rect 56577 14391 56579 14413
rect 56523 14361 56525 14367
rect 56525 14361 56577 14367
rect 56577 14361 56579 14367
rect 56523 14349 56579 14361
rect 56523 14311 56525 14349
rect 56525 14311 56577 14349
rect 56577 14311 56579 14349
rect 56523 14285 56579 14287
rect 56523 14233 56525 14285
rect 56525 14233 56577 14285
rect 56577 14233 56579 14285
rect 56523 14231 56579 14233
rect 56523 14169 56525 14207
rect 56525 14169 56577 14207
rect 56577 14169 56579 14207
rect 56523 14157 56579 14169
rect 56523 14151 56525 14157
rect 56525 14151 56577 14157
rect 56577 14151 56579 14157
rect 56523 14105 56525 14127
rect 56525 14105 56577 14127
rect 56577 14105 56579 14127
rect 56523 14093 56579 14105
rect 56523 14071 56525 14093
rect 56525 14071 56577 14093
rect 56577 14071 56579 14093
rect 56523 14041 56525 14047
rect 56525 14041 56577 14047
rect 56577 14041 56579 14047
rect 56523 14029 56579 14041
rect 56523 13991 56525 14029
rect 56525 13991 56577 14029
rect 56577 13991 56579 14029
rect 56523 13965 56579 13967
rect 56523 13913 56525 13965
rect 56525 13913 56577 13965
rect 56577 13913 56579 13965
rect 56523 13911 56579 13913
rect 54925 11912 55141 11930
rect 54925 11732 54943 11912
rect 54943 11732 55123 11912
rect 55123 11732 55141 11912
rect 54925 11714 55141 11732
<< metal3 >>
rect 40081 109629 40317 114463
rect 40081 109393 41920 109629
rect 41684 102167 41920 109393
rect 68084 109601 68320 114463
rect 80009 109774 80245 114463
rect 68084 109365 69937 109601
rect 80009 109538 81986 109774
rect 41674 102152 41930 102167
rect 41674 101936 41694 102152
rect 41910 101936 41930 102152
rect 69701 102138 69937 109365
rect 81750 102139 81986 109538
rect 41674 101921 41930 101936
rect 69690 102123 69946 102138
rect 69690 101907 69710 102123
rect 69926 101907 69946 102123
rect 69690 101892 69946 101907
rect 81740 102124 81996 102139
rect 81740 101908 81760 102124
rect 81976 101908 81996 102124
rect 81740 101893 81996 101908
rect 71228 100765 71376 100772
rect 40235 100714 40356 100750
rect 40235 100650 40263 100714
rect 40327 100650 40356 100714
rect 40235 100634 40356 100650
rect 40235 100570 40263 100634
rect 40327 100570 40356 100634
rect 40235 100554 40356 100570
rect 40235 100490 40263 100554
rect 40327 100490 40356 100554
rect 40235 100474 40356 100490
rect 40235 100410 40263 100474
rect 40327 100410 40356 100474
rect 40235 100394 40356 100410
rect 40235 100330 40263 100394
rect 40327 100330 40356 100394
rect 40235 100314 40356 100330
rect 40235 100250 40263 100314
rect 40327 100250 40356 100314
rect 40235 100234 40356 100250
rect 40235 100170 40263 100234
rect 40327 100170 40356 100234
rect 40235 100154 40356 100170
rect 40235 100090 40263 100154
rect 40327 100090 40356 100154
rect 40235 100074 40356 100090
rect 40235 100010 40263 100074
rect 40327 100010 40356 100074
rect 40235 99994 40356 100010
rect 40235 99930 40263 99994
rect 40327 99930 40356 99994
rect 40235 99914 40356 99930
rect 40235 99850 40263 99914
rect 40327 99850 40356 99914
rect 40235 99834 40356 99850
rect 40235 99770 40263 99834
rect 40327 99770 40356 99834
rect 40235 99754 40356 99770
rect 40235 99690 40263 99754
rect 40327 99690 40356 99754
rect 40235 99674 40356 99690
rect 40235 99610 40263 99674
rect 40327 99610 40356 99674
rect 40235 99594 40356 99610
rect 40235 99530 40263 99594
rect 40327 99530 40356 99594
rect 40235 99514 40356 99530
rect 40235 99450 40263 99514
rect 40327 99450 40356 99514
rect 40235 99434 40356 99450
rect 40235 99370 40263 99434
rect 40327 99370 40356 99434
rect 40235 99354 40356 99370
rect 40235 99290 40263 99354
rect 40327 99290 40356 99354
rect 40235 99274 40356 99290
rect 40235 99210 40263 99274
rect 40327 99210 40356 99274
rect 40235 99194 40356 99210
rect 40235 99130 40263 99194
rect 40327 99130 40356 99194
rect 40235 99114 40356 99130
rect 40235 99050 40263 99114
rect 40327 99050 40356 99114
rect 40235 99034 40356 99050
rect 40235 98970 40263 99034
rect 40327 98970 40356 99034
rect 40235 98954 40356 98970
rect 40235 98890 40263 98954
rect 40327 98890 40356 98954
rect 40235 98874 40356 98890
rect 40235 98810 40263 98874
rect 40327 98810 40356 98874
rect 40235 98794 40356 98810
rect 40235 98730 40263 98794
rect 40327 98730 40356 98794
rect 40235 98714 40356 98730
rect 40235 98650 40263 98714
rect 40327 98650 40356 98714
rect 40235 98634 40356 98650
rect 40235 98570 40263 98634
rect 40327 98570 40356 98634
rect 40235 98554 40356 98570
rect 40235 98490 40263 98554
rect 40327 98490 40356 98554
rect 40235 98474 40356 98490
rect 40235 98410 40263 98474
rect 40327 98410 40356 98474
rect 40235 98394 40356 98410
rect 40235 98330 40263 98394
rect 40327 98330 40356 98394
rect 40235 98314 40356 98330
rect 40235 98250 40263 98314
rect 40327 98250 40356 98314
rect 40235 98234 40356 98250
rect 40235 98170 40263 98234
rect 40327 98170 40356 98234
rect 40235 98154 40356 98170
rect 40235 98090 40263 98154
rect 40327 98090 40356 98154
rect 40235 98074 40356 98090
rect 40235 98010 40263 98074
rect 40327 98010 40356 98074
rect 40235 97994 40356 98010
rect 40235 97930 40263 97994
rect 40327 97930 40356 97994
rect 40235 97914 40356 97930
rect 40235 97850 40263 97914
rect 40327 97850 40356 97914
rect 40235 97834 40356 97850
rect 40235 97770 40263 97834
rect 40327 97770 40356 97834
rect 40235 97754 40356 97770
rect 40235 97690 40263 97754
rect 40327 97690 40356 97754
rect 40235 97674 40356 97690
rect 40235 97610 40263 97674
rect 40327 97610 40356 97674
rect 40235 97594 40356 97610
rect 40235 97530 40263 97594
rect 40327 97530 40356 97594
rect 40235 97514 40356 97530
rect 40235 97450 40263 97514
rect 40327 97450 40356 97514
rect 40235 97415 40356 97450
rect 43236 100720 43357 100756
rect 43236 100656 43264 100720
rect 43328 100656 43357 100720
rect 43236 100640 43357 100656
rect 43236 100576 43264 100640
rect 43328 100576 43357 100640
rect 43236 100560 43357 100576
rect 43236 100496 43264 100560
rect 43328 100496 43357 100560
rect 43236 100480 43357 100496
rect 43236 100416 43264 100480
rect 43328 100416 43357 100480
rect 43236 100400 43357 100416
rect 43236 100336 43264 100400
rect 43328 100336 43357 100400
rect 43236 100320 43357 100336
rect 43236 100256 43264 100320
rect 43328 100256 43357 100320
rect 43236 100240 43357 100256
rect 43236 100176 43264 100240
rect 43328 100176 43357 100240
rect 43236 100160 43357 100176
rect 43236 100096 43264 100160
rect 43328 100096 43357 100160
rect 43236 100080 43357 100096
rect 43236 100016 43264 100080
rect 43328 100016 43357 100080
rect 43236 100000 43357 100016
rect 43236 99936 43264 100000
rect 43328 99936 43357 100000
rect 43236 99920 43357 99936
rect 43236 99856 43264 99920
rect 43328 99856 43357 99920
rect 43236 99840 43357 99856
rect 43236 99776 43264 99840
rect 43328 99776 43357 99840
rect 43236 99760 43357 99776
rect 43236 99696 43264 99760
rect 43328 99696 43357 99760
rect 43236 99680 43357 99696
rect 43236 99616 43264 99680
rect 43328 99616 43357 99680
rect 43236 99600 43357 99616
rect 43236 99536 43264 99600
rect 43328 99536 43357 99600
rect 43236 99520 43357 99536
rect 43236 99456 43264 99520
rect 43328 99456 43357 99520
rect 43236 99440 43357 99456
rect 43236 99376 43264 99440
rect 43328 99376 43357 99440
rect 43236 99360 43357 99376
rect 43236 99296 43264 99360
rect 43328 99296 43357 99360
rect 43236 99280 43357 99296
rect 43236 99216 43264 99280
rect 43328 99216 43357 99280
rect 43236 99200 43357 99216
rect 43236 99136 43264 99200
rect 43328 99136 43357 99200
rect 43236 99120 43357 99136
rect 43236 99056 43264 99120
rect 43328 99056 43357 99120
rect 43236 99040 43357 99056
rect 43236 98976 43264 99040
rect 43328 98976 43357 99040
rect 43236 98960 43357 98976
rect 43236 98896 43264 98960
rect 43328 98896 43357 98960
rect 43236 98880 43357 98896
rect 43236 98816 43264 98880
rect 43328 98816 43357 98880
rect 43236 98800 43357 98816
rect 43236 98736 43264 98800
rect 43328 98736 43357 98800
rect 43236 98720 43357 98736
rect 43236 98656 43264 98720
rect 43328 98656 43357 98720
rect 43236 98640 43357 98656
rect 43236 98576 43264 98640
rect 43328 98576 43357 98640
rect 43236 98560 43357 98576
rect 43236 98496 43264 98560
rect 43328 98496 43357 98560
rect 43236 98480 43357 98496
rect 43236 98416 43264 98480
rect 43328 98416 43357 98480
rect 43236 98400 43357 98416
rect 43236 98336 43264 98400
rect 43328 98336 43357 98400
rect 43236 98320 43357 98336
rect 43236 98256 43264 98320
rect 43328 98256 43357 98320
rect 43236 98240 43357 98256
rect 43236 98176 43264 98240
rect 43328 98176 43357 98240
rect 43236 98160 43357 98176
rect 43236 98096 43264 98160
rect 43328 98096 43357 98160
rect 43236 98080 43357 98096
rect 43236 98016 43264 98080
rect 43328 98016 43357 98080
rect 43236 98000 43357 98016
rect 43236 97936 43264 98000
rect 43328 97936 43357 98000
rect 43236 97920 43357 97936
rect 43236 97856 43264 97920
rect 43328 97856 43357 97920
rect 43236 97840 43357 97856
rect 43236 97776 43264 97840
rect 43328 97776 43357 97840
rect 43236 97760 43357 97776
rect 43236 97696 43264 97760
rect 43328 97696 43357 97760
rect 43236 97680 43357 97696
rect 43236 97616 43264 97680
rect 43328 97616 43357 97680
rect 43236 97600 43357 97616
rect 43236 97536 43264 97600
rect 43328 97536 43357 97600
rect 43236 97520 43357 97536
rect 43236 97456 43264 97520
rect 43328 97456 43357 97520
rect 43236 97421 43357 97456
rect 68227 100752 68375 100759
rect 68227 100716 68273 100752
rect 68329 100716 68375 100752
rect 68227 100652 68269 100716
rect 68333 100652 68375 100716
rect 68227 100636 68273 100652
rect 68329 100636 68375 100652
rect 68227 100572 68269 100636
rect 68333 100572 68375 100636
rect 68227 100556 68273 100572
rect 68329 100556 68375 100572
rect 68227 100492 68269 100556
rect 68333 100492 68375 100556
rect 68227 100476 68273 100492
rect 68329 100476 68375 100492
rect 68227 100412 68269 100476
rect 68333 100412 68375 100476
rect 68227 100396 68273 100412
rect 68329 100396 68375 100412
rect 68227 100332 68269 100396
rect 68333 100332 68375 100396
rect 68227 100316 68273 100332
rect 68329 100316 68375 100332
rect 68227 100252 68269 100316
rect 68333 100252 68375 100316
rect 68227 100236 68273 100252
rect 68329 100236 68375 100252
rect 68227 100172 68269 100236
rect 68333 100172 68375 100236
rect 68227 100156 68273 100172
rect 68329 100156 68375 100172
rect 68227 100092 68269 100156
rect 68333 100092 68375 100156
rect 68227 100076 68273 100092
rect 68329 100076 68375 100092
rect 68227 100012 68269 100076
rect 68333 100012 68375 100076
rect 68227 99996 68273 100012
rect 68329 99996 68375 100012
rect 68227 99932 68269 99996
rect 68333 99932 68375 99996
rect 68227 99916 68273 99932
rect 68329 99916 68375 99932
rect 68227 99852 68269 99916
rect 68333 99852 68375 99916
rect 68227 99836 68273 99852
rect 68329 99836 68375 99852
rect 68227 99772 68269 99836
rect 68333 99772 68375 99836
rect 68227 99756 68273 99772
rect 68329 99756 68375 99772
rect 68227 99692 68269 99756
rect 68333 99692 68375 99756
rect 68227 99676 68273 99692
rect 68329 99676 68375 99692
rect 68227 99612 68269 99676
rect 68333 99612 68375 99676
rect 68227 99596 68273 99612
rect 68329 99596 68375 99612
rect 68227 99532 68269 99596
rect 68333 99532 68375 99596
rect 68227 99516 68273 99532
rect 68329 99516 68375 99532
rect 68227 99452 68269 99516
rect 68333 99452 68375 99516
rect 68227 99436 68273 99452
rect 68329 99436 68375 99452
rect 68227 99372 68269 99436
rect 68333 99372 68375 99436
rect 68227 99356 68273 99372
rect 68329 99356 68375 99372
rect 68227 99292 68269 99356
rect 68333 99292 68375 99356
rect 68227 99276 68273 99292
rect 68329 99276 68375 99292
rect 68227 99212 68269 99276
rect 68333 99212 68375 99276
rect 68227 99196 68273 99212
rect 68329 99196 68375 99212
rect 68227 99132 68269 99196
rect 68333 99132 68375 99196
rect 68227 99116 68273 99132
rect 68329 99116 68375 99132
rect 68227 99052 68269 99116
rect 68333 99052 68375 99116
rect 68227 99036 68273 99052
rect 68329 99036 68375 99052
rect 68227 98972 68269 99036
rect 68333 98972 68375 99036
rect 68227 98956 68273 98972
rect 68329 98956 68375 98972
rect 68227 98892 68269 98956
rect 68333 98892 68375 98956
rect 68227 98876 68273 98892
rect 68329 98876 68375 98892
rect 68227 98812 68269 98876
rect 68333 98812 68375 98876
rect 68227 98796 68273 98812
rect 68329 98796 68375 98812
rect 68227 98732 68269 98796
rect 68333 98732 68375 98796
rect 68227 98716 68273 98732
rect 68329 98716 68375 98732
rect 68227 98652 68269 98716
rect 68333 98652 68375 98716
rect 68227 98636 68273 98652
rect 68329 98636 68375 98652
rect 68227 98572 68269 98636
rect 68333 98572 68375 98636
rect 68227 98556 68273 98572
rect 68329 98556 68375 98572
rect 68227 98492 68269 98556
rect 68333 98492 68375 98556
rect 68227 98476 68273 98492
rect 68329 98476 68375 98492
rect 68227 98412 68269 98476
rect 68333 98412 68375 98476
rect 68227 98396 68273 98412
rect 68329 98396 68375 98412
rect 68227 98332 68269 98396
rect 68333 98332 68375 98396
rect 68227 98316 68273 98332
rect 68329 98316 68375 98332
rect 68227 98252 68269 98316
rect 68333 98252 68375 98316
rect 68227 98236 68273 98252
rect 68329 98236 68375 98252
rect 68227 98172 68269 98236
rect 68333 98172 68375 98236
rect 68227 98156 68273 98172
rect 68329 98156 68375 98172
rect 68227 98092 68269 98156
rect 68333 98092 68375 98156
rect 68227 98076 68273 98092
rect 68329 98076 68375 98092
rect 68227 98012 68269 98076
rect 68333 98012 68375 98076
rect 68227 97996 68273 98012
rect 68329 97996 68375 98012
rect 68227 97932 68269 97996
rect 68333 97932 68375 97996
rect 68227 97916 68273 97932
rect 68329 97916 68375 97932
rect 68227 97852 68269 97916
rect 68333 97852 68375 97916
rect 68227 97836 68273 97852
rect 68329 97836 68375 97852
rect 68227 97772 68269 97836
rect 68333 97772 68375 97836
rect 68227 97756 68273 97772
rect 68329 97756 68375 97772
rect 68227 97692 68269 97756
rect 68333 97692 68375 97756
rect 68227 97676 68273 97692
rect 68329 97676 68375 97692
rect 68227 97612 68269 97676
rect 68333 97612 68375 97676
rect 68227 97596 68273 97612
rect 68329 97596 68375 97612
rect 68227 97532 68269 97596
rect 68333 97532 68375 97596
rect 68227 97516 68273 97532
rect 68329 97516 68375 97532
rect 68227 97452 68269 97516
rect 68333 97452 68375 97516
rect 68227 97416 68273 97452
rect 68329 97416 68375 97452
rect 71228 100729 71274 100765
rect 71330 100729 71376 100765
rect 71228 100665 71270 100729
rect 71334 100665 71376 100729
rect 71228 100649 71274 100665
rect 71330 100649 71376 100665
rect 71228 100585 71270 100649
rect 71334 100585 71376 100649
rect 71228 100569 71274 100585
rect 71330 100569 71376 100585
rect 71228 100505 71270 100569
rect 71334 100505 71376 100569
rect 71228 100489 71274 100505
rect 71330 100489 71376 100505
rect 71228 100425 71270 100489
rect 71334 100425 71376 100489
rect 71228 100409 71274 100425
rect 71330 100409 71376 100425
rect 71228 100345 71270 100409
rect 71334 100345 71376 100409
rect 71228 100329 71274 100345
rect 71330 100329 71376 100345
rect 71228 100265 71270 100329
rect 71334 100265 71376 100329
rect 71228 100249 71274 100265
rect 71330 100249 71376 100265
rect 71228 100185 71270 100249
rect 71334 100185 71376 100249
rect 71228 100169 71274 100185
rect 71330 100169 71376 100185
rect 71228 100105 71270 100169
rect 71334 100105 71376 100169
rect 71228 100089 71274 100105
rect 71330 100089 71376 100105
rect 71228 100025 71270 100089
rect 71334 100025 71376 100089
rect 71228 100009 71274 100025
rect 71330 100009 71376 100025
rect 71228 99945 71270 100009
rect 71334 99945 71376 100009
rect 71228 99929 71274 99945
rect 71330 99929 71376 99945
rect 71228 99865 71270 99929
rect 71334 99865 71376 99929
rect 71228 99849 71274 99865
rect 71330 99849 71376 99865
rect 71228 99785 71270 99849
rect 71334 99785 71376 99849
rect 71228 99769 71274 99785
rect 71330 99769 71376 99785
rect 71228 99705 71270 99769
rect 71334 99705 71376 99769
rect 71228 99689 71274 99705
rect 71330 99689 71376 99705
rect 71228 99625 71270 99689
rect 71334 99625 71376 99689
rect 71228 99609 71274 99625
rect 71330 99609 71376 99625
rect 71228 99545 71270 99609
rect 71334 99545 71376 99609
rect 71228 99529 71274 99545
rect 71330 99529 71376 99545
rect 71228 99465 71270 99529
rect 71334 99465 71376 99529
rect 71228 99449 71274 99465
rect 71330 99449 71376 99465
rect 71228 99385 71270 99449
rect 71334 99385 71376 99449
rect 71228 99369 71274 99385
rect 71330 99369 71376 99385
rect 71228 99305 71270 99369
rect 71334 99305 71376 99369
rect 71228 99289 71274 99305
rect 71330 99289 71376 99305
rect 71228 99225 71270 99289
rect 71334 99225 71376 99289
rect 71228 99209 71274 99225
rect 71330 99209 71376 99225
rect 71228 99145 71270 99209
rect 71334 99145 71376 99209
rect 71228 99129 71274 99145
rect 71330 99129 71376 99145
rect 71228 99065 71270 99129
rect 71334 99065 71376 99129
rect 71228 99049 71274 99065
rect 71330 99049 71376 99065
rect 71228 98985 71270 99049
rect 71334 98985 71376 99049
rect 71228 98969 71274 98985
rect 71330 98969 71376 98985
rect 71228 98905 71270 98969
rect 71334 98905 71376 98969
rect 71228 98889 71274 98905
rect 71330 98889 71376 98905
rect 71228 98825 71270 98889
rect 71334 98825 71376 98889
rect 71228 98809 71274 98825
rect 71330 98809 71376 98825
rect 71228 98745 71270 98809
rect 71334 98745 71376 98809
rect 71228 98729 71274 98745
rect 71330 98729 71376 98745
rect 71228 98665 71270 98729
rect 71334 98665 71376 98729
rect 71228 98649 71274 98665
rect 71330 98649 71376 98665
rect 71228 98585 71270 98649
rect 71334 98585 71376 98649
rect 71228 98569 71274 98585
rect 71330 98569 71376 98585
rect 71228 98505 71270 98569
rect 71334 98505 71376 98569
rect 71228 98489 71274 98505
rect 71330 98489 71376 98505
rect 71228 98425 71270 98489
rect 71334 98425 71376 98489
rect 71228 98409 71274 98425
rect 71330 98409 71376 98425
rect 71228 98345 71270 98409
rect 71334 98345 71376 98409
rect 71228 98329 71274 98345
rect 71330 98329 71376 98345
rect 71228 98265 71270 98329
rect 71334 98265 71376 98329
rect 71228 98249 71274 98265
rect 71330 98249 71376 98265
rect 71228 98185 71270 98249
rect 71334 98185 71376 98249
rect 71228 98169 71274 98185
rect 71330 98169 71376 98185
rect 71228 98105 71270 98169
rect 71334 98105 71376 98169
rect 71228 98089 71274 98105
rect 71330 98089 71376 98105
rect 71228 98025 71270 98089
rect 71334 98025 71376 98089
rect 71228 98009 71274 98025
rect 71330 98009 71376 98025
rect 71228 97945 71270 98009
rect 71334 97945 71376 98009
rect 71228 97929 71274 97945
rect 71330 97929 71376 97945
rect 71228 97865 71270 97929
rect 71334 97865 71376 97929
rect 71228 97849 71274 97865
rect 71330 97849 71376 97865
rect 71228 97785 71270 97849
rect 71334 97785 71376 97849
rect 71228 97769 71274 97785
rect 71330 97769 71376 97785
rect 71228 97705 71270 97769
rect 71334 97705 71376 97769
rect 71228 97689 71274 97705
rect 71330 97689 71376 97705
rect 71228 97625 71270 97689
rect 71334 97625 71376 97689
rect 71228 97609 71274 97625
rect 71330 97609 71376 97625
rect 71228 97545 71270 97609
rect 71334 97545 71376 97609
rect 71228 97529 71274 97545
rect 71330 97529 71376 97545
rect 71228 97465 71270 97529
rect 71334 97465 71376 97529
rect 71228 97429 71274 97465
rect 71330 97429 71376 97465
rect 71228 97422 71376 97429
rect 114815 99997 120001 100233
rect 68227 97409 68375 97416
rect 40397 95824 40534 95854
rect 40397 95760 40430 95824
rect 40494 95760 40534 95824
rect 40397 95728 40534 95760
rect 41585 95820 41702 95842
rect 41585 95756 41608 95820
rect 41672 95756 41702 95820
rect 41585 95731 41702 95756
rect 41802 95827 41918 95857
rect 41802 95763 41825 95827
rect 41889 95763 41918 95827
rect 41802 95736 41918 95763
rect 42933 95824 43053 95848
rect 42933 95760 42959 95824
rect 43023 95760 43053 95824
rect 42933 95731 43053 95760
rect 40517 94320 40625 94341
rect 40517 94256 40540 94320
rect 40604 94256 40625 94320
rect 40517 94228 40625 94256
rect 41630 94306 41739 94326
rect 41630 94242 41654 94306
rect 41718 94242 41739 94306
rect 41630 94219 41739 94242
rect 41845 94307 41954 94332
rect 41845 94243 41867 94307
rect 41931 94243 41954 94307
rect 41845 94219 41954 94243
rect 43003 94307 43140 94333
rect 43003 94243 43031 94307
rect 43095 94243 43140 94307
rect 43003 94219 43140 94243
rect 114815 93442 115051 99997
rect 93649 93356 115051 93442
rect 93649 93292 93725 93356
rect 93789 93292 115051 93356
rect 93649 93206 115051 93292
rect 43131 92763 120001 92835
rect 40376 92725 40460 92730
rect 43131 92725 93160 92763
rect 40376 92721 93160 92725
rect 40376 92665 40390 92721
rect 40446 92699 93160 92721
rect 93224 92699 120001 92763
rect 40446 92665 120001 92699
rect 40376 92661 120001 92665
rect 40376 92656 40460 92661
rect 43131 92599 120001 92661
rect 41662 92514 41746 92542
rect 41662 92450 41672 92514
rect 41736 92450 41746 92514
rect 41662 92434 41746 92450
rect 41662 92370 41672 92434
rect 41736 92370 41746 92434
rect 41662 92354 41746 92370
rect 41662 92290 41672 92354
rect 41736 92290 41746 92354
rect 41121 92277 41214 92288
rect 41121 92213 41135 92277
rect 41199 92213 41214 92277
rect 41121 92197 41214 92213
rect 41121 92133 41135 92197
rect 41199 92133 41214 92197
rect 41662 92274 41746 92290
rect 41662 92210 41672 92274
rect 41736 92210 41746 92274
rect 41662 92183 41746 92210
rect 42205 92280 42298 92291
rect 42205 92216 42219 92280
rect 42283 92216 42298 92280
rect 42205 92200 42298 92216
rect 41121 92122 41214 92133
rect 42205 92136 42219 92200
rect 42283 92136 42298 92200
rect 42205 92125 42298 92136
rect 43128 92103 115126 92191
rect 42885 92095 42969 92100
rect 43128 92095 92571 92103
rect 42885 92091 92571 92095
rect 42885 92035 42899 92091
rect 42955 92039 92571 92091
rect 92635 92039 115126 92103
rect 42955 92035 115126 92039
rect 42885 92031 115126 92035
rect 42885 92026 42969 92031
rect 43128 91955 115126 92031
rect 40489 91635 40612 91665
rect 40489 91571 40517 91635
rect 40581 91571 40612 91635
rect 40489 91540 40612 91571
rect 41645 91629 41764 91655
rect 41645 91565 41672 91629
rect 41736 91565 41764 91629
rect 41645 91535 41764 91565
rect 42766 91640 42883 91663
rect 42766 91576 42790 91640
rect 42854 91576 42883 91640
rect 42766 91548 42883 91576
rect 43988 90727 43998 90791
rect 44062 90727 49021 90791
rect 49085 90727 49095 90791
rect 44769 90404 44779 90468
rect 44843 90404 49828 90468
rect 49892 90404 49902 90468
rect 45781 89971 45789 90035
rect 45853 89971 54421 90035
rect 54485 89971 54495 90035
rect 46550 89718 46558 89782
rect 46622 89718 55228 89782
rect 55292 89718 55302 89782
rect 49011 89287 49021 89351
rect 49085 89287 49095 89351
rect 54411 89287 54421 89351
rect 54485 89287 54495 89351
rect 49818 89034 49828 89098
rect 49892 89034 49902 89098
rect 55218 89034 55228 89098
rect 55292 89034 55302 89098
rect 74514 88750 74600 88770
rect 74514 88686 74525 88750
rect 74589 88686 74600 88750
rect 74514 88670 74600 88686
rect 74514 88606 74525 88670
rect 74589 88606 74600 88670
rect 74514 88590 74600 88606
rect 74514 88526 74525 88590
rect 74589 88526 74600 88590
rect 74514 88510 74600 88526
rect 74514 88446 74525 88510
rect 74589 88446 74600 88510
rect 74514 88430 74600 88446
rect 74514 88366 74525 88430
rect 74589 88366 74600 88430
rect 74514 88350 74600 88366
rect 74514 88286 74525 88350
rect 74589 88286 74600 88350
rect 74514 88270 74600 88286
rect 74514 88206 74525 88270
rect 74589 88206 74600 88270
rect 74514 88186 74600 88206
rect 81042 88750 81128 88770
rect 81042 88686 81053 88750
rect 81117 88686 81128 88750
rect 81042 88670 81128 88686
rect 81042 88606 81053 88670
rect 81117 88606 81128 88670
rect 81042 88590 81128 88606
rect 81042 88526 81053 88590
rect 81117 88526 81128 88590
rect 81042 88510 81128 88526
rect 81042 88446 81053 88510
rect 81117 88446 81128 88510
rect 81042 88430 81128 88446
rect 81042 88366 81053 88430
rect 81117 88366 81128 88430
rect 81042 88350 81128 88366
rect 81042 88286 81053 88350
rect 81117 88286 81128 88350
rect 81042 88270 81128 88286
rect 81042 88206 81053 88270
rect 81117 88206 81128 88270
rect 81042 88186 81128 88206
rect 88658 88750 88744 88770
rect 88658 88686 88669 88750
rect 88733 88686 88744 88750
rect 88658 88670 88744 88686
rect 88658 88606 88669 88670
rect 88733 88606 88744 88670
rect 88658 88590 88744 88606
rect 88658 88526 88669 88590
rect 88733 88526 88744 88590
rect 88658 88510 88744 88526
rect 88658 88446 88669 88510
rect 88733 88446 88744 88510
rect 88658 88430 88744 88446
rect 88658 88366 88669 88430
rect 88733 88366 88744 88430
rect 88658 88350 88744 88366
rect 88658 88286 88669 88350
rect 88733 88286 88744 88350
rect 88658 88270 88744 88286
rect 88658 88206 88669 88270
rect 88733 88206 88744 88270
rect 88658 88186 88744 88206
rect 46013 87555 46367 87579
rect 46013 87251 46038 87555
rect 46342 87424 46367 87555
rect 47200 87424 47662 87429
rect 46342 87360 46907 87424
rect 46971 87360 46981 87424
rect 47200 87360 47239 87424
rect 47303 87360 47319 87424
rect 47383 87360 47399 87424
rect 47463 87360 47479 87424
rect 47543 87360 47559 87424
rect 47623 87360 47662 87424
rect 46342 87251 46367 87360
rect 47200 87355 47662 87360
rect 49011 87426 49473 87431
rect 49011 87362 49050 87426
rect 49114 87362 49130 87426
rect 49194 87362 49210 87426
rect 49274 87362 49290 87426
rect 49354 87362 49370 87426
rect 49434 87362 49473 87426
rect 49011 87357 49473 87362
rect 50806 87422 51268 87427
rect 50806 87358 50845 87422
rect 50909 87358 50925 87422
rect 50989 87358 51005 87422
rect 51069 87358 51085 87422
rect 51149 87358 51165 87422
rect 51229 87358 51268 87422
rect 50806 87353 51268 87358
rect 52605 87420 53067 87425
rect 52605 87356 52644 87420
rect 52708 87356 52724 87420
rect 52788 87356 52804 87420
rect 52868 87356 52884 87420
rect 52948 87356 52964 87420
rect 53028 87356 53067 87420
rect 52605 87351 53067 87356
rect 54396 87424 54858 87429
rect 54396 87360 54435 87424
rect 54499 87360 54515 87424
rect 54579 87360 54595 87424
rect 54659 87360 54675 87424
rect 54739 87360 54755 87424
rect 54819 87360 54858 87424
rect 54396 87355 54858 87360
rect 56198 87420 56660 87425
rect 56198 87356 56237 87420
rect 56301 87356 56317 87420
rect 56381 87356 56397 87420
rect 56461 87356 56477 87420
rect 56541 87356 56557 87420
rect 56621 87356 56660 87420
rect 56198 87351 56660 87356
rect 46013 87227 46367 87251
rect 57841 87246 58391 87259
rect 50145 87220 50405 87233
rect 50145 86996 50163 87220
rect 50387 86996 50405 87220
rect 57841 87022 57884 87246
rect 58348 87022 58391 87246
rect 57841 87009 58391 87022
rect 50145 86983 50405 86996
rect 75059 86747 75145 86767
rect 75059 86683 75070 86747
rect 75134 86683 75145 86747
rect 75059 86667 75145 86683
rect 75059 86603 75070 86667
rect 75134 86603 75145 86667
rect 75059 86587 75145 86603
rect 75059 86523 75070 86587
rect 75134 86523 75145 86587
rect 75059 86507 75145 86523
rect 75059 86443 75070 86507
rect 75134 86443 75145 86507
rect 75059 86427 75145 86443
rect 75059 86363 75070 86427
rect 75134 86363 75145 86427
rect 75059 86347 75145 86363
rect 75059 86283 75070 86347
rect 75134 86283 75145 86347
rect 75059 86267 75145 86283
rect 75059 86203 75070 86267
rect 75134 86203 75145 86267
rect 75059 86183 75145 86203
rect 76147 86747 76233 86767
rect 76147 86683 76158 86747
rect 76222 86683 76233 86747
rect 76147 86667 76233 86683
rect 76147 86603 76158 86667
rect 76222 86603 76233 86667
rect 76147 86587 76233 86603
rect 76147 86523 76158 86587
rect 76222 86523 76233 86587
rect 76147 86507 76233 86523
rect 76147 86443 76158 86507
rect 76222 86443 76233 86507
rect 76147 86427 76233 86443
rect 76147 86363 76158 86427
rect 76222 86363 76233 86427
rect 76147 86347 76233 86363
rect 76147 86283 76158 86347
rect 76222 86283 76233 86347
rect 76147 86267 76233 86283
rect 76147 86203 76158 86267
rect 76222 86203 76233 86267
rect 76147 86183 76233 86203
rect 78323 86747 78409 86767
rect 78323 86683 78334 86747
rect 78398 86683 78409 86747
rect 78323 86667 78409 86683
rect 78323 86603 78334 86667
rect 78398 86603 78409 86667
rect 78323 86587 78409 86603
rect 78323 86523 78334 86587
rect 78398 86523 78409 86587
rect 78323 86507 78409 86523
rect 78323 86443 78334 86507
rect 78398 86443 78409 86507
rect 78323 86427 78409 86443
rect 78323 86363 78334 86427
rect 78398 86363 78409 86427
rect 78323 86347 78409 86363
rect 78323 86283 78334 86347
rect 78398 86283 78409 86347
rect 78323 86267 78409 86283
rect 78323 86203 78334 86267
rect 78398 86203 78409 86267
rect 78323 86183 78409 86203
rect 79411 86747 79497 86767
rect 79411 86683 79422 86747
rect 79486 86683 79497 86747
rect 79411 86667 79497 86683
rect 79411 86603 79422 86667
rect 79486 86603 79497 86667
rect 79411 86587 79497 86603
rect 79411 86523 79422 86587
rect 79486 86523 79497 86587
rect 79411 86507 79497 86523
rect 79411 86443 79422 86507
rect 79486 86443 79497 86507
rect 79411 86427 79497 86443
rect 79411 86363 79422 86427
rect 79486 86363 79497 86427
rect 79411 86347 79497 86363
rect 79411 86283 79422 86347
rect 79486 86283 79497 86347
rect 79411 86267 79497 86283
rect 79411 86203 79422 86267
rect 79486 86203 79497 86267
rect 79411 86183 79497 86203
rect 80499 86747 80585 86767
rect 80499 86683 80510 86747
rect 80574 86683 80585 86747
rect 80499 86667 80585 86683
rect 80499 86603 80510 86667
rect 80574 86603 80585 86667
rect 80499 86587 80585 86603
rect 80499 86523 80510 86587
rect 80574 86523 80585 86587
rect 80499 86507 80585 86523
rect 80499 86443 80510 86507
rect 80574 86443 80585 86507
rect 80499 86427 80585 86443
rect 80499 86363 80510 86427
rect 80574 86363 80585 86427
rect 80499 86347 80585 86363
rect 80499 86283 80510 86347
rect 80574 86283 80585 86347
rect 80499 86267 80585 86283
rect 80499 86203 80510 86267
rect 80574 86203 80585 86267
rect 80499 86183 80585 86203
rect 81587 86747 81673 86767
rect 81587 86683 81598 86747
rect 81662 86683 81673 86747
rect 81587 86667 81673 86683
rect 81587 86603 81598 86667
rect 81662 86603 81673 86667
rect 81587 86587 81673 86603
rect 81587 86523 81598 86587
rect 81662 86523 81673 86587
rect 81587 86507 81673 86523
rect 81587 86443 81598 86507
rect 81662 86443 81673 86507
rect 81587 86427 81673 86443
rect 81587 86363 81598 86427
rect 81662 86363 81673 86427
rect 81587 86347 81673 86363
rect 81587 86283 81598 86347
rect 81662 86283 81673 86347
rect 81587 86267 81673 86283
rect 81587 86203 81598 86267
rect 81662 86203 81673 86267
rect 81587 86183 81673 86203
rect 82675 86747 82761 86767
rect 82675 86683 82686 86747
rect 82750 86683 82761 86747
rect 82675 86667 82761 86683
rect 82675 86603 82686 86667
rect 82750 86603 82761 86667
rect 82675 86587 82761 86603
rect 82675 86523 82686 86587
rect 82750 86523 82761 86587
rect 82675 86507 82761 86523
rect 82675 86443 82686 86507
rect 82750 86443 82761 86507
rect 82675 86427 82761 86443
rect 82675 86363 82686 86427
rect 82750 86363 82761 86427
rect 82675 86347 82761 86363
rect 82675 86283 82686 86347
rect 82750 86283 82761 86347
rect 82675 86267 82761 86283
rect 82675 86203 82686 86267
rect 82750 86203 82761 86267
rect 82675 86183 82761 86203
rect 83763 86747 83849 86767
rect 83763 86683 83774 86747
rect 83838 86683 83849 86747
rect 83763 86667 83849 86683
rect 83763 86603 83774 86667
rect 83838 86603 83849 86667
rect 83763 86587 83849 86603
rect 83763 86523 83774 86587
rect 83838 86523 83849 86587
rect 83763 86507 83849 86523
rect 83763 86443 83774 86507
rect 83838 86443 83849 86507
rect 83763 86427 83849 86443
rect 83763 86363 83774 86427
rect 83838 86363 83849 86427
rect 83763 86347 83849 86363
rect 83763 86283 83774 86347
rect 83838 86283 83849 86347
rect 83763 86267 83849 86283
rect 83763 86203 83774 86267
rect 83838 86203 83849 86267
rect 83763 86183 83849 86203
rect 85939 86747 86025 86767
rect 85939 86683 85950 86747
rect 86014 86683 86025 86747
rect 85939 86667 86025 86683
rect 85939 86603 85950 86667
rect 86014 86603 86025 86667
rect 85939 86587 86025 86603
rect 85939 86523 85950 86587
rect 86014 86523 86025 86587
rect 85939 86507 86025 86523
rect 85939 86443 85950 86507
rect 86014 86443 86025 86507
rect 85939 86427 86025 86443
rect 85939 86363 85950 86427
rect 86014 86363 86025 86427
rect 85939 86347 86025 86363
rect 85939 86283 85950 86347
rect 86014 86283 86025 86347
rect 85939 86267 86025 86283
rect 85939 86203 85950 86267
rect 86014 86203 86025 86267
rect 85939 86183 86025 86203
rect 87027 86747 87113 86767
rect 87027 86683 87038 86747
rect 87102 86683 87113 86747
rect 87027 86667 87113 86683
rect 87027 86603 87038 86667
rect 87102 86603 87113 86667
rect 87027 86587 87113 86603
rect 87027 86523 87038 86587
rect 87102 86523 87113 86587
rect 87027 86507 87113 86523
rect 87027 86443 87038 86507
rect 87102 86443 87113 86507
rect 87027 86427 87113 86443
rect 87027 86363 87038 86427
rect 87102 86363 87113 86427
rect 87027 86347 87113 86363
rect 87027 86283 87038 86347
rect 87102 86283 87113 86347
rect 87027 86267 87113 86283
rect 87027 86203 87038 86267
rect 87102 86203 87113 86267
rect 87027 86183 87113 86203
rect 88115 86747 88201 86767
rect 88115 86683 88126 86747
rect 88190 86683 88201 86747
rect 88115 86667 88201 86683
rect 88115 86603 88126 86667
rect 88190 86603 88201 86667
rect 88115 86587 88201 86603
rect 88115 86523 88126 86587
rect 88190 86523 88201 86587
rect 88115 86507 88201 86523
rect 88115 86443 88126 86507
rect 88190 86443 88201 86507
rect 88115 86427 88201 86443
rect 88115 86363 88126 86427
rect 88190 86363 88201 86427
rect 88115 86347 88201 86363
rect 88115 86283 88126 86347
rect 88190 86283 88201 86347
rect 88115 86267 88201 86283
rect 88115 86203 88126 86267
rect 88190 86203 88201 86267
rect 88115 86183 88201 86203
rect 114890 85397 115126 91955
rect 114890 85161 120001 85397
rect 57431 84828 57623 84854
rect 48511 78617 48623 78641
rect 48511 78553 48537 78617
rect 48601 78553 48623 78617
rect 48511 78529 48623 78553
rect 50205 78618 50322 78647
rect 50205 78554 50228 78618
rect 50292 78554 50322 78618
rect 50205 78530 50322 78554
rect 51915 78617 52012 78636
rect 51915 78553 51933 78617
rect 51997 78553 52012 78617
rect 51915 78533 52012 78553
rect 53709 78617 53814 78644
rect 53709 78553 53729 78617
rect 53793 78553 53814 78617
rect 53709 78534 53814 78553
rect 55538 78617 55641 78637
rect 55538 78553 55558 78617
rect 55622 78553 55641 78617
rect 55538 78533 55641 78553
rect 47380 78425 47642 78430
rect 47380 78361 47399 78425
rect 47463 78361 47479 78425
rect 47543 78361 47559 78425
rect 47623 78361 47642 78425
rect 47380 78356 47642 78361
rect 49175 78424 49437 78429
rect 49175 78360 49194 78424
rect 49258 78360 49274 78424
rect 49338 78360 49354 78424
rect 49418 78360 49437 78424
rect 49175 78355 49437 78360
rect 50975 78426 51237 78431
rect 50975 78362 50994 78426
rect 51058 78362 51074 78426
rect 51138 78362 51154 78426
rect 51218 78362 51237 78426
rect 50975 78357 51237 78362
rect 52773 78425 53035 78430
rect 52773 78361 52792 78425
rect 52856 78361 52872 78425
rect 52936 78361 52952 78425
rect 53016 78361 53035 78425
rect 52773 78356 53035 78361
rect 54571 78426 54833 78431
rect 54571 78362 54590 78426
rect 54654 78362 54670 78426
rect 54734 78362 54750 78426
rect 54814 78362 54833 78426
rect 54571 78357 54833 78362
rect 56374 78425 56636 78430
rect 56374 78361 56393 78425
rect 56457 78361 56473 78425
rect 56537 78361 56553 78425
rect 56617 78361 56636 78425
rect 56374 78356 56636 78361
rect 57250 78426 57352 78446
rect 57250 78362 57270 78426
rect 57334 78362 57352 78426
rect 57250 78341 57352 78362
rect 49819 78041 49829 78105
rect 49893 78041 49903 78105
rect 55219 78041 55229 78105
rect 55293 78041 55303 78105
rect 49011 77788 49021 77852
rect 49085 77788 49095 77852
rect 54411 77788 54421 77852
rect 54485 77788 54495 77852
rect 46548 77360 46558 77424
rect 46622 77360 55229 77424
rect 55293 77360 55303 77424
rect 45779 77104 45789 77168
rect 45853 77104 54421 77168
rect 54485 77104 54495 77168
rect 57431 77164 57455 84828
rect 57599 77164 57623 84828
rect 57431 77138 57623 77164
rect 67261 84840 67655 84863
rect 44769 76671 44779 76735
rect 44843 76671 49829 76735
rect 49893 76671 49903 76735
rect 43988 76348 43998 76412
rect 44062 76348 49021 76412
rect 49085 76348 49095 76412
rect 48230 75265 48334 75276
rect 48230 75201 48250 75265
rect 48314 75201 48334 75265
rect 48230 75185 48334 75201
rect 48230 75121 48250 75185
rect 48314 75121 48334 75185
rect 49352 75269 49460 75294
rect 49352 75205 49372 75269
rect 49436 75205 49460 75269
rect 49352 75184 49460 75205
rect 48230 75105 48334 75121
rect 48230 75041 48250 75105
rect 48314 75041 48334 75105
rect 48230 75031 48334 75041
rect 51396 75068 53216 75093
rect 51396 74924 51434 75068
rect 53178 74924 53216 75068
rect 51396 74900 53216 74924
rect 53722 75079 54568 75101
rect 53722 74935 53753 75079
rect 54537 74935 54568 75079
rect 53722 74913 54568 74935
rect 55429 75069 56339 75091
rect 55429 74925 55452 75069
rect 56316 74925 56339 75069
rect 55429 74903 56339 74925
rect 48210 74798 48324 74818
rect 48210 74734 48235 74798
rect 48299 74734 48324 74798
rect 57006 74793 57225 74801
rect 57006 74757 57047 74793
rect 57183 74757 57225 74793
rect 48210 74718 48324 74734
rect 48210 74654 48235 74718
rect 48299 74654 48324 74718
rect 48210 74639 48324 74654
rect 37992 74638 48324 74639
rect 37992 74618 48235 74638
rect 37992 74554 38089 74618
rect 38153 74574 48235 74618
rect 48299 74574 48324 74638
rect 38153 74558 48324 74574
rect 38153 74554 48235 74558
rect 37992 74534 48235 74554
rect 48210 74494 48235 74534
rect 48299 74494 48324 74558
rect 48210 74478 48324 74494
rect 51152 74742 51356 74747
rect 48210 74414 48235 74478
rect 48299 74414 48324 74478
rect 48210 74395 48324 74414
rect 48597 74463 48696 74483
rect 48597 74399 48614 74463
rect 48678 74399 48696 74463
rect 48597 74379 48696 74399
rect 0 74094 29094 74177
rect 0 74030 48614 74094
rect 48678 74030 48688 74094
rect 0 73941 29094 74030
rect 30014 73742 30378 73747
rect 30014 73678 30044 73742
rect 30108 73678 30124 73742
rect 30188 73678 30204 73742
rect 30268 73678 30284 73742
rect 30348 73678 30378 73742
rect 30014 73673 30378 73678
rect 30622 73440 30686 74030
rect 31024 73446 31108 73451
rect 31024 73442 49372 73446
rect 30622 73431 30947 73440
rect 30622 73375 30703 73431
rect 30759 73375 30783 73431
rect 30839 73375 30863 73431
rect 30919 73375 30947 73431
rect 31024 73386 31038 73442
rect 31094 73386 49372 73442
rect 31024 73382 49372 73386
rect 49436 73382 49446 73446
rect 31024 73377 31108 73382
rect 30622 73371 30947 73375
rect 30676 73366 30947 73371
rect 31100 73200 31464 73205
rect 31100 73136 31130 73200
rect 31194 73136 31210 73200
rect 31274 73136 31290 73200
rect 31354 73136 31370 73200
rect 31434 73136 31464 73200
rect 31100 73131 31464 73136
rect 51152 71798 51182 74742
rect 51326 71798 51356 74742
rect 51152 71793 51356 71798
rect 57006 71813 57043 74757
rect 57187 71813 57225 74757
rect 57006 71777 57047 71813
rect 57183 71777 57225 71813
rect 57006 71769 57225 71777
rect 67261 71656 67306 84840
rect 67610 71656 67655 84840
rect 74514 84750 74600 84770
rect 74514 84686 74525 84750
rect 74589 84686 74600 84750
rect 74514 84670 74600 84686
rect 74514 84606 74525 84670
rect 74589 84606 74600 84670
rect 74514 84590 74600 84606
rect 74514 84526 74525 84590
rect 74589 84526 74600 84590
rect 74514 84510 74600 84526
rect 74514 84446 74525 84510
rect 74589 84446 74600 84510
rect 74514 84430 74600 84446
rect 74514 84366 74525 84430
rect 74589 84366 74600 84430
rect 74514 84350 74600 84366
rect 74514 84286 74525 84350
rect 74589 84286 74600 84350
rect 74514 84270 74600 84286
rect 74514 84206 74525 84270
rect 74589 84206 74600 84270
rect 74514 84186 74600 84206
rect 75602 84750 75688 84770
rect 75602 84686 75613 84750
rect 75677 84686 75688 84750
rect 75602 84670 75688 84686
rect 75602 84606 75613 84670
rect 75677 84606 75688 84670
rect 75602 84590 75688 84606
rect 75602 84526 75613 84590
rect 75677 84526 75688 84590
rect 75602 84510 75688 84526
rect 75602 84446 75613 84510
rect 75677 84446 75688 84510
rect 75602 84430 75688 84446
rect 75602 84366 75613 84430
rect 75677 84366 75688 84430
rect 75602 84350 75688 84366
rect 75602 84286 75613 84350
rect 75677 84286 75688 84350
rect 75602 84270 75688 84286
rect 75602 84206 75613 84270
rect 75677 84206 75688 84270
rect 75602 84186 75688 84206
rect 76690 84750 76776 84770
rect 76690 84686 76701 84750
rect 76765 84686 76776 84750
rect 76690 84670 76776 84686
rect 76690 84606 76701 84670
rect 76765 84606 76776 84670
rect 76690 84590 76776 84606
rect 76690 84526 76701 84590
rect 76765 84526 76776 84590
rect 76690 84510 76776 84526
rect 76690 84446 76701 84510
rect 76765 84446 76776 84510
rect 76690 84430 76776 84446
rect 76690 84366 76701 84430
rect 76765 84366 76776 84430
rect 76690 84350 76776 84366
rect 76690 84286 76701 84350
rect 76765 84286 76776 84350
rect 76690 84270 76776 84286
rect 76690 84206 76701 84270
rect 76765 84206 76776 84270
rect 76690 84186 76776 84206
rect 77778 84750 77864 84770
rect 77778 84686 77789 84750
rect 77853 84686 77864 84750
rect 77778 84670 77864 84686
rect 77778 84606 77789 84670
rect 77853 84606 77864 84670
rect 77778 84590 77864 84606
rect 77778 84526 77789 84590
rect 77853 84526 77864 84590
rect 77778 84510 77864 84526
rect 77778 84446 77789 84510
rect 77853 84446 77864 84510
rect 77778 84430 77864 84446
rect 77778 84366 77789 84430
rect 77853 84366 77864 84430
rect 77778 84350 77864 84366
rect 77778 84286 77789 84350
rect 77853 84286 77864 84350
rect 77778 84270 77864 84286
rect 77778 84206 77789 84270
rect 77853 84206 77864 84270
rect 77778 84186 77864 84206
rect 78866 84750 78952 84770
rect 78866 84686 78877 84750
rect 78941 84686 78952 84750
rect 78866 84670 78952 84686
rect 78866 84606 78877 84670
rect 78941 84606 78952 84670
rect 78866 84590 78952 84606
rect 78866 84526 78877 84590
rect 78941 84526 78952 84590
rect 78866 84510 78952 84526
rect 78866 84446 78877 84510
rect 78941 84446 78952 84510
rect 78866 84430 78952 84446
rect 78866 84366 78877 84430
rect 78941 84366 78952 84430
rect 78866 84350 78952 84366
rect 78866 84286 78877 84350
rect 78941 84286 78952 84350
rect 78866 84270 78952 84286
rect 78866 84206 78877 84270
rect 78941 84206 78952 84270
rect 78866 84186 78952 84206
rect 79954 84750 80040 84770
rect 79954 84686 79965 84750
rect 80029 84686 80040 84750
rect 79954 84670 80040 84686
rect 79954 84606 79965 84670
rect 80029 84606 80040 84670
rect 79954 84590 80040 84606
rect 79954 84526 79965 84590
rect 80029 84526 80040 84590
rect 79954 84510 80040 84526
rect 79954 84446 79965 84510
rect 80029 84446 80040 84510
rect 79954 84430 80040 84446
rect 79954 84366 79965 84430
rect 80029 84366 80040 84430
rect 79954 84350 80040 84366
rect 79954 84286 79965 84350
rect 80029 84286 80040 84350
rect 79954 84270 80040 84286
rect 79954 84206 79965 84270
rect 80029 84206 80040 84270
rect 79954 84186 80040 84206
rect 81042 84750 81128 84770
rect 81042 84686 81053 84750
rect 81117 84686 81128 84750
rect 81042 84670 81128 84686
rect 81042 84606 81053 84670
rect 81117 84606 81128 84670
rect 81042 84590 81128 84606
rect 81042 84526 81053 84590
rect 81117 84526 81128 84590
rect 81042 84510 81128 84526
rect 81042 84446 81053 84510
rect 81117 84446 81128 84510
rect 81042 84430 81128 84446
rect 81042 84366 81053 84430
rect 81117 84366 81128 84430
rect 81042 84350 81128 84366
rect 81042 84286 81053 84350
rect 81117 84286 81128 84350
rect 81042 84270 81128 84286
rect 81042 84206 81053 84270
rect 81117 84206 81128 84270
rect 81042 84186 81128 84206
rect 82130 84750 82216 84770
rect 82130 84686 82141 84750
rect 82205 84686 82216 84750
rect 82130 84670 82216 84686
rect 82130 84606 82141 84670
rect 82205 84606 82216 84670
rect 82130 84590 82216 84606
rect 82130 84526 82141 84590
rect 82205 84526 82216 84590
rect 82130 84510 82216 84526
rect 82130 84446 82141 84510
rect 82205 84446 82216 84510
rect 82130 84430 82216 84446
rect 82130 84366 82141 84430
rect 82205 84366 82216 84430
rect 82130 84350 82216 84366
rect 82130 84286 82141 84350
rect 82205 84286 82216 84350
rect 82130 84270 82216 84286
rect 82130 84206 82141 84270
rect 82205 84206 82216 84270
rect 82130 84186 82216 84206
rect 83218 84750 83304 84770
rect 83218 84686 83229 84750
rect 83293 84686 83304 84750
rect 83218 84670 83304 84686
rect 83218 84606 83229 84670
rect 83293 84606 83304 84670
rect 83218 84590 83304 84606
rect 83218 84526 83229 84590
rect 83293 84526 83304 84590
rect 83218 84510 83304 84526
rect 83218 84446 83229 84510
rect 83293 84446 83304 84510
rect 83218 84430 83304 84446
rect 83218 84366 83229 84430
rect 83293 84366 83304 84430
rect 83218 84350 83304 84366
rect 83218 84286 83229 84350
rect 83293 84286 83304 84350
rect 83218 84270 83304 84286
rect 83218 84206 83229 84270
rect 83293 84206 83304 84270
rect 83218 84186 83304 84206
rect 84306 84750 84392 84770
rect 84306 84686 84317 84750
rect 84381 84686 84392 84750
rect 84306 84670 84392 84686
rect 84306 84606 84317 84670
rect 84381 84606 84392 84670
rect 84306 84590 84392 84606
rect 84306 84526 84317 84590
rect 84381 84526 84392 84590
rect 84306 84510 84392 84526
rect 84306 84446 84317 84510
rect 84381 84446 84392 84510
rect 84306 84430 84392 84446
rect 84306 84366 84317 84430
rect 84381 84366 84392 84430
rect 84306 84350 84392 84366
rect 84306 84286 84317 84350
rect 84381 84286 84392 84350
rect 84306 84270 84392 84286
rect 84306 84206 84317 84270
rect 84381 84206 84392 84270
rect 84306 84186 84392 84206
rect 85394 84750 85480 84770
rect 85394 84686 85405 84750
rect 85469 84686 85480 84750
rect 85394 84670 85480 84686
rect 85394 84606 85405 84670
rect 85469 84606 85480 84670
rect 85394 84590 85480 84606
rect 85394 84526 85405 84590
rect 85469 84526 85480 84590
rect 85394 84510 85480 84526
rect 85394 84446 85405 84510
rect 85469 84446 85480 84510
rect 85394 84430 85480 84446
rect 85394 84366 85405 84430
rect 85469 84366 85480 84430
rect 85394 84350 85480 84366
rect 85394 84286 85405 84350
rect 85469 84286 85480 84350
rect 85394 84270 85480 84286
rect 85394 84206 85405 84270
rect 85469 84206 85480 84270
rect 85394 84186 85480 84206
rect 86482 84750 86568 84770
rect 86482 84686 86493 84750
rect 86557 84686 86568 84750
rect 86482 84670 86568 84686
rect 86482 84606 86493 84670
rect 86557 84606 86568 84670
rect 86482 84590 86568 84606
rect 86482 84526 86493 84590
rect 86557 84526 86568 84590
rect 86482 84510 86568 84526
rect 86482 84446 86493 84510
rect 86557 84446 86568 84510
rect 86482 84430 86568 84446
rect 86482 84366 86493 84430
rect 86557 84366 86568 84430
rect 86482 84350 86568 84366
rect 86482 84286 86493 84350
rect 86557 84286 86568 84350
rect 86482 84270 86568 84286
rect 86482 84206 86493 84270
rect 86557 84206 86568 84270
rect 86482 84186 86568 84206
rect 87570 84750 87656 84770
rect 87570 84686 87581 84750
rect 87645 84686 87656 84750
rect 87570 84670 87656 84686
rect 87570 84606 87581 84670
rect 87645 84606 87656 84670
rect 87570 84590 87656 84606
rect 87570 84526 87581 84590
rect 87645 84526 87656 84590
rect 87570 84510 87656 84526
rect 87570 84446 87581 84510
rect 87645 84446 87656 84510
rect 87570 84430 87656 84446
rect 87570 84366 87581 84430
rect 87645 84366 87656 84430
rect 87570 84350 87656 84366
rect 87570 84286 87581 84350
rect 87645 84286 87656 84350
rect 87570 84270 87656 84286
rect 87570 84206 87581 84270
rect 87645 84206 87656 84270
rect 87570 84186 87656 84206
rect 88658 84750 88744 84770
rect 88658 84686 88669 84750
rect 88733 84686 88744 84750
rect 88658 84670 88744 84686
rect 88658 84606 88669 84670
rect 88733 84606 88744 84670
rect 88658 84590 88744 84606
rect 88658 84526 88669 84590
rect 88733 84526 88744 84590
rect 88658 84510 88744 84526
rect 88658 84446 88669 84510
rect 88733 84446 88744 84510
rect 88658 84430 88744 84446
rect 88658 84366 88669 84430
rect 88733 84366 88744 84430
rect 88658 84350 88744 84366
rect 88658 84286 88669 84350
rect 88733 84286 88744 84350
rect 88658 84270 88744 84286
rect 88658 84206 88669 84270
rect 88733 84206 88744 84270
rect 88658 84186 88744 84206
rect 75059 82747 75145 82767
rect 75059 82683 75070 82747
rect 75134 82683 75145 82747
rect 75059 82667 75145 82683
rect 75059 82603 75070 82667
rect 75134 82603 75145 82667
rect 75059 82587 75145 82603
rect 75059 82523 75070 82587
rect 75134 82523 75145 82587
rect 75059 82507 75145 82523
rect 75059 82443 75070 82507
rect 75134 82443 75145 82507
rect 75059 82427 75145 82443
rect 75059 82363 75070 82427
rect 75134 82363 75145 82427
rect 75059 82347 75145 82363
rect 75059 82283 75070 82347
rect 75134 82283 75145 82347
rect 75059 82267 75145 82283
rect 75059 82203 75070 82267
rect 75134 82203 75145 82267
rect 75059 82183 75145 82203
rect 76147 82747 76233 82767
rect 76147 82683 76158 82747
rect 76222 82683 76233 82747
rect 76147 82667 76233 82683
rect 76147 82603 76158 82667
rect 76222 82603 76233 82667
rect 76147 82587 76233 82603
rect 76147 82523 76158 82587
rect 76222 82523 76233 82587
rect 76147 82507 76233 82523
rect 76147 82443 76158 82507
rect 76222 82443 76233 82507
rect 76147 82427 76233 82443
rect 76147 82363 76158 82427
rect 76222 82363 76233 82427
rect 76147 82347 76233 82363
rect 76147 82283 76158 82347
rect 76222 82283 76233 82347
rect 76147 82267 76233 82283
rect 76147 82203 76158 82267
rect 76222 82203 76233 82267
rect 76147 82183 76233 82203
rect 77235 82747 77321 82767
rect 77235 82683 77246 82747
rect 77310 82683 77321 82747
rect 77235 82667 77321 82683
rect 77235 82603 77246 82667
rect 77310 82603 77321 82667
rect 77235 82587 77321 82603
rect 77235 82523 77246 82587
rect 77310 82523 77321 82587
rect 77235 82507 77321 82523
rect 77235 82443 77246 82507
rect 77310 82443 77321 82507
rect 77235 82427 77321 82443
rect 77235 82363 77246 82427
rect 77310 82363 77321 82427
rect 77235 82347 77321 82363
rect 77235 82283 77246 82347
rect 77310 82283 77321 82347
rect 77235 82267 77321 82283
rect 77235 82203 77246 82267
rect 77310 82203 77321 82267
rect 77235 82183 77321 82203
rect 78323 82747 78409 82767
rect 78323 82683 78334 82747
rect 78398 82683 78409 82747
rect 78323 82667 78409 82683
rect 78323 82603 78334 82667
rect 78398 82603 78409 82667
rect 78323 82587 78409 82603
rect 78323 82523 78334 82587
rect 78398 82523 78409 82587
rect 78323 82507 78409 82523
rect 78323 82443 78334 82507
rect 78398 82443 78409 82507
rect 78323 82427 78409 82443
rect 78323 82363 78334 82427
rect 78398 82363 78409 82427
rect 78323 82347 78409 82363
rect 78323 82283 78334 82347
rect 78398 82283 78409 82347
rect 78323 82267 78409 82283
rect 78323 82203 78334 82267
rect 78398 82203 78409 82267
rect 78323 82183 78409 82203
rect 79411 82747 79497 82767
rect 79411 82683 79422 82747
rect 79486 82683 79497 82747
rect 79411 82667 79497 82683
rect 79411 82603 79422 82667
rect 79486 82603 79497 82667
rect 79411 82587 79497 82603
rect 79411 82523 79422 82587
rect 79486 82523 79497 82587
rect 79411 82507 79497 82523
rect 79411 82443 79422 82507
rect 79486 82443 79497 82507
rect 79411 82427 79497 82443
rect 79411 82363 79422 82427
rect 79486 82363 79497 82427
rect 79411 82347 79497 82363
rect 79411 82283 79422 82347
rect 79486 82283 79497 82347
rect 79411 82267 79497 82283
rect 79411 82203 79422 82267
rect 79486 82203 79497 82267
rect 79411 82183 79497 82203
rect 80499 82747 80585 82767
rect 80499 82683 80510 82747
rect 80574 82683 80585 82747
rect 80499 82667 80585 82683
rect 80499 82603 80510 82667
rect 80574 82603 80585 82667
rect 80499 82587 80585 82603
rect 80499 82523 80510 82587
rect 80574 82523 80585 82587
rect 80499 82507 80585 82523
rect 80499 82443 80510 82507
rect 80574 82443 80585 82507
rect 80499 82427 80585 82443
rect 80499 82363 80510 82427
rect 80574 82363 80585 82427
rect 80499 82347 80585 82363
rect 80499 82283 80510 82347
rect 80574 82283 80585 82347
rect 80499 82267 80585 82283
rect 80499 82203 80510 82267
rect 80574 82203 80585 82267
rect 80499 82183 80585 82203
rect 81587 82747 81673 82767
rect 81587 82683 81598 82747
rect 81662 82683 81673 82747
rect 81587 82667 81673 82683
rect 81587 82603 81598 82667
rect 81662 82603 81673 82667
rect 81587 82587 81673 82603
rect 81587 82523 81598 82587
rect 81662 82523 81673 82587
rect 81587 82507 81673 82523
rect 81587 82443 81598 82507
rect 81662 82443 81673 82507
rect 81587 82427 81673 82443
rect 81587 82363 81598 82427
rect 81662 82363 81673 82427
rect 81587 82347 81673 82363
rect 81587 82283 81598 82347
rect 81662 82283 81673 82347
rect 81587 82267 81673 82283
rect 81587 82203 81598 82267
rect 81662 82203 81673 82267
rect 81587 82183 81673 82203
rect 82675 82747 82761 82767
rect 82675 82683 82686 82747
rect 82750 82683 82761 82747
rect 82675 82667 82761 82683
rect 82675 82603 82686 82667
rect 82750 82603 82761 82667
rect 82675 82587 82761 82603
rect 82675 82523 82686 82587
rect 82750 82523 82761 82587
rect 82675 82507 82761 82523
rect 82675 82443 82686 82507
rect 82750 82443 82761 82507
rect 82675 82427 82761 82443
rect 82675 82363 82686 82427
rect 82750 82363 82761 82427
rect 82675 82347 82761 82363
rect 82675 82283 82686 82347
rect 82750 82283 82761 82347
rect 82675 82267 82761 82283
rect 82675 82203 82686 82267
rect 82750 82203 82761 82267
rect 82675 82183 82761 82203
rect 83763 82747 83849 82767
rect 83763 82683 83774 82747
rect 83838 82683 83849 82747
rect 83763 82667 83849 82683
rect 83763 82603 83774 82667
rect 83838 82603 83849 82667
rect 83763 82587 83849 82603
rect 83763 82523 83774 82587
rect 83838 82523 83849 82587
rect 83763 82507 83849 82523
rect 83763 82443 83774 82507
rect 83838 82443 83849 82507
rect 83763 82427 83849 82443
rect 83763 82363 83774 82427
rect 83838 82363 83849 82427
rect 83763 82347 83849 82363
rect 83763 82283 83774 82347
rect 83838 82283 83849 82347
rect 83763 82267 83849 82283
rect 83763 82203 83774 82267
rect 83838 82203 83849 82267
rect 83763 82183 83849 82203
rect 84851 82747 84937 82767
rect 84851 82683 84862 82747
rect 84926 82683 84937 82747
rect 84851 82667 84937 82683
rect 84851 82603 84862 82667
rect 84926 82603 84937 82667
rect 84851 82587 84937 82603
rect 84851 82523 84862 82587
rect 84926 82523 84937 82587
rect 84851 82507 84937 82523
rect 84851 82443 84862 82507
rect 84926 82443 84937 82507
rect 84851 82427 84937 82443
rect 84851 82363 84862 82427
rect 84926 82363 84937 82427
rect 84851 82347 84937 82363
rect 84851 82283 84862 82347
rect 84926 82283 84937 82347
rect 84851 82267 84937 82283
rect 84851 82203 84862 82267
rect 84926 82203 84937 82267
rect 84851 82183 84937 82203
rect 85939 82747 86025 82767
rect 85939 82683 85950 82747
rect 86014 82683 86025 82747
rect 85939 82667 86025 82683
rect 85939 82603 85950 82667
rect 86014 82603 86025 82667
rect 85939 82587 86025 82603
rect 85939 82523 85950 82587
rect 86014 82523 86025 82587
rect 85939 82507 86025 82523
rect 85939 82443 85950 82507
rect 86014 82443 86025 82507
rect 85939 82427 86025 82443
rect 85939 82363 85950 82427
rect 86014 82363 86025 82427
rect 85939 82347 86025 82363
rect 85939 82283 85950 82347
rect 86014 82283 86025 82347
rect 85939 82267 86025 82283
rect 85939 82203 85950 82267
rect 86014 82203 86025 82267
rect 85939 82183 86025 82203
rect 87027 82747 87113 82767
rect 87027 82683 87038 82747
rect 87102 82683 87113 82747
rect 87027 82667 87113 82683
rect 87027 82603 87038 82667
rect 87102 82603 87113 82667
rect 87027 82587 87113 82603
rect 87027 82523 87038 82587
rect 87102 82523 87113 82587
rect 87027 82507 87113 82523
rect 87027 82443 87038 82507
rect 87102 82443 87113 82507
rect 87027 82427 87113 82443
rect 87027 82363 87038 82427
rect 87102 82363 87113 82427
rect 87027 82347 87113 82363
rect 87027 82283 87038 82347
rect 87102 82283 87113 82347
rect 87027 82267 87113 82283
rect 87027 82203 87038 82267
rect 87102 82203 87113 82267
rect 87027 82183 87113 82203
rect 88115 82747 88201 82767
rect 88115 82683 88126 82747
rect 88190 82683 88201 82747
rect 88115 82667 88201 82683
rect 88115 82603 88126 82667
rect 88190 82603 88201 82667
rect 88115 82587 88201 82603
rect 88115 82523 88126 82587
rect 88190 82523 88201 82587
rect 88115 82507 88201 82523
rect 88115 82443 88126 82507
rect 88190 82443 88201 82507
rect 88115 82427 88201 82443
rect 88115 82363 88126 82427
rect 88190 82363 88201 82427
rect 88115 82347 88201 82363
rect 88115 82283 88126 82347
rect 88190 82283 88201 82347
rect 88115 82267 88201 82283
rect 88115 82203 88126 82267
rect 88190 82203 88201 82267
rect 88115 82183 88201 82203
rect 74514 80750 74600 80770
rect 74514 80686 74525 80750
rect 74589 80686 74600 80750
rect 74514 80670 74600 80686
rect 74514 80606 74525 80670
rect 74589 80606 74600 80670
rect 74514 80590 74600 80606
rect 74514 80526 74525 80590
rect 74589 80526 74600 80590
rect 74514 80510 74600 80526
rect 74514 80446 74525 80510
rect 74589 80446 74600 80510
rect 74514 80430 74600 80446
rect 74514 80366 74525 80430
rect 74589 80366 74600 80430
rect 74514 80350 74600 80366
rect 74514 80286 74525 80350
rect 74589 80286 74600 80350
rect 74514 80270 74600 80286
rect 74514 80206 74525 80270
rect 74589 80206 74600 80270
rect 74514 80186 74600 80206
rect 75602 80750 75688 80770
rect 75602 80686 75613 80750
rect 75677 80686 75688 80750
rect 75602 80670 75688 80686
rect 75602 80606 75613 80670
rect 75677 80606 75688 80670
rect 75602 80590 75688 80606
rect 75602 80526 75613 80590
rect 75677 80526 75688 80590
rect 75602 80510 75688 80526
rect 75602 80446 75613 80510
rect 75677 80446 75688 80510
rect 75602 80430 75688 80446
rect 75602 80366 75613 80430
rect 75677 80366 75688 80430
rect 75602 80350 75688 80366
rect 75602 80286 75613 80350
rect 75677 80286 75688 80350
rect 75602 80270 75688 80286
rect 75602 80206 75613 80270
rect 75677 80206 75688 80270
rect 75602 80186 75688 80206
rect 76690 80750 76776 80770
rect 76690 80686 76701 80750
rect 76765 80686 76776 80750
rect 76690 80670 76776 80686
rect 76690 80606 76701 80670
rect 76765 80606 76776 80670
rect 76690 80590 76776 80606
rect 76690 80526 76701 80590
rect 76765 80526 76776 80590
rect 76690 80510 76776 80526
rect 76690 80446 76701 80510
rect 76765 80446 76776 80510
rect 76690 80430 76776 80446
rect 76690 80366 76701 80430
rect 76765 80366 76776 80430
rect 76690 80350 76776 80366
rect 76690 80286 76701 80350
rect 76765 80286 76776 80350
rect 76690 80270 76776 80286
rect 76690 80206 76701 80270
rect 76765 80206 76776 80270
rect 76690 80186 76776 80206
rect 77778 80750 77864 80770
rect 77778 80686 77789 80750
rect 77853 80686 77864 80750
rect 77778 80670 77864 80686
rect 77778 80606 77789 80670
rect 77853 80606 77864 80670
rect 77778 80590 77864 80606
rect 77778 80526 77789 80590
rect 77853 80526 77864 80590
rect 77778 80510 77864 80526
rect 77778 80446 77789 80510
rect 77853 80446 77864 80510
rect 77778 80430 77864 80446
rect 77778 80366 77789 80430
rect 77853 80366 77864 80430
rect 77778 80350 77864 80366
rect 77778 80286 77789 80350
rect 77853 80286 77864 80350
rect 77778 80270 77864 80286
rect 77778 80206 77789 80270
rect 77853 80206 77864 80270
rect 77778 80186 77864 80206
rect 78866 80750 78952 80770
rect 78866 80686 78877 80750
rect 78941 80686 78952 80750
rect 78866 80670 78952 80686
rect 78866 80606 78877 80670
rect 78941 80606 78952 80670
rect 78866 80590 78952 80606
rect 78866 80526 78877 80590
rect 78941 80526 78952 80590
rect 78866 80510 78952 80526
rect 78866 80446 78877 80510
rect 78941 80446 78952 80510
rect 78866 80430 78952 80446
rect 78866 80366 78877 80430
rect 78941 80366 78952 80430
rect 78866 80350 78952 80366
rect 78866 80286 78877 80350
rect 78941 80286 78952 80350
rect 78866 80270 78952 80286
rect 78866 80206 78877 80270
rect 78941 80206 78952 80270
rect 78866 80186 78952 80206
rect 79954 80750 80040 80770
rect 79954 80686 79965 80750
rect 80029 80686 80040 80750
rect 79954 80670 80040 80686
rect 79954 80606 79965 80670
rect 80029 80606 80040 80670
rect 79954 80590 80040 80606
rect 79954 80526 79965 80590
rect 80029 80526 80040 80590
rect 79954 80510 80040 80526
rect 79954 80446 79965 80510
rect 80029 80446 80040 80510
rect 79954 80430 80040 80446
rect 79954 80366 79965 80430
rect 80029 80366 80040 80430
rect 79954 80350 80040 80366
rect 79954 80286 79965 80350
rect 80029 80286 80040 80350
rect 79954 80270 80040 80286
rect 79954 80206 79965 80270
rect 80029 80206 80040 80270
rect 79954 80186 80040 80206
rect 81042 80750 81128 80770
rect 81042 80686 81053 80750
rect 81117 80686 81128 80750
rect 81042 80670 81128 80686
rect 81042 80606 81053 80670
rect 81117 80606 81128 80670
rect 81042 80590 81128 80606
rect 81042 80526 81053 80590
rect 81117 80526 81128 80590
rect 81042 80510 81128 80526
rect 81042 80446 81053 80510
rect 81117 80446 81128 80510
rect 81042 80430 81128 80446
rect 81042 80366 81053 80430
rect 81117 80366 81128 80430
rect 81042 80350 81128 80366
rect 81042 80286 81053 80350
rect 81117 80286 81128 80350
rect 81042 80270 81128 80286
rect 81042 80206 81053 80270
rect 81117 80206 81128 80270
rect 81042 80186 81128 80206
rect 82130 80750 82216 80770
rect 82130 80686 82141 80750
rect 82205 80686 82216 80750
rect 82130 80670 82216 80686
rect 82130 80606 82141 80670
rect 82205 80606 82216 80670
rect 82130 80590 82216 80606
rect 82130 80526 82141 80590
rect 82205 80526 82216 80590
rect 82130 80510 82216 80526
rect 82130 80446 82141 80510
rect 82205 80446 82216 80510
rect 82130 80430 82216 80446
rect 82130 80366 82141 80430
rect 82205 80366 82216 80430
rect 82130 80350 82216 80366
rect 82130 80286 82141 80350
rect 82205 80286 82216 80350
rect 82130 80270 82216 80286
rect 82130 80206 82141 80270
rect 82205 80206 82216 80270
rect 82130 80186 82216 80206
rect 83218 80750 83304 80770
rect 83218 80686 83229 80750
rect 83293 80686 83304 80750
rect 83218 80670 83304 80686
rect 83218 80606 83229 80670
rect 83293 80606 83304 80670
rect 83218 80590 83304 80606
rect 83218 80526 83229 80590
rect 83293 80526 83304 80590
rect 83218 80510 83304 80526
rect 83218 80446 83229 80510
rect 83293 80446 83304 80510
rect 83218 80430 83304 80446
rect 83218 80366 83229 80430
rect 83293 80366 83304 80430
rect 83218 80350 83304 80366
rect 83218 80286 83229 80350
rect 83293 80286 83304 80350
rect 83218 80270 83304 80286
rect 83218 80206 83229 80270
rect 83293 80206 83304 80270
rect 83218 80186 83304 80206
rect 84306 80750 84392 80770
rect 84306 80686 84317 80750
rect 84381 80686 84392 80750
rect 84306 80670 84392 80686
rect 84306 80606 84317 80670
rect 84381 80606 84392 80670
rect 84306 80590 84392 80606
rect 84306 80526 84317 80590
rect 84381 80526 84392 80590
rect 84306 80510 84392 80526
rect 84306 80446 84317 80510
rect 84381 80446 84392 80510
rect 84306 80430 84392 80446
rect 84306 80366 84317 80430
rect 84381 80366 84392 80430
rect 84306 80350 84392 80366
rect 84306 80286 84317 80350
rect 84381 80286 84392 80350
rect 84306 80270 84392 80286
rect 84306 80206 84317 80270
rect 84381 80206 84392 80270
rect 84306 80186 84392 80206
rect 85394 80750 85480 80770
rect 85394 80686 85405 80750
rect 85469 80686 85480 80750
rect 85394 80670 85480 80686
rect 85394 80606 85405 80670
rect 85469 80606 85480 80670
rect 85394 80590 85480 80606
rect 85394 80526 85405 80590
rect 85469 80526 85480 80590
rect 85394 80510 85480 80526
rect 85394 80446 85405 80510
rect 85469 80446 85480 80510
rect 85394 80430 85480 80446
rect 85394 80366 85405 80430
rect 85469 80366 85480 80430
rect 85394 80350 85480 80366
rect 85394 80286 85405 80350
rect 85469 80286 85480 80350
rect 85394 80270 85480 80286
rect 85394 80206 85405 80270
rect 85469 80206 85480 80270
rect 85394 80186 85480 80206
rect 86482 80750 86568 80770
rect 86482 80686 86493 80750
rect 86557 80686 86568 80750
rect 86482 80670 86568 80686
rect 86482 80606 86493 80670
rect 86557 80606 86568 80670
rect 86482 80590 86568 80606
rect 86482 80526 86493 80590
rect 86557 80526 86568 80590
rect 86482 80510 86568 80526
rect 86482 80446 86493 80510
rect 86557 80446 86568 80510
rect 86482 80430 86568 80446
rect 86482 80366 86493 80430
rect 86557 80366 86568 80430
rect 86482 80350 86568 80366
rect 86482 80286 86493 80350
rect 86557 80286 86568 80350
rect 86482 80270 86568 80286
rect 86482 80206 86493 80270
rect 86557 80206 86568 80270
rect 86482 80186 86568 80206
rect 87570 80750 87656 80770
rect 87570 80686 87581 80750
rect 87645 80686 87656 80750
rect 87570 80670 87656 80686
rect 87570 80606 87581 80670
rect 87645 80606 87656 80670
rect 87570 80590 87656 80606
rect 87570 80526 87581 80590
rect 87645 80526 87656 80590
rect 87570 80510 87656 80526
rect 87570 80446 87581 80510
rect 87645 80446 87656 80510
rect 87570 80430 87656 80446
rect 87570 80366 87581 80430
rect 87645 80366 87656 80430
rect 87570 80350 87656 80366
rect 87570 80286 87581 80350
rect 87645 80286 87656 80350
rect 87570 80270 87656 80286
rect 87570 80206 87581 80270
rect 87645 80206 87656 80270
rect 87570 80186 87656 80206
rect 88658 80750 88744 80770
rect 88658 80686 88669 80750
rect 88733 80686 88744 80750
rect 88658 80670 88744 80686
rect 88658 80606 88669 80670
rect 88733 80606 88744 80670
rect 88658 80590 88744 80606
rect 88658 80526 88669 80590
rect 88733 80526 88744 80590
rect 88658 80510 88744 80526
rect 88658 80446 88669 80510
rect 88733 80446 88744 80510
rect 88658 80430 88744 80446
rect 88658 80366 88669 80430
rect 88733 80366 88744 80430
rect 88658 80350 88744 80366
rect 88658 80286 88669 80350
rect 88733 80286 88744 80350
rect 88658 80270 88744 80286
rect 88658 80206 88669 80270
rect 88733 80206 88744 80270
rect 88658 80186 88744 80206
rect 109850 79123 120001 79359
rect 75059 78747 75145 78767
rect 75059 78683 75070 78747
rect 75134 78683 75145 78747
rect 75059 78667 75145 78683
rect 75059 78603 75070 78667
rect 75134 78603 75145 78667
rect 75059 78587 75145 78603
rect 75059 78523 75070 78587
rect 75134 78523 75145 78587
rect 75059 78507 75145 78523
rect 75059 78443 75070 78507
rect 75134 78443 75145 78507
rect 75059 78427 75145 78443
rect 75059 78363 75070 78427
rect 75134 78363 75145 78427
rect 75059 78347 75145 78363
rect 75059 78283 75070 78347
rect 75134 78283 75145 78347
rect 75059 78267 75145 78283
rect 75059 78203 75070 78267
rect 75134 78203 75145 78267
rect 75059 78183 75145 78203
rect 76147 78747 76233 78767
rect 76147 78683 76158 78747
rect 76222 78683 76233 78747
rect 76147 78667 76233 78683
rect 76147 78603 76158 78667
rect 76222 78603 76233 78667
rect 76147 78587 76233 78603
rect 76147 78523 76158 78587
rect 76222 78523 76233 78587
rect 76147 78507 76233 78523
rect 76147 78443 76158 78507
rect 76222 78443 76233 78507
rect 76147 78427 76233 78443
rect 76147 78363 76158 78427
rect 76222 78363 76233 78427
rect 76147 78347 76233 78363
rect 76147 78283 76158 78347
rect 76222 78283 76233 78347
rect 76147 78267 76233 78283
rect 76147 78203 76158 78267
rect 76222 78203 76233 78267
rect 76147 78183 76233 78203
rect 77235 78747 77321 78767
rect 77235 78683 77246 78747
rect 77310 78683 77321 78747
rect 77235 78667 77321 78683
rect 77235 78603 77246 78667
rect 77310 78603 77321 78667
rect 77235 78587 77321 78603
rect 77235 78523 77246 78587
rect 77310 78523 77321 78587
rect 77235 78507 77321 78523
rect 77235 78443 77246 78507
rect 77310 78443 77321 78507
rect 77235 78427 77321 78443
rect 77235 78363 77246 78427
rect 77310 78363 77321 78427
rect 77235 78347 77321 78363
rect 77235 78283 77246 78347
rect 77310 78283 77321 78347
rect 77235 78267 77321 78283
rect 77235 78203 77246 78267
rect 77310 78203 77321 78267
rect 77235 78183 77321 78203
rect 78323 78747 78409 78767
rect 78323 78683 78334 78747
rect 78398 78683 78409 78747
rect 78323 78667 78409 78683
rect 78323 78603 78334 78667
rect 78398 78603 78409 78667
rect 78323 78587 78409 78603
rect 78323 78523 78334 78587
rect 78398 78523 78409 78587
rect 78323 78507 78409 78523
rect 78323 78443 78334 78507
rect 78398 78443 78409 78507
rect 78323 78427 78409 78443
rect 78323 78363 78334 78427
rect 78398 78363 78409 78427
rect 78323 78347 78409 78363
rect 78323 78283 78334 78347
rect 78398 78283 78409 78347
rect 78323 78267 78409 78283
rect 78323 78203 78334 78267
rect 78398 78203 78409 78267
rect 78323 78183 78409 78203
rect 79411 78747 79497 78767
rect 79411 78683 79422 78747
rect 79486 78683 79497 78747
rect 79411 78667 79497 78683
rect 79411 78603 79422 78667
rect 79486 78603 79497 78667
rect 79411 78587 79497 78603
rect 79411 78523 79422 78587
rect 79486 78523 79497 78587
rect 79411 78507 79497 78523
rect 79411 78443 79422 78507
rect 79486 78443 79497 78507
rect 79411 78427 79497 78443
rect 79411 78363 79422 78427
rect 79486 78363 79497 78427
rect 79411 78347 79497 78363
rect 79411 78283 79422 78347
rect 79486 78283 79497 78347
rect 79411 78267 79497 78283
rect 79411 78203 79422 78267
rect 79486 78203 79497 78267
rect 79411 78183 79497 78203
rect 80499 78747 80585 78767
rect 80499 78683 80510 78747
rect 80574 78683 80585 78747
rect 80499 78667 80585 78683
rect 80499 78603 80510 78667
rect 80574 78603 80585 78667
rect 80499 78587 80585 78603
rect 80499 78523 80510 78587
rect 80574 78523 80585 78587
rect 80499 78507 80585 78523
rect 80499 78443 80510 78507
rect 80574 78443 80585 78507
rect 80499 78427 80585 78443
rect 80499 78363 80510 78427
rect 80574 78363 80585 78427
rect 80499 78347 80585 78363
rect 80499 78283 80510 78347
rect 80574 78283 80585 78347
rect 80499 78267 80585 78283
rect 80499 78203 80510 78267
rect 80574 78203 80585 78267
rect 80499 78183 80585 78203
rect 81587 78747 81673 78767
rect 81587 78683 81598 78747
rect 81662 78683 81673 78747
rect 81587 78667 81673 78683
rect 81587 78603 81598 78667
rect 81662 78603 81673 78667
rect 81587 78587 81673 78603
rect 81587 78523 81598 78587
rect 81662 78523 81673 78587
rect 81587 78507 81673 78523
rect 81587 78443 81598 78507
rect 81662 78443 81673 78507
rect 81587 78427 81673 78443
rect 81587 78363 81598 78427
rect 81662 78363 81673 78427
rect 81587 78347 81673 78363
rect 81587 78283 81598 78347
rect 81662 78283 81673 78347
rect 81587 78267 81673 78283
rect 81587 78203 81598 78267
rect 81662 78203 81673 78267
rect 81587 78183 81673 78203
rect 82675 78747 82761 78767
rect 82675 78683 82686 78747
rect 82750 78683 82761 78747
rect 82675 78667 82761 78683
rect 82675 78603 82686 78667
rect 82750 78603 82761 78667
rect 82675 78587 82761 78603
rect 82675 78523 82686 78587
rect 82750 78523 82761 78587
rect 82675 78507 82761 78523
rect 82675 78443 82686 78507
rect 82750 78443 82761 78507
rect 82675 78427 82761 78443
rect 82675 78363 82686 78427
rect 82750 78363 82761 78427
rect 82675 78347 82761 78363
rect 82675 78283 82686 78347
rect 82750 78283 82761 78347
rect 82675 78267 82761 78283
rect 82675 78203 82686 78267
rect 82750 78203 82761 78267
rect 82675 78183 82761 78203
rect 83763 78747 83849 78767
rect 83763 78683 83774 78747
rect 83838 78683 83849 78747
rect 83763 78667 83849 78683
rect 83763 78603 83774 78667
rect 83838 78603 83849 78667
rect 83763 78587 83849 78603
rect 83763 78523 83774 78587
rect 83838 78523 83849 78587
rect 83763 78507 83849 78523
rect 83763 78443 83774 78507
rect 83838 78443 83849 78507
rect 83763 78427 83849 78443
rect 83763 78363 83774 78427
rect 83838 78363 83849 78427
rect 83763 78347 83849 78363
rect 83763 78283 83774 78347
rect 83838 78283 83849 78347
rect 83763 78267 83849 78283
rect 83763 78203 83774 78267
rect 83838 78203 83849 78267
rect 83763 78183 83849 78203
rect 84851 78747 84937 78767
rect 84851 78683 84862 78747
rect 84926 78683 84937 78747
rect 84851 78667 84937 78683
rect 84851 78603 84862 78667
rect 84926 78603 84937 78667
rect 84851 78587 84937 78603
rect 84851 78523 84862 78587
rect 84926 78523 84937 78587
rect 84851 78507 84937 78523
rect 84851 78443 84862 78507
rect 84926 78443 84937 78507
rect 84851 78427 84937 78443
rect 84851 78363 84862 78427
rect 84926 78363 84937 78427
rect 84851 78347 84937 78363
rect 84851 78283 84862 78347
rect 84926 78283 84937 78347
rect 84851 78267 84937 78283
rect 84851 78203 84862 78267
rect 84926 78203 84937 78267
rect 84851 78183 84937 78203
rect 85939 78747 86025 78767
rect 85939 78683 85950 78747
rect 86014 78683 86025 78747
rect 85939 78667 86025 78683
rect 85939 78603 85950 78667
rect 86014 78603 86025 78667
rect 85939 78587 86025 78603
rect 85939 78523 85950 78587
rect 86014 78523 86025 78587
rect 85939 78507 86025 78523
rect 85939 78443 85950 78507
rect 86014 78443 86025 78507
rect 85939 78427 86025 78443
rect 85939 78363 85950 78427
rect 86014 78363 86025 78427
rect 85939 78347 86025 78363
rect 85939 78283 85950 78347
rect 86014 78283 86025 78347
rect 85939 78267 86025 78283
rect 85939 78203 85950 78267
rect 86014 78203 86025 78267
rect 85939 78183 86025 78203
rect 87027 78747 87113 78767
rect 87027 78683 87038 78747
rect 87102 78683 87113 78747
rect 87027 78667 87113 78683
rect 87027 78603 87038 78667
rect 87102 78603 87113 78667
rect 87027 78587 87113 78603
rect 87027 78523 87038 78587
rect 87102 78523 87113 78587
rect 87027 78507 87113 78523
rect 87027 78443 87038 78507
rect 87102 78443 87113 78507
rect 87027 78427 87113 78443
rect 87027 78363 87038 78427
rect 87102 78363 87113 78427
rect 87027 78347 87113 78363
rect 87027 78283 87038 78347
rect 87102 78283 87113 78347
rect 87027 78267 87113 78283
rect 87027 78203 87038 78267
rect 87102 78203 87113 78267
rect 87027 78183 87113 78203
rect 88115 78747 88201 78767
rect 88115 78683 88126 78747
rect 88190 78683 88201 78747
rect 88115 78667 88201 78683
rect 88115 78603 88126 78667
rect 88190 78603 88201 78667
rect 88115 78587 88201 78603
rect 88115 78523 88126 78587
rect 88190 78523 88201 78587
rect 88115 78507 88201 78523
rect 88115 78443 88126 78507
rect 88190 78443 88201 78507
rect 88115 78427 88201 78443
rect 88115 78363 88126 78427
rect 88190 78363 88201 78427
rect 88115 78347 88201 78363
rect 88115 78283 88126 78347
rect 88190 78283 88201 78347
rect 88115 78267 88201 78283
rect 88115 78203 88126 78267
rect 88190 78203 88201 78267
rect 88115 78183 88201 78203
rect 74514 76750 74600 76770
rect 74514 76686 74525 76750
rect 74589 76686 74600 76750
rect 74514 76670 74600 76686
rect 74514 76606 74525 76670
rect 74589 76606 74600 76670
rect 74514 76590 74600 76606
rect 74514 76526 74525 76590
rect 74589 76526 74600 76590
rect 74514 76510 74600 76526
rect 74514 76446 74525 76510
rect 74589 76446 74600 76510
rect 74514 76430 74600 76446
rect 74514 76366 74525 76430
rect 74589 76366 74600 76430
rect 74514 76350 74600 76366
rect 74514 76286 74525 76350
rect 74589 76286 74600 76350
rect 74514 76270 74600 76286
rect 74514 76206 74525 76270
rect 74589 76206 74600 76270
rect 74514 76186 74600 76206
rect 75602 76750 75688 76770
rect 75602 76686 75613 76750
rect 75677 76686 75688 76750
rect 75602 76670 75688 76686
rect 75602 76606 75613 76670
rect 75677 76606 75688 76670
rect 75602 76590 75688 76606
rect 75602 76526 75613 76590
rect 75677 76526 75688 76590
rect 75602 76510 75688 76526
rect 75602 76446 75613 76510
rect 75677 76446 75688 76510
rect 75602 76430 75688 76446
rect 75602 76366 75613 76430
rect 75677 76366 75688 76430
rect 75602 76350 75688 76366
rect 75602 76286 75613 76350
rect 75677 76286 75688 76350
rect 75602 76270 75688 76286
rect 75602 76206 75613 76270
rect 75677 76206 75688 76270
rect 75602 76186 75688 76206
rect 76690 76750 76776 76770
rect 76690 76686 76701 76750
rect 76765 76686 76776 76750
rect 76690 76670 76776 76686
rect 76690 76606 76701 76670
rect 76765 76606 76776 76670
rect 76690 76590 76776 76606
rect 76690 76526 76701 76590
rect 76765 76526 76776 76590
rect 76690 76510 76776 76526
rect 76690 76446 76701 76510
rect 76765 76446 76776 76510
rect 76690 76430 76776 76446
rect 76690 76366 76701 76430
rect 76765 76366 76776 76430
rect 76690 76350 76776 76366
rect 76690 76286 76701 76350
rect 76765 76286 76776 76350
rect 76690 76270 76776 76286
rect 76690 76206 76701 76270
rect 76765 76206 76776 76270
rect 76690 76186 76776 76206
rect 77778 76750 77864 76770
rect 77778 76686 77789 76750
rect 77853 76686 77864 76750
rect 77778 76670 77864 76686
rect 77778 76606 77789 76670
rect 77853 76606 77864 76670
rect 77778 76590 77864 76606
rect 77778 76526 77789 76590
rect 77853 76526 77864 76590
rect 77778 76510 77864 76526
rect 77778 76446 77789 76510
rect 77853 76446 77864 76510
rect 77778 76430 77864 76446
rect 77778 76366 77789 76430
rect 77853 76366 77864 76430
rect 77778 76350 77864 76366
rect 77778 76286 77789 76350
rect 77853 76286 77864 76350
rect 77778 76270 77864 76286
rect 77778 76206 77789 76270
rect 77853 76206 77864 76270
rect 77778 76186 77864 76206
rect 78866 76750 78952 76770
rect 78866 76686 78877 76750
rect 78941 76686 78952 76750
rect 78866 76670 78952 76686
rect 78866 76606 78877 76670
rect 78941 76606 78952 76670
rect 78866 76590 78952 76606
rect 78866 76526 78877 76590
rect 78941 76526 78952 76590
rect 78866 76510 78952 76526
rect 78866 76446 78877 76510
rect 78941 76446 78952 76510
rect 78866 76430 78952 76446
rect 78866 76366 78877 76430
rect 78941 76366 78952 76430
rect 78866 76350 78952 76366
rect 78866 76286 78877 76350
rect 78941 76286 78952 76350
rect 78866 76270 78952 76286
rect 78866 76206 78877 76270
rect 78941 76206 78952 76270
rect 78866 76186 78952 76206
rect 79954 76750 80040 76770
rect 79954 76686 79965 76750
rect 80029 76686 80040 76750
rect 79954 76670 80040 76686
rect 79954 76606 79965 76670
rect 80029 76606 80040 76670
rect 79954 76590 80040 76606
rect 79954 76526 79965 76590
rect 80029 76526 80040 76590
rect 79954 76510 80040 76526
rect 79954 76446 79965 76510
rect 80029 76446 80040 76510
rect 79954 76430 80040 76446
rect 79954 76366 79965 76430
rect 80029 76366 80040 76430
rect 79954 76350 80040 76366
rect 79954 76286 79965 76350
rect 80029 76286 80040 76350
rect 79954 76270 80040 76286
rect 79954 76206 79965 76270
rect 80029 76206 80040 76270
rect 79954 76186 80040 76206
rect 81042 76750 81128 76770
rect 81042 76686 81053 76750
rect 81117 76686 81128 76750
rect 81042 76670 81128 76686
rect 81042 76606 81053 76670
rect 81117 76606 81128 76670
rect 81042 76590 81128 76606
rect 81042 76526 81053 76590
rect 81117 76526 81128 76590
rect 81042 76510 81128 76526
rect 81042 76446 81053 76510
rect 81117 76446 81128 76510
rect 81042 76430 81128 76446
rect 81042 76366 81053 76430
rect 81117 76366 81128 76430
rect 81042 76350 81128 76366
rect 81042 76286 81053 76350
rect 81117 76286 81128 76350
rect 81042 76270 81128 76286
rect 81042 76206 81053 76270
rect 81117 76206 81128 76270
rect 81042 76186 81128 76206
rect 82130 76750 82216 76770
rect 82130 76686 82141 76750
rect 82205 76686 82216 76750
rect 82130 76670 82216 76686
rect 82130 76606 82141 76670
rect 82205 76606 82216 76670
rect 82130 76590 82216 76606
rect 82130 76526 82141 76590
rect 82205 76526 82216 76590
rect 82130 76510 82216 76526
rect 82130 76446 82141 76510
rect 82205 76446 82216 76510
rect 82130 76430 82216 76446
rect 82130 76366 82141 76430
rect 82205 76366 82216 76430
rect 82130 76350 82216 76366
rect 82130 76286 82141 76350
rect 82205 76286 82216 76350
rect 82130 76270 82216 76286
rect 82130 76206 82141 76270
rect 82205 76206 82216 76270
rect 82130 76186 82216 76206
rect 83218 76750 83304 76770
rect 83218 76686 83229 76750
rect 83293 76686 83304 76750
rect 83218 76670 83304 76686
rect 83218 76606 83229 76670
rect 83293 76606 83304 76670
rect 83218 76590 83304 76606
rect 83218 76526 83229 76590
rect 83293 76526 83304 76590
rect 83218 76510 83304 76526
rect 83218 76446 83229 76510
rect 83293 76446 83304 76510
rect 83218 76430 83304 76446
rect 83218 76366 83229 76430
rect 83293 76366 83304 76430
rect 83218 76350 83304 76366
rect 83218 76286 83229 76350
rect 83293 76286 83304 76350
rect 83218 76270 83304 76286
rect 83218 76206 83229 76270
rect 83293 76206 83304 76270
rect 83218 76186 83304 76206
rect 84306 76750 84392 76770
rect 84306 76686 84317 76750
rect 84381 76686 84392 76750
rect 84306 76670 84392 76686
rect 84306 76606 84317 76670
rect 84381 76606 84392 76670
rect 84306 76590 84392 76606
rect 84306 76526 84317 76590
rect 84381 76526 84392 76590
rect 84306 76510 84392 76526
rect 84306 76446 84317 76510
rect 84381 76446 84392 76510
rect 84306 76430 84392 76446
rect 84306 76366 84317 76430
rect 84381 76366 84392 76430
rect 84306 76350 84392 76366
rect 84306 76286 84317 76350
rect 84381 76286 84392 76350
rect 84306 76270 84392 76286
rect 84306 76206 84317 76270
rect 84381 76206 84392 76270
rect 84306 76186 84392 76206
rect 85394 76750 85480 76770
rect 85394 76686 85405 76750
rect 85469 76686 85480 76750
rect 85394 76670 85480 76686
rect 85394 76606 85405 76670
rect 85469 76606 85480 76670
rect 85394 76590 85480 76606
rect 85394 76526 85405 76590
rect 85469 76526 85480 76590
rect 85394 76510 85480 76526
rect 85394 76446 85405 76510
rect 85469 76446 85480 76510
rect 85394 76430 85480 76446
rect 85394 76366 85405 76430
rect 85469 76366 85480 76430
rect 85394 76350 85480 76366
rect 85394 76286 85405 76350
rect 85469 76286 85480 76350
rect 85394 76270 85480 76286
rect 85394 76206 85405 76270
rect 85469 76206 85480 76270
rect 85394 76186 85480 76206
rect 86482 76750 86568 76770
rect 86482 76686 86493 76750
rect 86557 76686 86568 76750
rect 86482 76670 86568 76686
rect 86482 76606 86493 76670
rect 86557 76606 86568 76670
rect 86482 76590 86568 76606
rect 86482 76526 86493 76590
rect 86557 76526 86568 76590
rect 86482 76510 86568 76526
rect 86482 76446 86493 76510
rect 86557 76446 86568 76510
rect 86482 76430 86568 76446
rect 86482 76366 86493 76430
rect 86557 76366 86568 76430
rect 86482 76350 86568 76366
rect 86482 76286 86493 76350
rect 86557 76286 86568 76350
rect 86482 76270 86568 76286
rect 86482 76206 86493 76270
rect 86557 76206 86568 76270
rect 86482 76186 86568 76206
rect 87570 76750 87656 76770
rect 87570 76686 87581 76750
rect 87645 76686 87656 76750
rect 87570 76670 87656 76686
rect 87570 76606 87581 76670
rect 87645 76606 87656 76670
rect 87570 76590 87656 76606
rect 87570 76526 87581 76590
rect 87645 76526 87656 76590
rect 87570 76510 87656 76526
rect 87570 76446 87581 76510
rect 87645 76446 87656 76510
rect 87570 76430 87656 76446
rect 87570 76366 87581 76430
rect 87645 76366 87656 76430
rect 87570 76350 87656 76366
rect 87570 76286 87581 76350
rect 87645 76286 87656 76350
rect 87570 76270 87656 76286
rect 87570 76206 87581 76270
rect 87645 76206 87656 76270
rect 87570 76186 87656 76206
rect 88658 76750 88744 76770
rect 88658 76686 88669 76750
rect 88733 76686 88744 76750
rect 88658 76670 88744 76686
rect 88658 76606 88669 76670
rect 88733 76606 88744 76670
rect 88658 76590 88744 76606
rect 88658 76526 88669 76590
rect 88733 76526 88744 76590
rect 88658 76510 88744 76526
rect 88658 76446 88669 76510
rect 88733 76446 88744 76510
rect 88658 76430 88744 76446
rect 88658 76366 88669 76430
rect 88733 76366 88744 76430
rect 88658 76350 88744 76366
rect 88658 76286 88669 76350
rect 88733 76286 88744 76350
rect 88658 76270 88744 76286
rect 88658 76206 88669 76270
rect 88733 76206 88744 76270
rect 88658 76186 88744 76206
rect 75059 74747 75145 74767
rect 75059 74683 75070 74747
rect 75134 74683 75145 74747
rect 75059 74667 75145 74683
rect 75059 74603 75070 74667
rect 75134 74603 75145 74667
rect 75059 74587 75145 74603
rect 75059 74523 75070 74587
rect 75134 74523 75145 74587
rect 75059 74507 75145 74523
rect 75059 74443 75070 74507
rect 75134 74443 75145 74507
rect 75059 74427 75145 74443
rect 75059 74363 75070 74427
rect 75134 74363 75145 74427
rect 75059 74347 75145 74363
rect 75059 74283 75070 74347
rect 75134 74283 75145 74347
rect 75059 74267 75145 74283
rect 75059 74203 75070 74267
rect 75134 74203 75145 74267
rect 75059 74183 75145 74203
rect 77235 74747 77321 74767
rect 77235 74683 77246 74747
rect 77310 74683 77321 74747
rect 77235 74667 77321 74683
rect 77235 74603 77246 74667
rect 77310 74603 77321 74667
rect 77235 74587 77321 74603
rect 77235 74523 77246 74587
rect 77310 74523 77321 74587
rect 77235 74507 77321 74523
rect 77235 74443 77246 74507
rect 77310 74443 77321 74507
rect 77235 74427 77321 74443
rect 77235 74363 77246 74427
rect 77310 74363 77321 74427
rect 77235 74347 77321 74363
rect 77235 74283 77246 74347
rect 77310 74283 77321 74347
rect 77235 74267 77321 74283
rect 77235 74203 77246 74267
rect 77310 74203 77321 74267
rect 77235 74183 77321 74203
rect 78323 74747 78409 74767
rect 78323 74683 78334 74747
rect 78398 74683 78409 74747
rect 78323 74667 78409 74683
rect 78323 74603 78334 74667
rect 78398 74603 78409 74667
rect 78323 74587 78409 74603
rect 78323 74523 78334 74587
rect 78398 74523 78409 74587
rect 78323 74507 78409 74523
rect 78323 74443 78334 74507
rect 78398 74443 78409 74507
rect 78323 74427 78409 74443
rect 78323 74363 78334 74427
rect 78398 74363 78409 74427
rect 78323 74347 78409 74363
rect 78323 74283 78334 74347
rect 78398 74283 78409 74347
rect 78323 74267 78409 74283
rect 78323 74203 78334 74267
rect 78398 74203 78409 74267
rect 78323 74183 78409 74203
rect 80499 74747 80585 74767
rect 80499 74683 80510 74747
rect 80574 74683 80585 74747
rect 80499 74667 80585 74683
rect 80499 74603 80510 74667
rect 80574 74603 80585 74667
rect 80499 74587 80585 74603
rect 80499 74523 80510 74587
rect 80574 74523 80585 74587
rect 80499 74507 80585 74523
rect 80499 74443 80510 74507
rect 80574 74443 80585 74507
rect 80499 74427 80585 74443
rect 80499 74363 80510 74427
rect 80574 74363 80585 74427
rect 80499 74347 80585 74363
rect 80499 74283 80510 74347
rect 80574 74283 80585 74347
rect 80499 74267 80585 74283
rect 80499 74203 80510 74267
rect 80574 74203 80585 74267
rect 80499 74183 80585 74203
rect 81587 74747 81673 74767
rect 81587 74683 81598 74747
rect 81662 74683 81673 74747
rect 81587 74667 81673 74683
rect 81587 74603 81598 74667
rect 81662 74603 81673 74667
rect 81587 74587 81673 74603
rect 81587 74523 81598 74587
rect 81662 74523 81673 74587
rect 81587 74507 81673 74523
rect 81587 74443 81598 74507
rect 81662 74443 81673 74507
rect 81587 74427 81673 74443
rect 81587 74363 81598 74427
rect 81662 74363 81673 74427
rect 81587 74347 81673 74363
rect 81587 74283 81598 74347
rect 81662 74283 81673 74347
rect 81587 74267 81673 74283
rect 81587 74203 81598 74267
rect 81662 74203 81673 74267
rect 81587 74183 81673 74203
rect 82675 74747 82761 74767
rect 82675 74683 82686 74747
rect 82750 74683 82761 74747
rect 82675 74667 82761 74683
rect 82675 74603 82686 74667
rect 82750 74603 82761 74667
rect 82675 74587 82761 74603
rect 82675 74523 82686 74587
rect 82750 74523 82761 74587
rect 82675 74507 82761 74523
rect 82675 74443 82686 74507
rect 82750 74443 82761 74507
rect 82675 74427 82761 74443
rect 82675 74363 82686 74427
rect 82750 74363 82761 74427
rect 82675 74347 82761 74363
rect 82675 74283 82686 74347
rect 82750 74283 82761 74347
rect 82675 74267 82761 74283
rect 82675 74203 82686 74267
rect 82750 74203 82761 74267
rect 82675 74183 82761 74203
rect 84851 74747 84937 74767
rect 84851 74683 84862 74747
rect 84926 74683 84937 74747
rect 84851 74667 84937 74683
rect 84851 74603 84862 74667
rect 84926 74603 84937 74667
rect 84851 74587 84937 74603
rect 84851 74523 84862 74587
rect 84926 74523 84937 74587
rect 84851 74507 84937 74523
rect 84851 74443 84862 74507
rect 84926 74443 84937 74507
rect 84851 74427 84937 74443
rect 84851 74363 84862 74427
rect 84926 74363 84937 74427
rect 84851 74347 84937 74363
rect 84851 74283 84862 74347
rect 84926 74283 84937 74347
rect 84851 74267 84937 74283
rect 84851 74203 84862 74267
rect 84926 74203 84937 74267
rect 84851 74183 84937 74203
rect 85939 74747 86025 74767
rect 85939 74683 85950 74747
rect 86014 74683 86025 74747
rect 85939 74667 86025 74683
rect 85939 74603 85950 74667
rect 86014 74603 86025 74667
rect 85939 74587 86025 74603
rect 85939 74523 85950 74587
rect 86014 74523 86025 74587
rect 85939 74507 86025 74523
rect 85939 74443 85950 74507
rect 86014 74443 86025 74507
rect 85939 74427 86025 74443
rect 85939 74363 85950 74427
rect 86014 74363 86025 74427
rect 85939 74347 86025 74363
rect 85939 74283 85950 74347
rect 86014 74283 86025 74347
rect 85939 74267 86025 74283
rect 85939 74203 85950 74267
rect 86014 74203 86025 74267
rect 85939 74183 86025 74203
rect 88115 74747 88201 74767
rect 88115 74683 88126 74747
rect 88190 74683 88201 74747
rect 88115 74667 88201 74683
rect 88115 74603 88126 74667
rect 88190 74603 88201 74667
rect 88115 74587 88201 74603
rect 88115 74523 88126 74587
rect 88190 74523 88201 74587
rect 88115 74507 88201 74523
rect 88115 74443 88126 74507
rect 88190 74443 88201 74507
rect 88115 74427 88201 74443
rect 88115 74363 88126 74427
rect 88190 74363 88201 74427
rect 88115 74347 88201 74363
rect 88115 74283 88126 74347
rect 88190 74283 88201 74347
rect 88115 74267 88201 74283
rect 88115 74203 88126 74267
rect 88190 74203 88201 74267
rect 88115 74183 88201 74203
rect 74514 72750 74600 72770
rect 74514 72686 74525 72750
rect 74589 72686 74600 72750
rect 74514 72670 74600 72686
rect 74514 72606 74525 72670
rect 74589 72606 74600 72670
rect 74514 72590 74600 72606
rect 74514 72526 74525 72590
rect 74589 72526 74600 72590
rect 74514 72510 74600 72526
rect 74514 72446 74525 72510
rect 74589 72446 74600 72510
rect 74514 72430 74600 72446
rect 74514 72366 74525 72430
rect 74589 72366 74600 72430
rect 74514 72350 74600 72366
rect 74514 72286 74525 72350
rect 74589 72286 74600 72350
rect 74514 72270 74600 72286
rect 74514 72206 74525 72270
rect 74589 72206 74600 72270
rect 74514 72186 74600 72206
rect 75602 72750 75688 72770
rect 75602 72686 75613 72750
rect 75677 72686 75688 72750
rect 75602 72670 75688 72686
rect 75602 72606 75613 72670
rect 75677 72606 75688 72670
rect 75602 72590 75688 72606
rect 75602 72526 75613 72590
rect 75677 72526 75688 72590
rect 75602 72510 75688 72526
rect 75602 72446 75613 72510
rect 75677 72446 75688 72510
rect 75602 72430 75688 72446
rect 75602 72366 75613 72430
rect 75677 72366 75688 72430
rect 75602 72350 75688 72366
rect 75602 72286 75613 72350
rect 75677 72286 75688 72350
rect 75602 72270 75688 72286
rect 75602 72206 75613 72270
rect 75677 72206 75688 72270
rect 75602 72186 75688 72206
rect 76690 72750 76776 72770
rect 76690 72686 76701 72750
rect 76765 72686 76776 72750
rect 76690 72670 76776 72686
rect 76690 72606 76701 72670
rect 76765 72606 76776 72670
rect 76690 72590 76776 72606
rect 76690 72526 76701 72590
rect 76765 72526 76776 72590
rect 76690 72510 76776 72526
rect 76690 72446 76701 72510
rect 76765 72446 76776 72510
rect 76690 72430 76776 72446
rect 76690 72366 76701 72430
rect 76765 72366 76776 72430
rect 76690 72350 76776 72366
rect 76690 72286 76701 72350
rect 76765 72286 76776 72350
rect 76690 72270 76776 72286
rect 76690 72206 76701 72270
rect 76765 72206 76776 72270
rect 76690 72186 76776 72206
rect 77778 72750 77864 72770
rect 77778 72686 77789 72750
rect 77853 72686 77864 72750
rect 77778 72670 77864 72686
rect 77778 72606 77789 72670
rect 77853 72606 77864 72670
rect 77778 72590 77864 72606
rect 77778 72526 77789 72590
rect 77853 72526 77864 72590
rect 77778 72510 77864 72526
rect 77778 72446 77789 72510
rect 77853 72446 77864 72510
rect 77778 72430 77864 72446
rect 77778 72366 77789 72430
rect 77853 72366 77864 72430
rect 77778 72350 77864 72366
rect 77778 72286 77789 72350
rect 77853 72286 77864 72350
rect 77778 72270 77864 72286
rect 77778 72206 77789 72270
rect 77853 72206 77864 72270
rect 77778 72186 77864 72206
rect 78866 72750 78952 72770
rect 78866 72686 78877 72750
rect 78941 72686 78952 72750
rect 78866 72670 78952 72686
rect 78866 72606 78877 72670
rect 78941 72606 78952 72670
rect 78866 72590 78952 72606
rect 78866 72526 78877 72590
rect 78941 72526 78952 72590
rect 78866 72510 78952 72526
rect 78866 72446 78877 72510
rect 78941 72446 78952 72510
rect 78866 72430 78952 72446
rect 78866 72366 78877 72430
rect 78941 72366 78952 72430
rect 78866 72350 78952 72366
rect 78866 72286 78877 72350
rect 78941 72286 78952 72350
rect 78866 72270 78952 72286
rect 78866 72206 78877 72270
rect 78941 72206 78952 72270
rect 78866 72186 78952 72206
rect 79954 72750 80040 72770
rect 79954 72686 79965 72750
rect 80029 72686 80040 72750
rect 79954 72670 80040 72686
rect 79954 72606 79965 72670
rect 80029 72606 80040 72670
rect 79954 72590 80040 72606
rect 79954 72526 79965 72590
rect 80029 72526 80040 72590
rect 79954 72510 80040 72526
rect 79954 72446 79965 72510
rect 80029 72446 80040 72510
rect 79954 72430 80040 72446
rect 79954 72366 79965 72430
rect 80029 72366 80040 72430
rect 79954 72350 80040 72366
rect 79954 72286 79965 72350
rect 80029 72286 80040 72350
rect 79954 72270 80040 72286
rect 79954 72206 79965 72270
rect 80029 72206 80040 72270
rect 79954 72186 80040 72206
rect 81042 72750 81128 72770
rect 81042 72686 81053 72750
rect 81117 72686 81128 72750
rect 81042 72670 81128 72686
rect 81042 72606 81053 72670
rect 81117 72606 81128 72670
rect 81042 72590 81128 72606
rect 81042 72526 81053 72590
rect 81117 72526 81128 72590
rect 81042 72510 81128 72526
rect 81042 72446 81053 72510
rect 81117 72446 81128 72510
rect 81042 72430 81128 72446
rect 81042 72366 81053 72430
rect 81117 72366 81128 72430
rect 81042 72350 81128 72366
rect 81042 72286 81053 72350
rect 81117 72286 81128 72350
rect 81042 72270 81128 72286
rect 81042 72206 81053 72270
rect 81117 72206 81128 72270
rect 81042 72186 81128 72206
rect 86482 72750 86568 72770
rect 86482 72686 86493 72750
rect 86557 72686 86568 72750
rect 86482 72670 86568 72686
rect 86482 72606 86493 72670
rect 86557 72606 86568 72670
rect 86482 72590 86568 72606
rect 86482 72526 86493 72590
rect 86557 72526 86568 72590
rect 86482 72510 86568 72526
rect 86482 72446 86493 72510
rect 86557 72446 86568 72510
rect 86482 72430 86568 72446
rect 86482 72366 86493 72430
rect 86557 72366 86568 72430
rect 86482 72350 86568 72366
rect 86482 72286 86493 72350
rect 86557 72286 86568 72350
rect 86482 72270 86568 72286
rect 86482 72206 86493 72270
rect 86557 72206 86568 72270
rect 86482 72186 86568 72206
rect 87570 72750 87656 72770
rect 87570 72686 87581 72750
rect 87645 72686 87656 72750
rect 87570 72670 87656 72686
rect 87570 72606 87581 72670
rect 87645 72606 87656 72670
rect 87570 72590 87656 72606
rect 87570 72526 87581 72590
rect 87645 72526 87656 72590
rect 87570 72510 87656 72526
rect 87570 72446 87581 72510
rect 87645 72446 87656 72510
rect 87570 72430 87656 72446
rect 87570 72366 87581 72430
rect 87645 72366 87656 72430
rect 87570 72350 87656 72366
rect 87570 72286 87581 72350
rect 87645 72286 87656 72350
rect 87570 72270 87656 72286
rect 87570 72206 87581 72270
rect 87645 72206 87656 72270
rect 87570 72186 87656 72206
rect 88658 72750 88744 72770
rect 88658 72686 88669 72750
rect 88733 72686 88744 72750
rect 88658 72670 88744 72686
rect 88658 72606 88669 72670
rect 88733 72606 88744 72670
rect 88658 72590 88744 72606
rect 88658 72526 88669 72590
rect 88733 72526 88744 72590
rect 88658 72510 88744 72526
rect 88658 72446 88669 72510
rect 88733 72446 88744 72510
rect 88658 72430 88744 72446
rect 88658 72366 88669 72430
rect 88733 72366 88744 72430
rect 88658 72350 88744 72366
rect 88658 72286 88669 72350
rect 88733 72286 88744 72350
rect 88658 72270 88744 72286
rect 88658 72206 88669 72270
rect 88733 72206 88744 72270
rect 88658 72186 88744 72206
rect 67261 71634 67655 71656
rect 33596 71214 45733 71278
rect 45797 71214 50683 71278
rect 50747 71214 50757 71278
rect 29997 67300 30114 67340
rect 29997 67236 30023 67300
rect 30087 67236 30114 67300
rect 29997 67220 30114 67236
rect 29997 67156 30023 67220
rect 30087 67156 30114 67220
rect 29997 67140 30114 67156
rect 29997 67076 30023 67140
rect 30087 67076 30114 67140
rect 29997 67060 30114 67076
rect 29997 66996 30023 67060
rect 30087 66996 30114 67060
rect 29997 66980 30114 66996
rect 29997 66916 30023 66980
rect 30087 66916 30114 66980
rect 29997 66900 30114 66916
rect 29997 66836 30023 66900
rect 30087 66836 30114 66900
rect 29997 66796 30114 66836
rect 30002 66159 30109 66196
rect 30002 66095 30023 66159
rect 30087 66095 30109 66159
rect 30002 66079 30109 66095
rect 30002 66015 30023 66079
rect 30087 66015 30109 66079
rect 30002 65999 30109 66015
rect 30002 65935 30023 65999
rect 30087 65935 30109 65999
rect 30002 65919 30109 65935
rect 30002 65855 30023 65919
rect 30087 65855 30109 65919
rect 30002 65839 30109 65855
rect 30002 65775 30023 65839
rect 30087 65775 30109 65839
rect 30002 65759 30109 65775
rect 30002 65695 30023 65759
rect 30087 65695 30109 65759
rect 30002 65679 30109 65695
rect 30002 65615 30023 65679
rect 30087 65615 30109 65679
rect 30002 65599 30109 65615
rect 30002 65535 30023 65599
rect 30087 65535 30109 65599
rect 30002 65519 30109 65535
rect 30002 65455 30023 65519
rect 30087 65455 30109 65519
rect 30002 65439 30109 65455
rect 30002 65375 30023 65439
rect 30087 65375 30109 65439
rect 30002 65359 30109 65375
rect 30002 65295 30023 65359
rect 30087 65295 30109 65359
rect 30002 65279 30109 65295
rect 30002 65215 30023 65279
rect 30087 65215 30109 65279
rect 30002 65199 30109 65215
rect 30002 65135 30023 65199
rect 30087 65135 30109 65199
rect 30002 65119 30109 65135
rect 30002 65055 30023 65119
rect 30087 65055 30109 65119
rect 30002 65019 30109 65055
rect 30007 64633 30114 64670
rect 30007 64569 30028 64633
rect 30092 64569 30114 64633
rect 30007 64553 30114 64569
rect 30007 64489 30028 64553
rect 30092 64489 30114 64553
rect 30007 64473 30114 64489
rect 30007 64409 30028 64473
rect 30092 64409 30114 64473
rect 30007 64393 30114 64409
rect 30007 64329 30028 64393
rect 30092 64329 30114 64393
rect 30007 64313 30114 64329
rect 30007 64249 30028 64313
rect 30092 64249 30114 64313
rect 30007 64233 30114 64249
rect 30007 64169 30028 64233
rect 30092 64169 30114 64233
rect 30007 64153 30114 64169
rect 30007 64089 30028 64153
rect 30092 64089 30114 64153
rect 30007 64073 30114 64089
rect 30007 64009 30028 64073
rect 30092 64009 30114 64073
rect 30007 63993 30114 64009
rect 30007 63929 30028 63993
rect 30092 63929 30114 63993
rect 30007 63913 30114 63929
rect 30007 63849 30028 63913
rect 30092 63849 30114 63913
rect 30007 63833 30114 63849
rect 30007 63769 30028 63833
rect 30092 63769 30114 63833
rect 30007 63753 30114 63769
rect 30007 63689 30028 63753
rect 30092 63689 30114 63753
rect 30007 63673 30114 63689
rect 30007 63609 30028 63673
rect 30092 63609 30114 63673
rect 30007 63593 30114 63609
rect 30007 63529 30028 63593
rect 30092 63529 30114 63593
rect 30007 63493 30114 63529
rect 25272 63170 25356 63193
rect 25272 63106 25282 63170
rect 25346 63106 25356 63170
rect 25272 63090 25356 63106
rect 25272 63026 25282 63090
rect 25346 63026 25356 63090
rect 25272 63010 25356 63026
rect 25272 62946 25282 63010
rect 25346 62946 25356 63010
rect 25272 62930 25356 62946
rect 25272 62866 25282 62930
rect 25346 62866 25356 62930
rect 25272 62844 25356 62866
rect 30002 63130 30106 63147
rect 30002 63066 30022 63130
rect 30086 63066 30106 63130
rect 30002 63050 30106 63066
rect 30002 62986 30022 63050
rect 30086 62986 30106 63050
rect 30002 62970 30106 62986
rect 30002 62906 30022 62970
rect 30086 62906 30106 62970
rect 30002 62890 30106 62906
rect 30002 62826 30022 62890
rect 30086 62826 30106 62890
rect 30002 62810 30106 62826
rect 30002 62746 30022 62810
rect 30086 62746 30106 62810
rect 30002 62730 30106 62746
rect 30002 62666 30022 62730
rect 30086 62666 30106 62730
rect 30002 62650 30106 62666
rect 25273 62631 25357 62640
rect 25273 62567 25283 62631
rect 25347 62567 25357 62631
rect 25273 62551 25357 62567
rect 25273 62487 25283 62551
rect 25347 62487 25357 62551
rect 25273 62471 25357 62487
rect 25273 62407 25283 62471
rect 25347 62407 25357 62471
rect 30002 62586 30022 62650
rect 30086 62586 30106 62650
rect 30002 62570 30106 62586
rect 30002 62506 30022 62570
rect 30086 62506 30106 62570
rect 30002 62490 30106 62506
rect 25273 62391 25357 62407
rect 25273 62327 25283 62391
rect 25347 62327 25357 62391
rect 27470 62435 27954 62440
rect 27470 62371 27480 62435
rect 27544 62371 27560 62435
rect 27624 62371 27640 62435
rect 27704 62371 27720 62435
rect 27784 62371 27800 62435
rect 27864 62371 27880 62435
rect 27944 62371 27954 62435
rect 27470 62366 27954 62371
rect 30002 62426 30022 62490
rect 30086 62426 30106 62490
rect 30002 62410 30106 62426
rect 25273 62311 25357 62327
rect 25273 62247 25283 62311
rect 25347 62247 25357 62311
rect 30002 62346 30022 62410
rect 30086 62346 30106 62410
rect 30002 62330 30106 62346
rect 30002 62266 30022 62330
rect 30086 62266 30106 62330
rect 30002 62249 30106 62266
rect 25273 62231 25357 62247
rect 25273 62167 25283 62231
rect 25347 62167 25357 62231
rect 25273 62158 25357 62167
rect 33596 61824 33660 71214
rect 75059 70747 75145 70767
rect 75059 70683 75070 70747
rect 75134 70683 75145 70747
rect 75059 70667 75145 70683
rect 46597 70591 46607 70655
rect 46671 70591 50683 70655
rect 50747 70591 50759 70655
rect 75059 70603 75070 70667
rect 75134 70603 75145 70667
rect 75059 70587 75145 70603
rect 75059 70523 75070 70587
rect 75134 70523 75145 70587
rect 75059 70507 75145 70523
rect 75059 70443 75070 70507
rect 75134 70443 75145 70507
rect 75059 70427 75145 70443
rect 75059 70363 75070 70427
rect 75134 70363 75145 70427
rect 75059 70347 75145 70363
rect 51160 70260 51382 70301
rect 43615 67083 43699 67088
rect 43615 67019 43625 67083
rect 43689 67019 47886 67083
rect 47950 67019 47960 67083
rect 43615 67014 43699 67019
rect 44391 66420 44475 66425
rect 44391 66356 44401 66420
rect 44465 66356 47025 66420
rect 47089 66356 47099 66420
rect 44391 66351 44475 66356
rect 35593 66185 35708 66212
rect 35593 66121 35619 66185
rect 35683 66121 35708 66185
rect 35593 66096 35708 66121
rect 51160 63939 51199 70260
rect 51127 63876 51199 63939
rect 51343 63939 51382 70260
rect 75059 70283 75070 70347
rect 75134 70283 75145 70347
rect 75059 70267 75145 70283
rect 75059 70203 75070 70267
rect 75134 70203 75145 70267
rect 75059 70183 75145 70203
rect 76147 70747 76233 70767
rect 76147 70683 76158 70747
rect 76222 70683 76233 70747
rect 76147 70667 76233 70683
rect 76147 70603 76158 70667
rect 76222 70603 76233 70667
rect 76147 70587 76233 70603
rect 76147 70523 76158 70587
rect 76222 70523 76233 70587
rect 76147 70507 76233 70523
rect 76147 70443 76158 70507
rect 76222 70443 76233 70507
rect 76147 70427 76233 70443
rect 76147 70363 76158 70427
rect 76222 70363 76233 70427
rect 76147 70347 76233 70363
rect 76147 70283 76158 70347
rect 76222 70283 76233 70347
rect 76147 70267 76233 70283
rect 76147 70203 76158 70267
rect 76222 70203 76233 70267
rect 76147 70183 76233 70203
rect 77235 70747 77321 70767
rect 77235 70683 77246 70747
rect 77310 70683 77321 70747
rect 77235 70667 77321 70683
rect 77235 70603 77246 70667
rect 77310 70603 77321 70667
rect 77235 70587 77321 70603
rect 77235 70523 77246 70587
rect 77310 70523 77321 70587
rect 77235 70507 77321 70523
rect 77235 70443 77246 70507
rect 77310 70443 77321 70507
rect 77235 70427 77321 70443
rect 77235 70363 77246 70427
rect 77310 70363 77321 70427
rect 77235 70347 77321 70363
rect 77235 70283 77246 70347
rect 77310 70283 77321 70347
rect 77235 70267 77321 70283
rect 77235 70203 77246 70267
rect 77310 70203 77321 70267
rect 77235 70183 77321 70203
rect 78323 70747 78409 70767
rect 78323 70683 78334 70747
rect 78398 70683 78409 70747
rect 78323 70667 78409 70683
rect 78323 70603 78334 70667
rect 78398 70603 78409 70667
rect 78323 70587 78409 70603
rect 78323 70523 78334 70587
rect 78398 70523 78409 70587
rect 78323 70507 78409 70523
rect 78323 70443 78334 70507
rect 78398 70443 78409 70507
rect 78323 70427 78409 70443
rect 78323 70363 78334 70427
rect 78398 70363 78409 70427
rect 78323 70347 78409 70363
rect 78323 70283 78334 70347
rect 78398 70283 78409 70347
rect 78323 70267 78409 70283
rect 78323 70203 78334 70267
rect 78398 70203 78409 70267
rect 78323 70183 78409 70203
rect 79411 70747 79497 70767
rect 79411 70683 79422 70747
rect 79486 70683 79497 70747
rect 79411 70667 79497 70683
rect 79411 70603 79422 70667
rect 79486 70603 79497 70667
rect 79411 70587 79497 70603
rect 79411 70523 79422 70587
rect 79486 70523 79497 70587
rect 79411 70507 79497 70523
rect 79411 70443 79422 70507
rect 79486 70443 79497 70507
rect 79411 70427 79497 70443
rect 79411 70363 79422 70427
rect 79486 70363 79497 70427
rect 79411 70347 79497 70363
rect 79411 70283 79422 70347
rect 79486 70283 79497 70347
rect 79411 70267 79497 70283
rect 79411 70203 79422 70267
rect 79486 70203 79497 70267
rect 79411 70183 79497 70203
rect 81587 70747 81673 70767
rect 81587 70683 81598 70747
rect 81662 70683 81673 70747
rect 81587 70667 81673 70683
rect 81587 70603 81598 70667
rect 81662 70603 81673 70667
rect 81587 70587 81673 70603
rect 81587 70523 81598 70587
rect 81662 70523 81673 70587
rect 81587 70507 81673 70523
rect 81587 70443 81598 70507
rect 81662 70443 81673 70507
rect 81587 70427 81673 70443
rect 81587 70363 81598 70427
rect 81662 70363 81673 70427
rect 81587 70347 81673 70363
rect 81587 70283 81598 70347
rect 81662 70283 81673 70347
rect 81587 70267 81673 70283
rect 81587 70203 81598 70267
rect 81662 70203 81673 70267
rect 81587 70183 81673 70203
rect 82675 70747 82761 70767
rect 82675 70683 82686 70747
rect 82750 70683 82761 70747
rect 82675 70667 82761 70683
rect 82675 70603 82686 70667
rect 82750 70603 82761 70667
rect 82675 70587 82761 70603
rect 82675 70523 82686 70587
rect 82750 70523 82761 70587
rect 82675 70507 82761 70523
rect 82675 70443 82686 70507
rect 82750 70443 82761 70507
rect 82675 70427 82761 70443
rect 82675 70363 82686 70427
rect 82750 70363 82761 70427
rect 82675 70347 82761 70363
rect 82675 70283 82686 70347
rect 82750 70283 82761 70347
rect 82675 70267 82761 70283
rect 82675 70203 82686 70267
rect 82750 70203 82761 70267
rect 82675 70183 82761 70203
rect 83763 70747 83849 70767
rect 83763 70683 83774 70747
rect 83838 70683 83849 70747
rect 83763 70667 83849 70683
rect 83763 70603 83774 70667
rect 83838 70603 83849 70667
rect 83763 70587 83849 70603
rect 83763 70523 83774 70587
rect 83838 70523 83849 70587
rect 83763 70507 83849 70523
rect 83763 70443 83774 70507
rect 83838 70443 83849 70507
rect 83763 70427 83849 70443
rect 83763 70363 83774 70427
rect 83838 70363 83849 70427
rect 83763 70347 83849 70363
rect 83763 70283 83774 70347
rect 83838 70283 83849 70347
rect 83763 70267 83849 70283
rect 83763 70203 83774 70267
rect 83838 70203 83849 70267
rect 83763 70183 83849 70203
rect 84851 70747 84937 70767
rect 84851 70683 84862 70747
rect 84926 70683 84937 70747
rect 84851 70667 84937 70683
rect 84851 70603 84862 70667
rect 84926 70603 84937 70667
rect 84851 70587 84937 70603
rect 84851 70523 84862 70587
rect 84926 70523 84937 70587
rect 84851 70507 84937 70523
rect 84851 70443 84862 70507
rect 84926 70443 84937 70507
rect 84851 70427 84937 70443
rect 84851 70363 84862 70427
rect 84926 70363 84937 70427
rect 84851 70347 84937 70363
rect 84851 70283 84862 70347
rect 84926 70283 84937 70347
rect 84851 70267 84937 70283
rect 84851 70203 84862 70267
rect 84926 70203 84937 70267
rect 84851 70183 84937 70203
rect 85939 70747 86025 70767
rect 85939 70683 85950 70747
rect 86014 70683 86025 70747
rect 85939 70667 86025 70683
rect 85939 70603 85950 70667
rect 86014 70603 86025 70667
rect 85939 70587 86025 70603
rect 85939 70523 85950 70587
rect 86014 70523 86025 70587
rect 85939 70507 86025 70523
rect 85939 70443 85950 70507
rect 86014 70443 86025 70507
rect 85939 70427 86025 70443
rect 85939 70363 85950 70427
rect 86014 70363 86025 70427
rect 85939 70347 86025 70363
rect 85939 70283 85950 70347
rect 86014 70283 86025 70347
rect 85939 70267 86025 70283
rect 85939 70203 85950 70267
rect 86014 70203 86025 70267
rect 85939 70183 86025 70203
rect 87027 70747 87113 70767
rect 87027 70683 87038 70747
rect 87102 70683 87113 70747
rect 87027 70667 87113 70683
rect 87027 70603 87038 70667
rect 87102 70603 87113 70667
rect 87027 70587 87113 70603
rect 87027 70523 87038 70587
rect 87102 70523 87113 70587
rect 87027 70507 87113 70523
rect 87027 70443 87038 70507
rect 87102 70443 87113 70507
rect 87027 70427 87113 70443
rect 87027 70363 87038 70427
rect 87102 70363 87113 70427
rect 87027 70347 87113 70363
rect 87027 70283 87038 70347
rect 87102 70283 87113 70347
rect 87027 70267 87113 70283
rect 87027 70203 87038 70267
rect 87102 70203 87113 70267
rect 87027 70183 87113 70203
rect 88115 70747 88201 70767
rect 88115 70683 88126 70747
rect 88190 70683 88201 70747
rect 88115 70667 88201 70683
rect 88115 70603 88126 70667
rect 88190 70603 88201 70667
rect 88115 70587 88201 70603
rect 88115 70523 88126 70587
rect 88190 70523 88201 70587
rect 88115 70507 88201 70523
rect 88115 70443 88126 70507
rect 88190 70443 88201 70507
rect 109850 70486 110086 79123
rect 88115 70427 88201 70443
rect 88115 70363 88126 70427
rect 88190 70363 88201 70427
rect 88115 70347 88201 70363
rect 88115 70283 88126 70347
rect 88190 70283 88201 70347
rect 97673 70397 97757 70402
rect 104863 70397 110086 70486
rect 97673 70393 110086 70397
rect 97673 70337 97687 70393
rect 97743 70337 110086 70393
rect 97673 70333 110086 70337
rect 97673 70328 97757 70333
rect 88115 70267 88201 70283
rect 88115 70203 88126 70267
rect 88190 70203 88201 70267
rect 104863 70250 110086 70333
rect 112280 74908 120001 75144
rect 88115 70183 88201 70203
rect 67264 70131 67655 70155
rect 57428 69855 57662 69871
rect 57428 68351 57473 69855
rect 57617 68351 57662 69855
rect 57428 68335 57662 68351
rect 57436 65393 57616 65410
rect 51343 63876 51443 63939
rect 51127 63873 51443 63876
rect 57436 63889 57454 65393
rect 57598 63889 57616 65393
rect 51127 63850 56956 63873
rect 57436 63872 57616 63889
rect 67264 63907 67307 70131
rect 67611 63907 67655 70131
rect 112280 69924 112516 74908
rect 98230 69841 98314 69846
rect 104863 69841 112516 69924
rect 98230 69837 112516 69841
rect 75315 69770 75433 69796
rect 75315 69706 75339 69770
rect 75403 69706 75433 69770
rect 75315 69681 75433 69706
rect 75860 69770 75978 69795
rect 75860 69706 75885 69770
rect 75949 69706 75978 69770
rect 75860 69680 75978 69706
rect 76402 69761 76520 69791
rect 76402 69697 76431 69761
rect 76495 69697 76520 69761
rect 76402 69676 76520 69697
rect 76950 69760 77068 69789
rect 76950 69696 76976 69760
rect 77040 69696 77068 69760
rect 76950 69674 77068 69696
rect 78580 69748 78692 69773
rect 78580 69684 78607 69748
rect 78671 69684 78692 69748
rect 78580 69659 78692 69684
rect 79127 69745 79236 69764
rect 79127 69681 79150 69745
rect 79214 69681 79236 69745
rect 79127 69659 79236 69681
rect 79669 69744 79790 69767
rect 79669 69680 79692 69744
rect 79756 69680 79790 69744
rect 79669 69655 79790 69680
rect 80208 69749 80331 69772
rect 80208 69685 80239 69749
rect 80303 69685 80331 69749
rect 80208 69656 80331 69685
rect 82931 69760 83049 69788
rect 82931 69696 82957 69760
rect 83021 69696 83049 69760
rect 82931 69673 83049 69696
rect 83475 69764 83593 69788
rect 83475 69700 83500 69764
rect 83564 69700 83593 69764
rect 83475 69673 83593 69700
rect 84014 69758 84132 69786
rect 84014 69694 84042 69758
rect 84106 69694 84132 69758
rect 84014 69671 84132 69694
rect 84573 69749 84691 69775
rect 84573 69685 84599 69749
rect 84663 69685 84691 69749
rect 84573 69660 84691 69685
rect 86197 69760 86315 69787
rect 86197 69696 86223 69760
rect 86287 69696 86315 69760
rect 86197 69672 86315 69696
rect 86739 69753 86857 69778
rect 86739 69689 86767 69753
rect 86831 69689 86857 69753
rect 86739 69663 86857 69689
rect 87292 69757 87410 69782
rect 87292 69693 87317 69757
rect 87381 69693 87410 69757
rect 87292 69667 87410 69693
rect 87822 69757 87940 69784
rect 98230 69781 98244 69837
rect 98300 69781 112516 69837
rect 98230 69777 112516 69781
rect 98230 69772 98314 69777
rect 87822 69693 87850 69757
rect 87914 69693 87940 69757
rect 87822 69669 87940 69693
rect 104863 69688 112516 69777
rect 114815 71169 120001 71405
rect 101838 69094 102410 69101
rect 75856 69030 75885 69094
rect 75949 69030 96869 69094
rect 96805 69013 96869 69030
rect 101838 69030 101852 69094
rect 101916 69030 101932 69094
rect 101996 69030 102012 69094
rect 102076 69030 102092 69094
rect 102156 69030 102172 69094
rect 102236 69030 102252 69094
rect 102316 69030 102332 69094
rect 102396 69030 102410 69094
rect 101838 69024 102410 69030
rect 98072 69013 98156 69018
rect 96805 69009 98156 69013
rect 96805 68953 98086 69009
rect 98142 68953 98156 69009
rect 96805 68949 98156 68953
rect 98072 68944 98156 68949
rect 103378 68961 103634 68966
rect 114815 68961 115051 71169
rect 103378 68951 115051 68961
rect 96641 68913 96725 68918
rect 82938 68849 82957 68913
rect 83021 68909 96725 68913
rect 83021 68853 96655 68909
rect 96711 68853 96725 68909
rect 83021 68849 96725 68853
rect 96641 68844 96725 68849
rect 103378 68735 103398 68951
rect 103614 68735 115051 68951
rect 96641 68723 96725 68728
rect 75325 68659 75339 68723
rect 75403 68719 96725 68723
rect 103378 68725 115051 68735
rect 103378 68720 103634 68725
rect 75403 68663 96655 68719
rect 96711 68663 96725 68719
rect 75403 68659 96725 68663
rect 96641 68654 96725 68659
rect 97972 68629 98056 68634
rect 96805 68625 98056 68629
rect 96805 68569 97986 68625
rect 98042 68569 98056 68625
rect 96805 68565 98056 68569
rect 96805 68548 96869 68565
rect 97972 68560 98056 68565
rect 83486 68484 83500 68548
rect 83564 68484 96869 68548
rect 98600 68548 98978 68554
rect 98600 68484 98637 68548
rect 98701 68484 98717 68548
rect 98781 68484 98797 68548
rect 98861 68484 98877 68548
rect 98941 68484 98978 68548
rect 98600 68479 98978 68484
rect 79681 67880 79691 67944
rect 79755 67880 96869 67944
rect 96805 67863 96869 67880
rect 101850 67943 102397 67952
rect 101850 67879 101891 67943
rect 101955 67879 101971 67943
rect 102035 67879 102051 67943
rect 102115 67879 102131 67943
rect 102195 67879 102211 67943
rect 102275 67879 102291 67943
rect 102355 67879 102397 67943
rect 101850 67871 102397 67879
rect 98072 67863 98156 67868
rect 96805 67859 98156 67863
rect 96805 67803 98086 67859
rect 98142 67803 98156 67859
rect 96805 67799 98156 67803
rect 98072 67794 98156 67799
rect 103366 67810 103622 67815
rect 103366 67800 120001 67810
rect 96641 67763 96725 67768
rect 87840 67699 87850 67763
rect 87914 67759 96725 67763
rect 87914 67703 96655 67759
rect 96711 67703 96725 67759
rect 87914 67699 96725 67703
rect 96641 67694 96725 67699
rect 103366 67584 103386 67800
rect 103602 67584 120001 67800
rect 96641 67573 96725 67578
rect 80229 67509 80239 67573
rect 80303 67569 96725 67573
rect 103366 67574 120001 67584
rect 103366 67569 103622 67574
rect 80303 67513 96655 67569
rect 96711 67513 96725 67569
rect 80303 67509 96725 67513
rect 96641 67504 96725 67509
rect 97972 67479 98056 67484
rect 96805 67475 98056 67479
rect 96805 67419 97986 67475
rect 98042 67419 98056 67475
rect 96805 67415 98056 67419
rect 96805 67398 96869 67415
rect 97972 67410 98056 67415
rect 87308 67397 96869 67398
rect 87306 67333 87316 67397
rect 87380 67334 96869 67397
rect 98598 67398 98976 67404
rect 98598 67334 98635 67398
rect 98699 67334 98715 67398
rect 98779 67334 98795 67398
rect 98859 67334 98875 67398
rect 98939 67334 98976 67398
rect 87380 67333 87390 67334
rect 98598 67329 98976 67334
rect 97673 66707 97757 66712
rect 104854 66707 115059 66799
rect 97673 66703 115059 66707
rect 97673 66647 97687 66703
rect 97743 66647 115059 66703
rect 97673 66643 115059 66647
rect 97673 66638 97757 66643
rect 104854 66563 115059 66643
rect 98230 66151 98314 66156
rect 104845 66151 112476 66245
rect 98230 66147 112476 66151
rect 98230 66091 98244 66147
rect 98300 66091 112476 66147
rect 98230 66087 112476 66091
rect 98230 66082 98314 66087
rect 104845 66009 112476 66087
rect 76966 65340 76976 65404
rect 77040 65340 96869 65404
rect 96805 65323 96869 65340
rect 101840 65401 102387 65410
rect 101840 65337 101881 65401
rect 101945 65337 101961 65401
rect 102025 65337 102041 65401
rect 102105 65337 102121 65401
rect 102185 65337 102201 65401
rect 102265 65337 102281 65401
rect 102345 65337 102387 65401
rect 101840 65329 102387 65337
rect 98072 65323 98156 65328
rect 96805 65319 98156 65323
rect 96805 65263 98086 65319
rect 98142 65263 98156 65319
rect 96805 65259 98156 65263
rect 98072 65254 98156 65259
rect 103224 65278 103480 65283
rect 103224 65268 110131 65278
rect 96641 65223 96725 65228
rect 84032 65159 84042 65223
rect 84106 65219 96725 65223
rect 84106 65163 96655 65219
rect 96711 65163 96725 65219
rect 84106 65159 96725 65163
rect 96641 65154 96725 65159
rect 103224 65052 103244 65268
rect 103460 65052 110131 65268
rect 103224 65042 110131 65052
rect 96641 65033 96725 65038
rect 103224 65037 103480 65042
rect 76399 64969 76431 65033
rect 76495 65029 96725 65033
rect 76495 64973 96655 65029
rect 96711 64973 96725 65029
rect 76495 64969 96725 64973
rect 96641 64964 96725 64969
rect 97972 64939 98056 64944
rect 96805 64935 98056 64939
rect 96805 64879 97986 64935
rect 98042 64879 98056 64935
rect 96805 64875 98056 64879
rect 96805 64858 96869 64875
rect 97972 64870 98056 64875
rect 84584 64794 84599 64858
rect 84663 64794 96869 64858
rect 98516 64857 98894 64863
rect 98516 64793 98553 64857
rect 98617 64793 98633 64857
rect 98697 64793 98713 64857
rect 98777 64793 98793 64857
rect 98857 64793 98894 64857
rect 98516 64788 98894 64793
rect 78597 64070 78607 64134
rect 78671 64070 96869 64134
rect 96805 64053 96869 64070
rect 101840 64131 102387 64140
rect 101840 64067 101881 64131
rect 101945 64067 101961 64131
rect 102025 64067 102041 64131
rect 102105 64067 102121 64131
rect 102185 64067 102201 64131
rect 102265 64067 102281 64131
rect 102345 64067 102387 64131
rect 101840 64059 102387 64067
rect 98072 64053 98156 64058
rect 96805 64049 98156 64053
rect 96805 63993 98086 64049
rect 98142 63993 98156 64049
rect 96805 63989 98156 63993
rect 98072 63984 98156 63989
rect 103195 63988 103451 63993
rect 103195 63978 107936 63988
rect 96641 63953 96725 63958
rect 67264 63884 67655 63907
rect 86757 63889 86767 63953
rect 86831 63949 96725 63953
rect 86831 63893 96655 63949
rect 96711 63893 96725 63949
rect 86831 63889 96725 63893
rect 96641 63884 96725 63889
rect 51127 63706 51426 63850
rect 56930 63706 56956 63850
rect 96641 63763 96725 63768
rect 51127 63683 56956 63706
rect 79141 63699 79151 63763
rect 79215 63759 96725 63763
rect 79215 63703 96655 63759
rect 96711 63703 96725 63759
rect 103195 63762 103215 63978
rect 103431 63762 107936 63978
rect 103195 63752 107936 63762
rect 103195 63747 103451 63752
rect 79215 63699 96725 63703
rect 96641 63694 96725 63699
rect 51127 63672 51443 63683
rect 97972 63669 98056 63674
rect 96805 63665 98056 63669
rect 96805 63609 97986 63665
rect 98042 63609 98056 63665
rect 96805 63605 98056 63609
rect 96805 63588 96869 63605
rect 97972 63600 98056 63605
rect 38201 63524 38297 63564
rect 86213 63524 86223 63588
rect 86287 63524 96869 63588
rect 98514 63588 98892 63594
rect 98514 63524 98551 63588
rect 98615 63524 98631 63588
rect 98695 63524 98711 63588
rect 98775 63524 98791 63588
rect 98855 63524 98892 63588
rect 38201 63460 38217 63524
rect 38281 63460 38297 63524
rect 98514 63519 98892 63524
rect 38201 63444 38297 63460
rect 38201 63380 38217 63444
rect 38281 63380 38297 63444
rect 38201 63364 38297 63380
rect 38201 63300 38217 63364
rect 38281 63300 38297 63364
rect 38201 63284 38297 63300
rect 38201 63220 38217 63284
rect 38281 63220 38297 63284
rect 38201 63204 38297 63220
rect 38201 63140 38217 63204
rect 38281 63140 38297 63204
rect 38201 63124 38297 63140
rect 38201 63060 38217 63124
rect 38281 63060 38297 63124
rect 38201 63044 38297 63060
rect 38201 62980 38217 63044
rect 38281 62980 38297 63044
rect 38201 62964 38297 62980
rect 38201 62900 38217 62964
rect 38281 62900 38297 62964
rect 58567 62905 58631 62909
rect 38201 62884 38297 62900
rect 38201 62820 38217 62884
rect 38281 62820 38297 62884
rect 58557 62896 58641 62905
rect 58557 62840 58571 62896
rect 58627 62840 58641 62896
rect 58557 62831 58641 62840
rect 59597 62895 59699 62908
rect 59597 62831 59616 62895
rect 59680 62831 59699 62895
rect 38201 62804 38297 62820
rect 38201 62740 38217 62804
rect 38281 62740 38297 62804
rect 45371 62748 45381 62812
rect 45445 62748 52381 62812
rect 52445 62748 52455 62812
rect 38201 62724 38297 62740
rect 38201 62660 38217 62724
rect 38281 62660 38297 62724
rect 38201 62644 38297 62660
rect 38201 62580 38217 62644
rect 38281 62580 38297 62644
rect 38201 62564 38297 62580
rect 38201 62500 38217 62564
rect 38281 62500 38297 62564
rect 38201 62484 38297 62500
rect 38201 62420 38217 62484
rect 38281 62420 38297 62484
rect 38201 62404 38297 62420
rect 38201 62340 38217 62404
rect 38281 62340 38297 62404
rect 38201 62324 38297 62340
rect 38201 62260 38217 62324
rect 38281 62260 38297 62324
rect 38201 62244 38297 62260
rect 38201 62180 38217 62244
rect 38281 62180 38297 62244
rect 38201 62164 38297 62180
rect 38201 62100 38217 62164
rect 38281 62100 38297 62164
rect 38201 62084 38297 62100
rect 38201 62020 38217 62084
rect 38281 62020 38297 62084
rect 38201 62004 38297 62020
rect 38201 61940 38217 62004
rect 38281 61940 38297 62004
rect 38201 61924 38297 61940
rect 38201 61860 38217 61924
rect 38281 61860 38297 61924
rect 38201 61844 38297 61860
rect 38201 61780 38217 61844
rect 38281 61780 38297 61844
rect 38201 61764 38297 61780
rect 38201 61700 38217 61764
rect 38281 61700 38297 61764
rect 38201 61684 38297 61700
rect 38201 61620 38217 61684
rect 38281 61620 38297 61684
rect 38201 61604 38297 61620
rect 41082 62203 41234 62568
rect 46182 62405 46189 62469
rect 46253 62405 52971 62469
rect 53035 62405 53045 62469
rect 41868 62303 42372 62321
rect 41868 62203 41888 62303
rect 41082 61921 41888 62203
rect 41082 61619 41234 61921
rect 41868 61839 41888 61921
rect 42352 61839 42372 62303
rect 58567 61921 58631 62831
rect 59597 62815 59699 62831
rect 59597 62751 59616 62815
rect 59680 62751 59699 62815
rect 59597 62735 59699 62751
rect 59597 62671 59616 62735
rect 59680 62671 59699 62735
rect 59597 62659 59699 62671
rect 59599 62422 59718 62447
rect 59599 62358 59626 62422
rect 59690 62358 59718 62422
rect 70915 62394 70925 62458
rect 70989 62394 75339 62458
rect 75403 62394 75413 62458
rect 82947 62376 82957 62440
rect 83021 62376 89508 62440
rect 89572 62376 89582 62440
rect 59599 62342 59718 62358
rect 59599 62278 59626 62342
rect 59690 62278 59718 62342
rect 59599 62262 59718 62278
rect 59599 62198 59626 62262
rect 59690 62198 59718 62262
rect 59599 62182 59718 62198
rect 59599 62118 59626 62182
rect 59690 62118 59718 62182
rect 59090 62096 59154 62105
rect 59599 62102 59718 62118
rect 59080 62087 59164 62096
rect 59080 62031 59094 62087
rect 59150 62031 59164 62087
rect 59080 62022 59164 62031
rect 59599 62038 59626 62102
rect 59690 62038 59718 62102
rect 49362 61857 49372 61921
rect 49436 61857 54696 61921
rect 54760 61857 56334 61921
rect 56398 61857 56408 61921
rect 58557 61857 58567 61921
rect 58631 61857 58641 61921
rect 41868 61821 42372 61839
rect 21566 61591 21822 61595
rect 0 61580 21822 61591
rect 0 61364 21586 61580
rect 21802 61364 21822 61580
rect 38201 61540 38217 61604
rect 38281 61540 38297 61604
rect 38201 61524 38297 61540
rect 38201 61460 38217 61524
rect 38281 61460 38297 61524
rect 38201 61444 38297 61460
rect 38201 61380 38217 61444
rect 38281 61380 38297 61444
rect 0 61355 21822 61364
rect 21566 61349 21822 61355
rect 30005 61363 30109 61380
rect 27432 61345 27961 61350
rect 27432 61281 27464 61345
rect 27528 61281 27544 61345
rect 27608 61281 27624 61345
rect 27688 61281 27704 61345
rect 27768 61281 27784 61345
rect 27848 61281 27864 61345
rect 27928 61281 27961 61345
rect 27432 61276 27961 61281
rect 30005 61299 30025 61363
rect 30089 61299 30109 61363
rect 30005 61283 30109 61299
rect 30005 61219 30025 61283
rect 30089 61219 30109 61283
rect 30005 61203 30109 61219
rect 30005 61139 30025 61203
rect 30089 61139 30109 61203
rect 30005 61123 30109 61139
rect 30005 61059 30025 61123
rect 30089 61059 30109 61123
rect 30005 61043 30109 61059
rect 30005 60979 30025 61043
rect 30089 60979 30109 61043
rect 30005 60963 30109 60979
rect 30005 60899 30025 60963
rect 30089 60899 30109 60963
rect 30005 60883 30109 60899
rect 30005 60819 30025 60883
rect 30089 60819 30109 60883
rect 30005 60803 30109 60819
rect 30005 60739 30025 60803
rect 30089 60739 30109 60803
rect 30005 60723 30109 60739
rect 30005 60659 30025 60723
rect 30089 60659 30109 60723
rect 30005 60643 30109 60659
rect 30005 60579 30025 60643
rect 30089 60579 30109 60643
rect 30005 60563 30109 60579
rect 30005 60499 30025 60563
rect 30089 60499 30109 60563
rect 30005 60482 30109 60499
rect 38201 61364 38297 61380
rect 38201 61300 38217 61364
rect 38281 61300 38297 61364
rect 48604 61329 48614 61393
rect 48678 61329 54279 61393
rect 54343 61392 56365 61393
rect 54343 61329 56334 61392
rect 56324 61328 56334 61329
rect 56398 61328 56408 61392
rect 38201 61284 38297 61300
rect 38201 61220 38217 61284
rect 38281 61220 38297 61284
rect 38201 61204 38297 61220
rect 38201 61140 38217 61204
rect 38281 61140 38297 61204
rect 58567 61156 58631 61857
rect 59090 61392 59154 62022
rect 59599 62013 59718 62038
rect 71670 61819 71680 61883
rect 71744 61819 75885 61883
rect 75949 61819 75959 61883
rect 83490 61796 83500 61860
rect 83564 61796 88918 61860
rect 88982 61796 88992 61860
rect 59080 61328 59090 61392
rect 59154 61328 59164 61392
rect 38201 61124 38297 61140
rect 38201 61060 38217 61124
rect 38281 61060 38297 61124
rect 58557 61147 58641 61156
rect 58557 61091 58571 61147
rect 58627 61091 58641 61147
rect 58557 61082 58641 61091
rect 38201 61044 38297 61060
rect 38201 60980 38217 61044
rect 38281 60980 38297 61044
rect 38201 60964 38297 60980
rect 38201 60900 38217 60964
rect 38281 60900 38297 60964
rect 38201 60884 38297 60900
rect 38201 60820 38217 60884
rect 38281 60820 38297 60884
rect 38201 60804 38297 60820
rect 38201 60740 38217 60804
rect 38281 60740 38297 60804
rect 38201 60724 38297 60740
rect 38201 60660 38217 60724
rect 38281 60660 38297 60724
rect 38201 60644 38297 60660
rect 38201 60580 38217 60644
rect 38281 60580 38297 60644
rect 38201 60564 38297 60580
rect 38201 60500 38217 60564
rect 38281 60500 38297 60564
rect 38201 60484 38297 60500
rect 38201 60420 38217 60484
rect 38281 60420 38297 60484
rect 38201 60404 38297 60420
rect 38201 60340 38217 60404
rect 38281 60340 38297 60404
rect 59090 60346 59154 61328
rect 72314 61268 72324 61332
rect 72388 61268 76431 61332
rect 76495 61268 76505 61332
rect 87840 61187 87850 61251
rect 87914 61187 88325 61251
rect 88389 61187 88399 61251
rect 59252 61157 59336 61176
rect 59252 61093 59262 61157
rect 59326 61093 59336 61157
rect 59252 61077 59336 61093
rect 59252 61013 59262 61077
rect 59326 61013 59336 61077
rect 59252 60997 59336 61013
rect 59252 60933 59262 60997
rect 59326 60933 59336 60997
rect 59252 60915 59336 60933
rect 59253 60673 59337 60695
rect 73074 60686 73084 60750
rect 73148 60686 76976 60750
rect 77040 60686 77050 60750
rect 59253 60609 59263 60673
rect 59327 60609 59337 60673
rect 63429 60619 63513 60624
rect 59253 60593 59337 60609
rect 59253 60529 59263 60593
rect 59327 60529 59337 60593
rect 59253 60513 59337 60529
rect 59253 60449 59263 60513
rect 59327 60449 59337 60513
rect 59253 60433 59337 60449
rect 59253 60369 59263 60433
rect 59327 60369 59337 60433
rect 59253 60353 59337 60369
rect 38201 60324 38297 60340
rect 38201 60260 38217 60324
rect 38281 60260 38297 60324
rect 59080 60337 59164 60346
rect 59080 60281 59094 60337
rect 59150 60281 59164 60337
rect 59080 60272 59164 60281
rect 59253 60289 59263 60353
rect 59327 60289 59337 60353
rect 59253 60267 59337 60289
rect 59555 60615 63513 60619
rect 59555 60559 63443 60615
rect 63499 60559 63513 60615
rect 59555 60555 63513 60559
rect 38201 60244 38297 60260
rect 30007 60146 30108 60187
rect 30007 60082 30025 60146
rect 30089 60082 30108 60146
rect 38201 60180 38217 60244
rect 38281 60180 38297 60244
rect 38201 60141 38297 60180
rect 30007 60066 30108 60082
rect 30007 60002 30025 60066
rect 30089 60002 30108 60066
rect 30007 59986 30108 60002
rect 30007 59922 30025 59986
rect 30089 59922 30108 59986
rect 59555 59963 59619 60555
rect 63429 60550 63513 60555
rect 87306 60551 87316 60615
rect 87380 60551 87678 60615
rect 87742 60551 87752 60615
rect 63439 60545 63503 60550
rect 63439 60280 63503 60286
rect 63429 60271 63513 60280
rect 63429 60215 63443 60271
rect 63499 60215 63513 60271
rect 63429 60206 63513 60215
rect 60216 60115 60335 60157
rect 60666 60116 60915 60121
rect 60022 60109 60447 60115
rect 60022 60053 60046 60109
rect 60102 60053 60126 60109
rect 60182 60053 60206 60109
rect 60262 60053 60286 60109
rect 60342 60053 60366 60109
rect 60422 60053 60447 60109
rect 60022 60047 60447 60053
rect 60666 60052 60678 60116
rect 60742 60052 60758 60116
rect 60822 60052 60838 60116
rect 60902 60052 60915 60116
rect 60666 60047 60915 60052
rect 62139 60115 62455 60131
rect 62139 60111 62185 60115
rect 62249 60111 62265 60115
rect 62329 60111 62345 60115
rect 62409 60111 62455 60115
rect 62139 60055 62149 60111
rect 62445 60055 62455 60111
rect 62139 60051 62185 60055
rect 62249 60051 62265 60055
rect 62329 60051 62345 60055
rect 62409 60051 62455 60055
rect 30007 59906 30108 59922
rect 30007 59842 30025 59906
rect 30089 59842 30108 59906
rect 47876 59899 47886 59963
rect 47950 59899 59619 59963
rect 30007 59826 30108 59842
rect 30007 59762 30025 59826
rect 30089 59762 30108 59826
rect 30007 59746 30108 59762
rect 30007 59682 30025 59746
rect 30089 59682 30108 59746
rect 60216 59694 60335 60047
rect 62139 60035 62455 60051
rect 62658 60116 62905 60124
rect 62658 60052 62669 60116
rect 62733 60052 62749 60116
rect 62813 60052 62829 60116
rect 62893 60052 62905 60116
rect 62658 60044 62905 60052
rect 30007 59666 30108 59682
rect 30007 59602 30025 59666
rect 30089 59602 30108 59666
rect 30007 59586 30108 59602
rect 30007 59522 30025 59586
rect 30089 59522 30108 59586
rect 60205 59666 60344 59694
rect 60205 59602 60242 59666
rect 60306 59602 60344 59666
rect 60205 59575 60344 59602
rect 30007 59506 30108 59522
rect 30007 59442 30025 59506
rect 30089 59442 30108 59506
rect 30007 59426 30108 59442
rect 30007 59362 30025 59426
rect 30089 59362 30108 59426
rect 63439 59373 63503 60206
rect 64597 60121 64716 60143
rect 64020 60108 64261 60116
rect 64020 60104 64068 60108
rect 64132 60104 64148 60108
rect 64212 60104 64261 60108
rect 64020 60048 64032 60104
rect 64248 60048 64261 60104
rect 64020 60044 64068 60048
rect 64132 60044 64148 60048
rect 64212 60044 64261 60048
rect 64467 60111 64785 60121
rect 64467 60055 64478 60111
rect 64534 60055 64558 60111
rect 64614 60055 64638 60111
rect 64694 60055 64718 60111
rect 64774 60055 64785 60111
rect 64467 60045 64785 60055
rect 66005 60110 66452 60120
rect 66005 60054 66040 60110
rect 66096 60054 66120 60110
rect 66176 60054 66200 60110
rect 66256 60054 66280 60110
rect 66336 60054 66360 60110
rect 66416 60054 66452 60110
rect 66005 60045 66452 60054
rect 66659 60111 66906 60118
rect 66659 60047 66670 60111
rect 66734 60047 66750 60111
rect 66814 60047 66830 60111
rect 66894 60047 66906 60111
rect 64020 60037 64261 60044
rect 64597 59663 64716 60045
rect 66164 59672 66283 60045
rect 66659 60040 66906 60047
rect 73805 60008 73815 60072
rect 73879 60008 80239 60072
rect 80303 60008 80313 60072
rect 86757 59928 86767 59992
rect 86831 59928 87084 59992
rect 87148 59928 87158 59992
rect 64587 59635 64726 59663
rect 64587 59571 64624 59635
rect 64688 59571 64726 59635
rect 64587 59544 64726 59571
rect 66154 59644 66293 59672
rect 66154 59580 66191 59644
rect 66255 59580 66293 59644
rect 66154 59553 66293 59580
rect 30007 59346 30108 59362
rect 30007 59282 30025 59346
rect 30089 59282 30108 59346
rect 47015 59309 47025 59373
rect 47089 59309 63503 59373
rect 74496 59301 74506 59365
rect 74570 59301 79692 59365
rect 79756 59301 79766 59365
rect 30007 59266 30108 59282
rect 30007 59202 30025 59266
rect 30089 59202 30108 59266
rect 86213 59216 86223 59280
rect 86287 59216 86501 59280
rect 86565 59216 86575 59280
rect 30007 59186 30108 59202
rect 30007 59122 30025 59186
rect 30089 59122 30108 59186
rect 30007 59106 30108 59122
rect 30007 59042 30025 59106
rect 30089 59042 30108 59106
rect 30007 59002 30108 59042
rect 30005 58708 30104 58718
rect 30005 58644 30022 58708
rect 30086 58644 30104 58708
rect 47715 58698 47799 58703
rect 30005 58628 30104 58644
rect 43689 58634 43699 58698
rect 43763 58694 47799 58698
rect 43763 58638 47729 58694
rect 47785 58638 47799 58694
rect 43763 58634 47799 58638
rect 47715 58629 47799 58634
rect 30005 58564 30022 58628
rect 30086 58564 30104 58628
rect 30005 58548 30104 58564
rect 30005 58484 30022 58548
rect 30086 58484 30104 58548
rect 75336 58541 75346 58605
rect 75410 58541 79150 58605
rect 79214 58541 79224 58605
rect 30005 58468 30104 58484
rect 84032 58480 84042 58544
rect 84106 58480 85922 58544
rect 85986 58480 85996 58544
rect 30005 58404 30022 58468
rect 30086 58404 30104 58468
rect 30005 58388 30104 58404
rect 30005 58324 30022 58388
rect 30086 58324 30104 58388
rect 30005 58308 30104 58324
rect 30005 58244 30022 58308
rect 30086 58244 30104 58308
rect 30005 58228 30104 58244
rect 30005 58164 30022 58228
rect 30086 58164 30104 58228
rect 63016 58217 63100 58222
rect 30005 58148 30104 58164
rect 52371 58153 52381 58217
rect 52445 58213 63100 58217
rect 52445 58157 63030 58213
rect 63086 58157 63100 58213
rect 52445 58153 63100 58157
rect 63016 58148 63100 58153
rect 30005 58084 30022 58148
rect 30086 58084 30104 58148
rect 30005 58068 30104 58084
rect 30005 58004 30022 58068
rect 30086 58004 30104 58068
rect 30005 57988 30104 58004
rect 30005 57924 30022 57988
rect 30086 57924 30104 57988
rect 30005 57908 30104 57924
rect 30005 57844 30022 57908
rect 30086 57844 30104 57908
rect 63822 57872 63906 57877
rect 30005 57828 30104 57844
rect 30005 57764 30022 57828
rect 30086 57764 30104 57828
rect 52961 57808 52971 57872
rect 53035 57868 63906 57872
rect 53035 57812 63836 57868
rect 63892 57812 63906 57868
rect 53035 57808 63906 57812
rect 63822 57803 63906 57808
rect 84589 57771 84599 57835
rect 84663 57771 85409 57835
rect 85473 57771 85483 57835
rect 30005 57748 30104 57764
rect 30005 57684 30022 57748
rect 30086 57684 30104 57748
rect 76339 57704 76349 57768
rect 76413 57704 78607 57768
rect 78671 57704 78682 57768
rect 30005 57668 30104 57684
rect 30005 57604 30022 57668
rect 30086 57604 30104 57668
rect 30005 57588 30104 57604
rect 30005 57524 30022 57588
rect 30086 57524 30104 57588
rect 30005 57515 30104 57524
rect 35554 57573 35660 57597
rect 35554 57509 35576 57573
rect 35640 57509 35660 57573
rect 35554 57488 35660 57509
rect 50136 57201 50220 57206
rect 41945 57137 41955 57201
rect 42019 57197 50220 57201
rect 42019 57141 50150 57197
rect 50206 57141 50220 57197
rect 42019 57137 50220 57141
rect 50136 57132 50220 57137
rect 30000 56886 30099 56926
rect 30000 56822 30017 56886
rect 30081 56822 30099 56886
rect 30000 56806 30099 56822
rect 30000 56742 30017 56806
rect 30081 56742 30099 56806
rect 30000 56726 30099 56742
rect 30000 56662 30017 56726
rect 30081 56662 30099 56726
rect 30000 56646 30099 56662
rect 30000 56582 30017 56646
rect 30081 56582 30099 56646
rect 30000 56566 30099 56582
rect 30000 56502 30017 56566
rect 30081 56502 30099 56566
rect 30000 56486 30099 56502
rect 30000 56422 30017 56486
rect 30081 56422 30099 56486
rect 30000 56382 30099 56422
rect 64448 56374 64532 56379
rect 62401 56367 62485 56372
rect 62215 56363 62485 56367
rect 62215 56307 62415 56363
rect 62471 56307 62485 56363
rect 62215 56303 62485 56307
rect 64448 56370 64701 56374
rect 64448 56314 64462 56370
rect 64518 56314 64701 56370
rect 64448 56310 64701 56314
rect 64448 56305 64532 56310
rect 62401 56298 62485 56303
rect 62058 55474 62122 56195
rect 64796 55474 64860 56195
rect 65036 55833 65147 55863
rect 65036 55769 65059 55833
rect 65123 55769 65147 55833
rect 65036 55745 65147 55769
rect 62058 55397 62122 55410
rect 64796 55397 64860 55410
rect 68431 55349 68441 55413
rect 68505 55349 70925 55413
rect 70989 55349 70999 55413
rect 62796 55213 62860 55214
rect 61038 55145 61836 55209
rect 62035 55149 62860 55213
rect 61055 54411 61119 55145
rect 61419 54454 61534 54482
rect 61419 54390 61448 54454
rect 61512 54390 61534 54454
rect 62796 54416 62860 55149
rect 64058 55213 64122 55214
rect 64058 55149 64883 55213
rect 64058 54416 64122 55149
rect 65082 55145 65880 55209
rect 65394 54459 65509 54486
rect 61419 54364 61534 54390
rect 65394 54395 65422 54459
rect 65486 54395 65509 54459
rect 65799 54411 65863 55145
rect 69050 54730 69060 54794
rect 69124 54730 71680 54794
rect 71744 54730 71754 54794
rect 107700 54491 107936 63752
rect 109895 57654 110131 65042
rect 112240 61116 112476 66009
rect 114823 64424 115059 66563
rect 114823 64188 120001 64424
rect 112240 60880 120001 61116
rect 109895 57418 120001 57654
rect 65394 54370 65509 54395
rect 60392 54327 60512 54357
rect 60392 54263 60420 54327
rect 60484 54263 60512 54327
rect 60392 54234 60512 54263
rect 107700 54255 120001 54491
rect 44391 53774 44475 53779
rect 58997 53774 59081 53779
rect 44391 53770 53176 53774
rect 44391 53714 44405 53770
rect 44461 53714 53176 53770
rect 44391 53710 53176 53714
rect 53240 53770 59081 53774
rect 53240 53714 59011 53770
rect 59067 53714 59081 53770
rect 53240 53710 59081 53714
rect 44391 53705 44475 53710
rect 58997 53705 59081 53710
rect 61055 53411 61119 54209
rect 61422 54004 61703 54068
rect 43615 53351 43699 53356
rect 58997 53351 59081 53356
rect 43615 53347 51815 53351
rect 43615 53291 43629 53347
rect 43685 53291 51815 53347
rect 43615 53287 51815 53291
rect 51879 53347 59081 53351
rect 51879 53291 59011 53347
rect 59067 53291 59081 53347
rect 51879 53287 59081 53291
rect 43615 53282 43699 53287
rect 58997 53282 59081 53287
rect 61055 52411 61119 53209
rect 61422 52622 61486 54004
rect 62796 53416 62860 54214
rect 64058 53416 64122 54214
rect 65215 54004 65496 54068
rect 61795 52835 61859 53034
rect 61785 52826 61869 52835
rect 61785 52770 61799 52826
rect 61855 52770 61869 52826
rect 61785 52761 61869 52770
rect 61412 52615 61496 52622
rect 61412 52613 61673 52615
rect 61412 52557 61426 52613
rect 61482 52557 61673 52613
rect 61412 52551 61673 52557
rect 61412 52548 61496 52551
rect 62796 52416 62860 53214
rect 64058 52416 64122 53214
rect 65054 52873 65118 53043
rect 65044 52864 65128 52873
rect 65044 52808 65058 52864
rect 65114 52808 65128 52864
rect 65044 52799 65128 52808
rect 65432 52619 65496 54004
rect 65799 53411 65863 54209
rect 73786 53774 73905 53803
rect 73786 53710 73815 53774
rect 73879 53710 73905 53774
rect 73786 53681 73905 53710
rect 74472 53351 74600 53388
rect 74472 53287 74506 53351
rect 74570 53287 74600 53351
rect 74472 53254 74600 53287
rect 65422 52615 65506 52619
rect 65245 52610 65506 52615
rect 65245 52554 65436 52610
rect 65492 52554 65506 52610
rect 65245 52551 65506 52554
rect 65422 52545 65506 52551
rect 65799 52411 65863 53209
rect 67717 52762 67727 52826
rect 67791 52762 69060 52826
rect 69124 52762 69134 52826
rect 41372 52085 41491 52125
rect 41372 52021 41399 52085
rect 41463 52021 41491 52085
rect 41372 52005 41491 52021
rect 41372 51941 41399 52005
rect 41463 51941 41491 52005
rect 41372 51925 41491 51941
rect 41372 51861 41399 51925
rect 41463 51861 41491 51925
rect 41372 51845 41491 51861
rect 41372 51781 41399 51845
rect 41463 51781 41491 51845
rect 41372 51765 41491 51781
rect 41372 51701 41399 51765
rect 41463 51701 41491 51765
rect 39449 51634 39597 51671
rect 41372 51662 41491 51701
rect 44695 52087 44788 52103
rect 44695 52023 44709 52087
rect 44773 52023 44788 52087
rect 44695 52007 44788 52023
rect 44695 51943 44709 52007
rect 44773 51943 44788 52007
rect 44695 51927 44788 51943
rect 44695 51863 44709 51927
rect 44773 51863 44788 51927
rect 44695 51847 44788 51863
rect 44695 51783 44709 51847
rect 44773 51783 44788 51847
rect 44695 51767 44788 51783
rect 44695 51703 44709 51767
rect 44773 51703 44788 51767
rect 44695 51687 44788 51703
rect 39449 51570 39491 51634
rect 39555 51570 39597 51634
rect 39449 51533 39597 51570
rect 51785 51554 51908 51587
rect 51785 51490 51815 51554
rect 51879 51490 51908 51554
rect 51785 51462 51908 51490
rect 61055 51473 61119 52209
rect 62796 51473 62860 52214
rect 44690 51446 44807 51454
rect 44690 51382 44716 51446
rect 44780 51382 44807 51446
rect 61055 51411 61858 51473
rect 61060 51409 61858 51411
rect 62060 51416 62860 51473
rect 64058 51473 64122 52214
rect 65799 51473 65863 52209
rect 64058 51416 64858 51473
rect 62060 51409 62858 51416
rect 64060 51409 64858 51416
rect 65060 51411 65863 51473
rect 65060 51409 65858 51411
rect 44690 51366 44807 51382
rect 44690 51302 44716 51366
rect 44780 51302 44807 51366
rect 44690 51286 44807 51302
rect 44690 51222 44716 51286
rect 44780 51222 44807 51286
rect 44690 51215 44807 51222
rect 53146 50877 53269 50911
rect 53146 50813 53176 50877
rect 53240 50813 53269 50877
rect 53146 50786 53269 50813
rect 18894 50616 22248 50638
rect 18894 50552 18939 50616
rect 19003 50552 19019 50616
rect 19083 50552 19099 50616
rect 19163 50552 19179 50616
rect 19243 50552 19259 50616
rect 19323 50552 19339 50616
rect 19403 50552 19419 50616
rect 19483 50552 19499 50616
rect 19563 50552 19579 50616
rect 19643 50552 19659 50616
rect 19723 50552 19739 50616
rect 19803 50552 19819 50616
rect 19883 50552 19899 50616
rect 19963 50552 19979 50616
rect 20043 50552 20059 50616
rect 20123 50552 20139 50616
rect 20203 50552 20219 50616
rect 20283 50552 20299 50616
rect 20363 50552 20379 50616
rect 20443 50552 20459 50616
rect 20523 50552 20539 50616
rect 20603 50552 20619 50616
rect 20683 50552 20699 50616
rect 20763 50552 20779 50616
rect 20843 50552 20859 50616
rect 20923 50552 20939 50616
rect 21003 50552 21019 50616
rect 21083 50552 21099 50616
rect 21163 50552 21179 50616
rect 21243 50552 21259 50616
rect 21323 50552 21339 50616
rect 21403 50552 21419 50616
rect 21483 50552 21499 50616
rect 21563 50552 21579 50616
rect 21643 50552 21659 50616
rect 21723 50552 21739 50616
rect 21803 50552 21819 50616
rect 21883 50552 21899 50616
rect 21963 50552 21979 50616
rect 22043 50552 22059 50616
rect 22123 50552 22139 50616
rect 22203 50552 22248 50616
rect 18894 50531 22248 50552
rect 44688 50485 44803 50513
rect 39449 50405 39597 50442
rect 39449 50341 39491 50405
rect 39555 50341 39597 50405
rect 39449 50304 39597 50341
rect 44688 50421 44713 50485
rect 44777 50421 44803 50485
rect 62060 50424 62124 51222
rect 64794 50424 64858 51222
rect 44688 50405 44803 50421
rect 44688 50341 44713 50405
rect 44777 50341 44803 50405
rect 44688 50325 44803 50341
rect 41359 50296 41468 50308
rect 41359 50232 41381 50296
rect 41445 50232 41468 50296
rect 41359 50216 41468 50232
rect 41359 50152 41381 50216
rect 41445 50152 41468 50216
rect 41359 50136 41468 50152
rect 41359 50072 41381 50136
rect 41445 50072 41468 50136
rect 44688 50261 44713 50325
rect 44777 50261 44803 50325
rect 68431 50308 68441 50372
rect 68505 50308 68931 50372
rect 68995 50308 69005 50372
rect 44688 50245 44803 50261
rect 44688 50181 44713 50245
rect 44777 50181 44803 50245
rect 44688 50165 44803 50181
rect 44688 50101 44713 50165
rect 44777 50101 44803 50165
rect 44688 50074 44803 50101
rect 41359 50061 41468 50072
rect 76955 50031 77039 50036
rect 70934 49967 70944 50031
rect 71008 50027 82973 50031
rect 71008 49971 76969 50027
rect 77025 49971 82973 50027
rect 71008 49967 82973 49971
rect 83037 49967 83044 50031
rect 76955 49962 77039 49967
rect 44700 49843 44783 49850
rect 37996 49821 41589 49826
rect 37996 49597 38010 49821
rect 38234 49597 41589 49821
rect 44700 49787 44713 49843
rect 44769 49787 44783 49843
rect 44700 49763 44783 49787
rect 44700 49707 44713 49763
rect 44769 49707 44783 49763
rect 43095 49686 43179 49691
rect 43095 49682 44550 49686
rect 43095 49626 43109 49682
rect 43165 49626 44550 49682
rect 43095 49622 44550 49626
rect 43095 49617 43179 49622
rect 37996 49593 41589 49597
rect 38534 49592 38767 49593
rect 31635 49502 31735 49509
rect 31635 49438 31653 49502
rect 31717 49438 31735 49502
rect 31635 49422 31735 49438
rect 31635 49358 31653 49422
rect 31717 49358 31735 49422
rect 31635 49342 31735 49358
rect 31635 49278 31653 49342
rect 31717 49278 31735 49342
rect 31635 49262 31735 49278
rect 31635 49198 31653 49262
rect 31717 49198 31735 49262
rect 16491 49193 16747 49198
rect 0 49183 16747 49193
rect 31635 49192 31735 49198
rect 41356 49442 41589 49593
rect 41356 49386 41386 49442
rect 41442 49386 41589 49442
rect 41356 49362 41589 49386
rect 44486 49441 44550 49622
rect 44700 49683 44783 49707
rect 44700 49627 44713 49683
rect 44769 49627 44783 49683
rect 44700 49621 44783 49627
rect 44917 49622 45770 49686
rect 45834 49622 45844 49686
rect 44917 49441 44981 49622
rect 76957 49620 77041 49625
rect 70350 49556 70360 49620
rect 70424 49616 83557 49620
rect 70424 49560 76971 49616
rect 77027 49560 83557 49616
rect 70424 49556 83557 49560
rect 83621 49556 83631 49620
rect 76957 49551 77041 49556
rect 44486 49377 44981 49441
rect 41356 49306 41386 49362
rect 41442 49306 41589 49362
rect 41356 49282 41589 49306
rect 41356 49226 41386 49282
rect 41442 49226 41589 49282
rect 41356 49202 41589 49226
rect 0 48967 16511 49183
rect 16727 48967 16747 49183
rect 41356 49146 41386 49202
rect 41442 49146 41589 49202
rect 41356 49122 41589 49146
rect 41356 49066 41386 49122
rect 41442 49066 41589 49122
rect 41356 49033 41589 49066
rect 39449 48992 39597 49029
rect 0 48957 16747 48967
rect 16491 48952 16747 48957
rect 31632 48963 31739 48972
rect 31632 48899 31653 48963
rect 31717 48899 31739 48963
rect 31632 48883 31739 48899
rect 39449 48928 39491 48992
rect 39555 48928 39597 48992
rect 39449 48891 39597 48928
rect 42674 48894 42758 48899
rect 31632 48819 31653 48883
rect 31717 48819 31739 48883
rect 42674 48890 45117 48894
rect 42674 48834 42688 48890
rect 42744 48834 45117 48890
rect 42674 48830 45117 48834
rect 45181 48830 45191 48894
rect 42674 48825 42758 48830
rect 31632 48803 31739 48819
rect 64685 48806 64695 48870
rect 64759 48806 72324 48870
rect 72388 48806 72398 48870
rect 31632 48739 31653 48803
rect 31717 48739 31739 48803
rect 31632 48731 31739 48739
rect 44691 48719 44776 48739
rect 44691 48655 44701 48719
rect 44765 48655 44776 48719
rect 44691 48639 44776 48655
rect 44691 48575 44701 48639
rect 44765 48575 44776 48639
rect 44691 48559 44776 48575
rect 44691 48495 44701 48559
rect 44765 48495 44776 48559
rect 44691 48475 44776 48495
rect 62799 48604 62887 48621
rect 62799 48540 62811 48604
rect 62875 48540 62887 48604
rect 64152 48614 64236 48619
rect 64350 48614 64360 48615
rect 64152 48610 64360 48614
rect 64152 48554 64166 48610
rect 64222 48554 64360 48610
rect 64152 48551 64360 48554
rect 64424 48551 64434 48615
rect 64152 48550 64384 48551
rect 64152 48545 64236 48550
rect 62799 48524 62887 48540
rect 62799 48460 62811 48524
rect 62875 48460 62887 48524
rect 65213 48488 65223 48552
rect 65287 48488 73084 48552
rect 73148 48488 73158 48552
rect 62799 48444 62887 48460
rect 62799 48380 62811 48444
rect 62875 48380 62887 48444
rect 62799 48364 62887 48380
rect 62799 48300 62811 48364
rect 62875 48300 62887 48364
rect 62799 48284 62887 48300
rect 44686 48255 44788 48266
rect 44686 48191 44705 48255
rect 44769 48191 44788 48255
rect 62799 48220 62811 48284
rect 62875 48220 62887 48284
rect 62799 48203 62887 48220
rect 44686 48175 44788 48191
rect 44686 48111 44705 48175
rect 44769 48111 44788 48175
rect 68167 48160 68174 48224
rect 68238 48160 77023 48224
rect 44686 48095 44788 48111
rect 44686 48031 44705 48095
rect 44769 48031 44788 48095
rect 44686 48020 44788 48031
rect 45760 47845 45770 47909
rect 45834 47845 64360 47909
rect 64424 47845 76349 47909
rect 76413 47845 76423 47909
rect 39449 47763 39597 47800
rect 39449 47699 39491 47763
rect 39555 47699 39597 47763
rect 39449 47662 39597 47699
rect 64175 47670 64259 47679
rect 41359 47655 41446 47664
rect 18902 47608 22252 47632
rect 18902 47544 18945 47608
rect 19009 47544 19025 47608
rect 19089 47544 19105 47608
rect 19169 47544 19185 47608
rect 19249 47544 19265 47608
rect 19329 47544 19345 47608
rect 19409 47544 19425 47608
rect 19489 47544 19505 47608
rect 19569 47544 19585 47608
rect 19649 47544 19665 47608
rect 19729 47544 19745 47608
rect 19809 47544 19825 47608
rect 19889 47544 19905 47608
rect 19969 47544 19985 47608
rect 20049 47544 20065 47608
rect 20129 47544 20145 47608
rect 20209 47544 20225 47608
rect 20289 47544 20305 47608
rect 20369 47544 20385 47608
rect 20449 47544 20465 47608
rect 20529 47544 20545 47608
rect 20609 47544 20625 47608
rect 20689 47544 20705 47608
rect 20769 47544 20785 47608
rect 20849 47544 20865 47608
rect 20929 47544 20945 47608
rect 21009 47544 21025 47608
rect 21089 47544 21105 47608
rect 21169 47544 21185 47608
rect 21249 47544 21265 47608
rect 21329 47544 21345 47608
rect 21409 47544 21425 47608
rect 21489 47544 21505 47608
rect 21569 47544 21585 47608
rect 21649 47544 21665 47608
rect 21729 47544 21745 47608
rect 21809 47544 21825 47608
rect 21889 47544 21905 47608
rect 21969 47544 21985 47608
rect 22049 47544 22065 47608
rect 22129 47544 22145 47608
rect 22209 47544 22252 47608
rect 18902 47520 22252 47544
rect 41359 47591 41370 47655
rect 41434 47591 41446 47655
rect 64175 47614 64189 47670
rect 64245 47614 64259 47670
rect 64175 47605 64259 47614
rect 41359 47575 41446 47591
rect 41359 47511 41370 47575
rect 41434 47511 41446 47575
rect 64185 47540 64249 47605
rect 41359 47495 41446 47511
rect 41359 47431 41370 47495
rect 41434 47431 41446 47495
rect 45107 47476 45117 47540
rect 45181 47476 75346 47540
rect 75410 47476 75420 47540
rect 41359 47422 41446 47431
rect 65871 47355 66047 47383
rect 44695 47281 44785 47304
rect 44695 47217 44708 47281
rect 44772 47217 44785 47281
rect 65871 47291 65887 47355
rect 65951 47291 65967 47355
rect 66031 47291 66047 47355
rect 65871 47263 66047 47291
rect 76959 47232 77023 48160
rect 99940 48173 103294 48201
rect 99940 48109 99985 48173
rect 100049 48109 100065 48173
rect 100129 48109 100145 48173
rect 100209 48109 100225 48173
rect 100289 48109 100305 48173
rect 100369 48109 100385 48173
rect 100449 48109 100465 48173
rect 100529 48109 100545 48173
rect 100609 48109 100625 48173
rect 100689 48109 100705 48173
rect 100769 48109 100785 48173
rect 100849 48109 100865 48173
rect 100929 48109 100945 48173
rect 101009 48109 101025 48173
rect 101089 48109 101105 48173
rect 101169 48109 101185 48173
rect 101249 48109 101265 48173
rect 101329 48109 101345 48173
rect 101409 48109 101425 48173
rect 101489 48109 101505 48173
rect 101569 48109 101585 48173
rect 101649 48109 101665 48173
rect 101729 48109 101745 48173
rect 101809 48109 101825 48173
rect 101889 48109 101905 48173
rect 101969 48109 101985 48173
rect 102049 48109 102065 48173
rect 102129 48109 102145 48173
rect 102209 48109 102225 48173
rect 102289 48109 102305 48173
rect 102369 48109 102385 48173
rect 102449 48109 102465 48173
rect 102529 48109 102545 48173
rect 102609 48109 102625 48173
rect 102689 48109 102705 48173
rect 102769 48109 102785 48173
rect 102849 48109 102865 48173
rect 102929 48109 102945 48173
rect 103009 48109 103025 48173
rect 103089 48109 103105 48173
rect 103169 48109 103185 48173
rect 103249 48109 103294 48173
rect 99940 48082 103294 48109
rect 93139 48040 93242 48060
rect 93139 47976 93160 48040
rect 93224 47976 93242 48040
rect 93139 47956 93242 47976
rect 92220 47888 92335 47915
rect 92220 47824 92246 47888
rect 92310 47824 92335 47888
rect 92220 47794 92335 47824
rect 96430 47733 96524 47741
rect 96430 47697 96449 47733
rect 96505 47697 96524 47733
rect 94903 47605 94996 47638
rect 94903 47541 94917 47605
rect 94981 47541 94996 47605
rect 94903 47509 94996 47541
rect 96430 47633 96445 47697
rect 96509 47633 96524 47697
rect 96430 47617 96449 47633
rect 96505 47617 96524 47633
rect 96430 47553 96445 47617
rect 96509 47553 96524 47617
rect 96430 47517 96449 47553
rect 96505 47517 96524 47553
rect 96430 47510 96524 47517
rect 44695 47201 44785 47217
rect 44695 47137 44708 47201
rect 44772 47137 44785 47201
rect 44695 47121 44785 47137
rect 44695 47057 44708 47121
rect 44772 47057 44785 47121
rect 61864 47173 62347 47181
rect 44695 47041 44785 47057
rect 44695 46977 44708 47041
rect 44772 46977 44785 47041
rect 59634 47085 59718 47090
rect 61864 47085 61913 47173
rect 59634 47081 61913 47085
rect 59634 47025 59648 47081
rect 59704 47025 61913 47081
rect 59634 47021 61913 47025
rect 59634 47016 59718 47021
rect 44695 46961 44785 46977
rect 44695 46897 44708 46961
rect 44772 46897 44785 46961
rect 61864 46949 61913 47021
rect 62297 47085 62347 47173
rect 69672 47168 69682 47232
rect 69746 47168 84205 47232
rect 84269 47168 84280 47232
rect 94903 47204 95009 47221
rect 94903 47140 94924 47204
rect 94988 47140 95009 47204
rect 94903 47124 95009 47140
rect 67286 47085 67370 47090
rect 62297 47021 62812 47085
rect 62876 47081 67370 47085
rect 62876 47025 67300 47081
rect 67356 47025 67370 47081
rect 62876 47021 67370 47025
rect 62297 46949 62347 47021
rect 67286 47016 67370 47021
rect 94903 47060 94924 47124
rect 94988 47060 95009 47124
rect 94903 47044 95009 47060
rect 61864 46941 62347 46949
rect 68930 46938 68994 47001
rect 94903 46980 94924 47044
rect 94988 46980 95009 47044
rect 94903 46963 95009 46980
rect 96419 47210 96525 47227
rect 96419 47146 96440 47210
rect 96504 47146 96525 47210
rect 96419 47130 96525 47146
rect 96419 47066 96440 47130
rect 96504 47066 96525 47130
rect 96419 47050 96525 47066
rect 96419 46986 96440 47050
rect 96504 46986 96525 47050
rect 96419 46969 96525 46986
rect 68921 46937 68931 46938
rect 44695 46874 44785 46897
rect 68560 46873 68570 46937
rect 68634 46874 68931 46937
rect 68995 46937 69005 46938
rect 68995 46874 71683 46937
rect 68634 46873 71683 46874
rect 44332 46746 45007 46799
rect 40485 46682 40495 46746
rect 40559 46735 65223 46746
rect 40559 46682 44407 46735
rect 44943 46682 65223 46735
rect 65287 46682 65297 46746
rect 44693 46645 44781 46651
rect 44693 46581 44705 46645
rect 44769 46581 44781 46645
rect 44693 46565 44781 46581
rect 44693 46501 44705 46565
rect 44769 46501 44781 46565
rect 44693 46485 44781 46501
rect 44693 46421 44705 46485
rect 44769 46421 44781 46485
rect 44693 46416 44781 46421
rect 40048 46231 64695 46295
rect 64759 46231 64769 46295
rect 40048 45119 40112 46231
rect 71619 46113 71683 46873
rect 72575 46873 73494 46937
rect 72575 46113 72639 46873
rect 71619 46049 72639 46113
rect 73430 46106 73494 46873
rect 74499 46873 75483 46937
rect 74499 46106 74563 46873
rect 75419 46515 75483 46873
rect 75994 46873 77024 46937
rect 75994 46515 76058 46873
rect 75419 46451 76058 46515
rect 73430 46042 74563 46106
rect 76960 45677 77024 46873
rect 93998 46831 94260 46837
rect 92184 46812 92384 46817
rect 93998 46812 94017 46831
rect 92184 46790 94017 46812
rect 92184 46654 92216 46790
rect 92352 46749 94017 46790
rect 92352 46693 92876 46749
rect 92932 46693 92956 46749
rect 93012 46693 93036 46749
rect 93092 46693 94017 46749
rect 92352 46654 94017 46693
rect 92184 46632 94017 46654
rect 92184 46627 92384 46632
rect 93998 46607 94017 46632
rect 94241 46607 94260 46831
rect 93998 46601 94260 46607
rect 104640 46756 104896 46761
rect 104640 46746 120001 46756
rect 104640 46530 104660 46746
rect 104876 46530 120001 46746
rect 104640 46520 120001 46530
rect 104640 46515 104896 46520
rect 96430 46407 96524 46415
rect 96430 46371 96449 46407
rect 96505 46371 96524 46407
rect 96430 46307 96445 46371
rect 96509 46307 96524 46371
rect 94910 46269 95000 46307
rect 94910 46205 94923 46269
rect 94987 46205 95000 46269
rect 94910 46168 95000 46205
rect 96430 46291 96449 46307
rect 96505 46291 96524 46307
rect 96430 46227 96445 46291
rect 96509 46227 96524 46291
rect 96430 46191 96449 46227
rect 96505 46191 96524 46227
rect 96430 46184 96524 46191
rect 94898 45816 95003 45850
rect 94898 45752 94918 45816
rect 94982 45752 95003 45816
rect 94898 45736 95003 45752
rect 56113 45647 56197 45652
rect 63391 45647 63475 45652
rect 56113 45643 63475 45647
rect 56113 45587 56127 45643
rect 56183 45587 63405 45643
rect 63461 45587 63475 45643
rect 69156 45613 69166 45677
rect 69230 45613 84751 45677
rect 84815 45613 84825 45677
rect 94898 45672 94918 45736
rect 94982 45672 95003 45736
rect 94898 45638 95003 45672
rect 96425 45844 96531 45861
rect 96425 45780 96446 45844
rect 96510 45780 96531 45844
rect 96425 45764 96531 45780
rect 96425 45700 96446 45764
rect 96510 45700 96531 45764
rect 96425 45684 96531 45700
rect 56113 45583 63475 45587
rect 56113 45578 56197 45583
rect 63391 45578 63475 45583
rect 92220 45607 92338 45637
rect 92220 45543 92246 45607
rect 92310 45543 92338 45607
rect 96425 45620 96446 45684
rect 96510 45620 96531 45684
rect 96425 45603 96531 45620
rect 92220 45510 92338 45543
rect 92551 45401 92658 45424
rect 92551 45337 92571 45401
rect 92635 45337 92658 45401
rect 92551 45315 92658 45337
rect 99938 45177 103292 45205
rect 29174 45055 63468 45119
rect 99938 45113 99983 45177
rect 100047 45113 100063 45177
rect 100127 45113 100143 45177
rect 100207 45113 100223 45177
rect 100287 45113 100303 45177
rect 100367 45113 100383 45177
rect 100447 45113 100463 45177
rect 100527 45113 100543 45177
rect 100607 45113 100623 45177
rect 100687 45113 100703 45177
rect 100767 45113 100783 45177
rect 100847 45113 100863 45177
rect 100927 45113 100943 45177
rect 101007 45113 101023 45177
rect 101087 45113 101103 45177
rect 101167 45113 101183 45177
rect 101247 45113 101263 45177
rect 101327 45113 101343 45177
rect 101407 45113 101423 45177
rect 101487 45113 101503 45177
rect 101567 45113 101583 45177
rect 101647 45113 101663 45177
rect 101727 45113 101743 45177
rect 101807 45113 101823 45177
rect 101887 45113 101903 45177
rect 101967 45113 101983 45177
rect 102047 45113 102063 45177
rect 102127 45113 102143 45177
rect 102207 45113 102223 45177
rect 102287 45113 102303 45177
rect 102367 45113 102383 45177
rect 102447 45113 102463 45177
rect 102527 45113 102543 45177
rect 102607 45113 102623 45177
rect 102687 45113 102703 45177
rect 102767 45113 102783 45177
rect 102847 45113 102863 45177
rect 102927 45113 102943 45177
rect 103007 45113 103023 45177
rect 103087 45113 103103 45177
rect 103167 45113 103183 45177
rect 103247 45113 103292 45177
rect 99938 45086 103292 45113
rect 18916 43080 22243 43092
rect 18916 43016 18947 43080
rect 19011 43016 19027 43080
rect 19091 43016 19107 43080
rect 19171 43016 19187 43080
rect 19251 43016 19267 43080
rect 19331 43016 19347 43080
rect 19411 43016 19427 43080
rect 19491 43016 19507 43080
rect 19571 43016 19587 43080
rect 19651 43016 19667 43080
rect 19731 43016 19747 43080
rect 19811 43016 19827 43080
rect 19891 43016 19907 43080
rect 19971 43016 19987 43080
rect 20051 43016 20067 43080
rect 20131 43016 20147 43080
rect 20211 43016 20227 43080
rect 20291 43016 20307 43080
rect 20371 43016 20387 43080
rect 20451 43016 20467 43080
rect 20531 43016 20547 43080
rect 20611 43016 20627 43080
rect 20691 43016 20707 43080
rect 20771 43016 20787 43080
rect 20851 43016 20867 43080
rect 20931 43016 20947 43080
rect 21011 43016 21027 43080
rect 21091 43016 21107 43080
rect 21171 43016 21187 43080
rect 21251 43016 21267 43080
rect 21331 43016 21347 43080
rect 21411 43016 21427 43080
rect 21491 43016 21507 43080
rect 21571 43016 21587 43080
rect 21651 43016 21667 43080
rect 21731 43016 21747 43080
rect 21811 43016 21827 43080
rect 21891 43016 21907 43080
rect 21971 43016 21987 43080
rect 22051 43016 22067 43080
rect 22131 43016 22147 43080
rect 22211 43016 22243 43080
rect 18916 43004 22243 43016
rect 16488 41652 16744 41657
rect 0 41642 16744 41652
rect 0 41426 16508 41642
rect 16724 41426 16744 41642
rect 0 41416 16744 41426
rect 16488 41411 16744 41416
rect 18910 40085 22252 40102
rect 18910 40021 18949 40085
rect 19013 40021 19029 40085
rect 19093 40021 19109 40085
rect 19173 40021 19189 40085
rect 19253 40021 19269 40085
rect 19333 40021 19349 40085
rect 19413 40021 19429 40085
rect 19493 40021 19509 40085
rect 19573 40021 19589 40085
rect 19653 40021 19669 40085
rect 19733 40021 19749 40085
rect 19813 40021 19829 40085
rect 19893 40021 19909 40085
rect 19973 40021 19989 40085
rect 20053 40021 20069 40085
rect 20133 40021 20149 40085
rect 20213 40021 20229 40085
rect 20293 40021 20309 40085
rect 20373 40021 20389 40085
rect 20453 40021 20469 40085
rect 20533 40021 20549 40085
rect 20613 40021 20629 40085
rect 20693 40021 20709 40085
rect 20773 40021 20789 40085
rect 20853 40021 20869 40085
rect 20933 40021 20949 40085
rect 21013 40021 21029 40085
rect 21093 40021 21109 40085
rect 21173 40021 21189 40085
rect 21253 40021 21269 40085
rect 21333 40021 21349 40085
rect 21413 40021 21429 40085
rect 21493 40021 21509 40085
rect 21573 40021 21589 40085
rect 21653 40021 21669 40085
rect 21733 40021 21749 40085
rect 21813 40021 21829 40085
rect 21893 40021 21909 40085
rect 21973 40021 21989 40085
rect 22053 40021 22069 40085
rect 22133 40021 22149 40085
rect 22213 40021 22252 40085
rect 18910 40004 22252 40021
rect 29174 39468 29238 45055
rect 63404 44984 63468 45055
rect 71772 45049 71856 45054
rect 70020 44985 70030 45049
rect 70094 45045 71856 45049
rect 70094 44989 71786 45045
rect 71842 44989 71856 45045
rect 70094 44985 71856 44989
rect 63394 44975 63478 44984
rect 71772 44980 71856 44985
rect 63394 44919 63408 44975
rect 63464 44919 63478 44975
rect 63394 44910 63478 44919
rect 56113 44737 56197 44742
rect 32924 44733 56197 44737
rect 32924 44677 56127 44733
rect 56183 44677 56197 44733
rect 32924 44673 56197 44677
rect 31632 41908 31717 41949
rect 31632 41844 31642 41908
rect 31706 41844 31717 41908
rect 31632 41828 31717 41844
rect 31632 41764 31642 41828
rect 31706 41764 31717 41828
rect 31632 41748 31717 41764
rect 31632 41684 31642 41748
rect 31706 41684 31717 41748
rect 31632 41644 31717 41684
rect 31634 41420 31726 41431
rect 31634 41356 31648 41420
rect 31712 41356 31726 41420
rect 31634 41340 31726 41356
rect 31634 41276 31648 41340
rect 31712 41276 31726 41340
rect 31634 41260 31726 41276
rect 31634 41196 31648 41260
rect 31712 41196 31726 41260
rect 31634 41186 31726 41196
rect 32924 40276 32988 44673
rect 40485 44609 40495 44673
rect 40559 44609 40569 44673
rect 56113 44668 56197 44673
rect 49652 44292 68174 44356
rect 68238 44292 68248 44356
rect 46649 41179 46773 41216
rect 46649 41115 46678 41179
rect 46742 41115 46773 41179
rect 46649 41083 46773 41115
rect 46669 40310 46753 40315
rect 46309 40306 46753 40310
rect 32914 40267 32998 40276
rect 32914 40211 32928 40267
rect 32984 40211 32998 40267
rect 38375 40225 39395 40289
rect 40975 40225 41995 40289
rect 43575 40225 44595 40289
rect 46309 40250 46683 40306
rect 46739 40250 46753 40306
rect 46309 40246 46753 40250
rect 46669 40241 46753 40246
rect 32914 40202 32998 40211
rect 29164 39459 29248 39468
rect 29164 39403 29178 39459
rect 29234 39403 29248 39459
rect 29164 39394 29248 39403
rect 38023 38902 38087 39922
rect 42900 39392 43048 39429
rect 42900 39328 42942 39392
rect 43006 39328 43048 39392
rect 42900 39291 43048 39328
rect 44897 38895 44961 39915
rect 41129 38494 41862 38558
rect 31567 38435 31660 38473
rect 31567 38371 31581 38435
rect 31645 38371 31660 38435
rect 31567 38355 31660 38371
rect 31567 38291 31581 38355
rect 31645 38291 31660 38355
rect 31567 38275 31660 38291
rect 31567 38211 31581 38275
rect 31645 38211 31660 38275
rect 31567 38174 31660 38211
rect 44020 38163 44104 38168
rect 43763 38159 44104 38163
rect 38854 38095 38955 38119
rect 43763 38103 44034 38159
rect 44090 38103 44104 38159
rect 43763 38099 44104 38103
rect 38854 38031 38871 38095
rect 38935 38031 38955 38095
rect 44020 38094 44104 38099
rect 38854 38008 38955 38031
rect 31566 37941 31658 37952
rect 31566 37877 31580 37941
rect 31644 37877 31658 37941
rect 31566 37861 31658 37877
rect 31566 37797 31580 37861
rect 31644 37797 31658 37861
rect 31566 37781 31658 37797
rect 31566 37717 31580 37781
rect 31644 37717 31658 37781
rect 31566 37707 31658 37717
rect 38023 36302 38087 37322
rect 44897 36295 44961 37315
rect 38372 35959 39392 36023
rect 40972 35959 41992 36023
rect 43572 35959 44592 36023
rect 46095 34245 46213 34272
rect 46095 34181 46124 34245
rect 46188 34181 46213 34245
rect 46095 34160 46213 34181
rect 49652 33841 49716 44292
rect 50335 43761 68570 43825
rect 68634 43761 68644 43825
rect 50335 34668 50399 43761
rect 57135 43535 57219 43540
rect 54269 43471 54279 43535
rect 54343 43531 57219 43535
rect 54343 43475 57149 43531
rect 57205 43475 57219 43531
rect 54343 43471 57219 43475
rect 51805 43001 51815 43065
rect 51879 43001 51889 43065
rect 53166 43001 53176 43065
rect 53240 43001 53250 43065
rect 51815 42893 51879 43001
rect 51815 42829 52369 42893
rect 53176 42892 53240 43001
rect 51279 39730 51404 39766
rect 51279 39666 51308 39730
rect 51372 39666 51404 39730
rect 51279 39635 51404 39666
rect 52305 38659 52369 42829
rect 52646 42828 53240 42892
rect 52305 38595 52542 38659
rect 52182 38435 52272 38473
rect 52182 38371 52195 38435
rect 52259 38371 52272 38435
rect 52182 38355 52272 38371
rect 52182 38291 52195 38355
rect 52259 38291 52272 38355
rect 52182 38253 52272 38291
rect 52180 38025 52244 38033
rect 52167 37982 52271 38025
rect 52167 37926 52191 37982
rect 52247 37926 52271 37982
rect 52167 37902 52271 37926
rect 52167 37846 52191 37902
rect 52247 37846 52271 37902
rect 52167 37822 52271 37846
rect 52167 37766 52191 37822
rect 52247 37766 52271 37822
rect 52167 37723 52271 37766
rect 52180 37301 52244 37723
rect 52080 37237 52244 37301
rect 51377 34860 51703 34865
rect 52080 34860 52144 37237
rect 52478 36402 52542 38595
rect 50922 34849 51167 34860
rect 50922 34785 50932 34849
rect 50996 34785 51012 34849
rect 51076 34785 51092 34849
rect 51156 34785 51167 34849
rect 51359 34844 52144 34860
rect 51359 34796 51392 34844
rect 50922 34775 51167 34785
rect 51377 34788 51392 34796
rect 51448 34788 51472 34844
rect 51528 34788 51552 34844
rect 51608 34788 51632 34844
rect 51688 34796 52144 34844
rect 51688 34788 51703 34796
rect 51377 34768 51703 34788
rect 50335 34604 51002 34668
rect 50938 34231 51002 34604
rect 50928 34222 51012 34231
rect 50928 34166 50942 34222
rect 50998 34166 51012 34222
rect 50928 34157 51012 34166
rect 51723 34222 51807 34231
rect 51723 34166 51737 34222
rect 51793 34166 51807 34222
rect 51723 34157 51807 34166
rect 51733 33841 51797 34157
rect 49652 33777 51797 33841
rect 50917 33606 51175 33619
rect 50917 33542 50934 33606
rect 50998 33542 51014 33606
rect 51078 33542 51094 33606
rect 51158 33542 51175 33606
rect 50917 33530 51175 33542
rect 51376 33602 51705 33622
rect 51376 33546 51392 33602
rect 51448 33546 51472 33602
rect 51528 33546 51552 33602
rect 51608 33546 51632 33602
rect 51688 33594 51705 33602
rect 52080 33594 52144 34796
rect 52305 36338 52542 36402
rect 52305 34260 52369 36338
rect 52646 34260 52710 42828
rect 54279 42321 54343 43471
rect 57135 43466 57219 43471
rect 80761 43404 80870 43426
rect 71755 43349 71871 43373
rect 71755 43285 71781 43349
rect 71845 43285 71871 43349
rect 80761 43340 80783 43404
rect 80847 43340 80870 43404
rect 80761 43314 80870 43340
rect 71755 43264 71871 43285
rect 56328 43234 56412 43239
rect 54686 43170 54696 43234
rect 54760 43230 56412 43234
rect 54760 43174 56342 43230
rect 56398 43174 56412 43230
rect 54760 43170 56412 43174
rect 56328 43165 56412 43170
rect 61941 43194 62298 43200
rect 60145 43128 60229 43133
rect 61941 43128 61967 43194
rect 60145 43124 61967 43128
rect 60145 43068 60159 43124
rect 60215 43068 61967 43124
rect 60145 43064 61967 43068
rect 60145 43059 60229 43064
rect 61941 43050 61967 43064
rect 62271 43128 62298 43194
rect 64169 43128 64253 43133
rect 66065 43128 66149 43133
rect 62271 43124 66183 43128
rect 62271 43068 64183 43124
rect 64239 43068 66079 43124
rect 66135 43068 66183 43124
rect 62271 43064 66183 43068
rect 67297 43080 67421 43105
rect 62271 43050 62298 43064
rect 64169 43059 64253 43064
rect 66065 43059 66149 43064
rect 61941 43044 62298 43050
rect 67297 43016 67326 43080
rect 67390 43016 67421 43080
rect 67297 42990 67421 43016
rect 78022 43084 78173 43128
rect 78022 43020 78065 43084
rect 78129 43020 78173 43084
rect 78022 42973 78173 43020
rect 62791 42932 62875 42937
rect 64790 42932 64874 42937
rect 55580 42868 55590 42932
rect 55654 42928 64874 42932
rect 55654 42872 62805 42928
rect 62861 42872 64804 42928
rect 64860 42872 64874 42928
rect 55654 42868 64874 42872
rect 62791 42863 62875 42868
rect 64790 42863 64874 42868
rect 65333 42740 65467 42780
rect 61983 42673 62067 42678
rect 63981 42673 64065 42678
rect 55951 42609 55961 42673
rect 56025 42669 64065 42673
rect 56025 42613 61997 42669
rect 62053 42613 63995 42669
rect 64051 42613 64065 42669
rect 65333 42676 65374 42740
rect 65438 42676 65467 42740
rect 70658 42710 70742 42715
rect 65333 42639 65467 42676
rect 70014 42646 70024 42710
rect 70088 42706 70742 42710
rect 70088 42650 70672 42706
rect 70728 42650 70742 42706
rect 70088 42646 70742 42650
rect 70658 42641 70742 42646
rect 56025 42609 64065 42613
rect 61983 42604 62067 42609
rect 63981 42604 64065 42609
rect 71199 42529 71209 42593
rect 71273 42529 71283 42593
rect 82698 42529 82708 42593
rect 82772 42529 82782 42593
rect 60791 42334 60875 42339
rect 66790 42334 66874 42339
rect 53585 42257 54343 42321
rect 56404 42270 56414 42334
rect 56478 42330 66874 42334
rect 56478 42274 60805 42330
rect 60861 42274 66804 42330
rect 66860 42274 66874 42330
rect 56478 42270 66874 42274
rect 60791 42265 60875 42270
rect 66790 42265 66874 42270
rect 53585 40227 53649 42257
rect 59982 42053 60066 42058
rect 65983 42053 66067 42058
rect 56800 41989 56810 42053
rect 56874 42049 66067 42053
rect 56874 41993 59996 42049
rect 60052 41993 65997 42049
rect 66053 41993 66067 42049
rect 56874 41989 66067 41993
rect 59982 41984 60066 41989
rect 65983 41984 66067 41989
rect 53873 41878 54356 41886
rect 53873 41654 53922 41878
rect 54306 41794 54356 41878
rect 57317 41794 57401 41799
rect 54306 41790 57401 41794
rect 54306 41734 57331 41790
rect 57387 41734 57401 41790
rect 54306 41730 57401 41734
rect 54306 41654 54356 41730
rect 57317 41725 57401 41730
rect 71452 41721 71462 41785
rect 71526 41721 71536 41785
rect 82445 41722 82455 41786
rect 82519 41722 82529 41786
rect 53873 41646 54356 41654
rect 71756 41564 71876 41588
rect 56263 41547 56347 41552
rect 56247 41543 58075 41547
rect 56247 41487 56277 41543
rect 56333 41487 58075 41543
rect 56247 41483 58075 41487
rect 58139 41483 58171 41547
rect 71756 41500 71783 41564
rect 71847 41500 71876 41564
rect 56263 41478 56347 41483
rect 71756 41471 71876 41500
rect 80759 41574 80872 41597
rect 80759 41510 80783 41574
rect 80847 41510 80872 41574
rect 80759 41480 80872 41510
rect 61362 41311 61481 41335
rect 61362 41247 61389 41311
rect 61453 41247 61481 41311
rect 61362 41216 61481 41247
rect 63294 41311 63413 41336
rect 63294 41247 63321 41311
rect 63385 41247 63413 41311
rect 63294 41217 63413 41247
rect 70687 41105 70771 41110
rect 70040 41041 70050 41105
rect 70114 41101 70771 41105
rect 70114 41045 70701 41101
rect 70757 41045 70771 41101
rect 70114 41041 70771 41045
rect 70687 41036 70771 41041
rect 57112 40436 68243 40473
rect 57112 40435 57357 40436
rect 54162 40292 57357 40435
rect 68221 40292 68243 40436
rect 54162 40274 68243 40292
rect 57112 40255 68243 40274
rect 53575 40163 53585 40227
rect 53649 40163 53659 40227
rect 57112 40206 57342 40255
rect 57112 40184 57291 40206
rect 54076 39476 54160 39481
rect 53156 39412 53166 39476
rect 53230 39472 54160 39476
rect 53230 39416 54090 39472
rect 54146 39416 54160 39472
rect 53230 39412 54160 39416
rect 54076 39407 54160 39412
rect 53940 38992 54043 39025
rect 53940 38928 53959 38992
rect 54023 38928 54043 38992
rect 53940 38912 54043 38928
rect 53940 38848 53959 38912
rect 54023 38848 54043 38912
rect 53940 38832 54043 38848
rect 53940 38768 53959 38832
rect 54023 38768 54043 38832
rect 53940 38736 54043 38768
rect 54061 38666 54145 38671
rect 53575 38602 53585 38666
rect 53649 38662 54145 38666
rect 53649 38606 54075 38662
rect 54131 38606 54145 38662
rect 53649 38602 54145 38606
rect 54061 38597 54145 38602
rect 57112 38015 57133 40184
rect 54138 37854 57133 38015
rect 54486 37155 54570 37164
rect 54486 37099 54500 37155
rect 54556 37099 54570 37155
rect 54486 37090 54570 37099
rect 55276 37143 55379 37160
rect 54199 36346 54283 36355
rect 54199 36290 54213 36346
rect 54269 36290 54283 36346
rect 54199 36281 54283 36290
rect 52295 34251 52379 34260
rect 52295 34195 52309 34251
rect 52365 34195 52379 34251
rect 52295 34186 52379 34195
rect 52636 34251 52720 34260
rect 52636 34195 52650 34251
rect 52706 34195 52720 34251
rect 52636 34186 52720 34195
rect 51688 33546 52144 33594
rect 51376 33530 52144 33546
rect 51376 33526 51705 33530
rect 52080 32729 52144 33530
rect 52080 32665 53909 32729
rect 53973 32665 53983 32729
rect 38375 32425 39395 32489
rect 40975 32425 41995 32489
rect 43575 32425 44595 32489
rect 38023 31102 38087 32122
rect 40303 31629 40451 31666
rect 40303 31565 40345 31629
rect 40409 31565 40451 31629
rect 40303 31528 40451 31565
rect 44897 31095 44961 32115
rect 54209 31554 54273 36281
rect 54496 32362 54560 37090
rect 55276 37079 55295 37143
rect 55359 37079 55379 37143
rect 55276 37063 55379 37079
rect 55276 36999 55295 37063
rect 55359 36999 55379 37063
rect 55276 36983 55379 36999
rect 55276 36919 55295 36983
rect 55359 36919 55379 36983
rect 55276 36903 55379 36919
rect 55276 36839 55295 36903
rect 55359 36839 55379 36903
rect 55276 36823 55379 36839
rect 55276 36759 55295 36823
rect 55359 36759 55379 36823
rect 55276 36743 55379 36759
rect 55586 36427 55670 36436
rect 55586 36371 55600 36427
rect 55656 36371 55670 36427
rect 55586 36362 55670 36371
rect 55158 35553 55242 35562
rect 55158 35497 55172 35553
rect 55228 35497 55242 35553
rect 55158 35488 55242 35497
rect 55325 35548 55411 35556
rect 54872 34747 54956 34756
rect 54872 34691 54886 34747
rect 54942 34691 54956 34747
rect 54872 34682 54956 34691
rect 54882 33156 54946 34682
rect 55168 33964 55232 35488
rect 55325 35484 55336 35548
rect 55400 35484 55411 35548
rect 55325 35468 55411 35484
rect 55325 35404 55336 35468
rect 55400 35404 55411 35468
rect 55325 35388 55411 35404
rect 55325 35324 55336 35388
rect 55400 35324 55411 35388
rect 55325 35308 55411 35324
rect 55325 35244 55336 35308
rect 55400 35244 55411 35308
rect 55325 35228 55411 35244
rect 55325 35164 55336 35228
rect 55400 35164 55411 35228
rect 55325 35157 55411 35164
rect 55596 34810 55660 36362
rect 55586 34801 55670 34810
rect 55586 34745 55600 34801
rect 55656 34745 55670 34801
rect 55586 34736 55670 34745
rect 55158 33955 55242 33964
rect 55158 33899 55172 33955
rect 55228 33899 55242 33955
rect 55158 33890 55242 33899
rect 55325 33945 55409 33957
rect 54872 33147 54956 33156
rect 54872 33091 54886 33147
rect 54942 33091 54956 33147
rect 54872 33082 54956 33091
rect 54486 32353 54570 32362
rect 54486 32297 54500 32353
rect 54556 32297 54570 32353
rect 54486 32288 54570 32297
rect 54199 31545 54283 31554
rect 54199 31489 54213 31545
rect 54269 31489 54283 31545
rect 54199 31480 54283 31489
rect 49870 31257 50353 31270
rect 49870 31253 49919 31257
rect 50303 31253 50353 31257
rect 49870 31037 49883 31253
rect 50339 31037 50353 31253
rect 49870 31033 49919 31037
rect 50303 31033 50353 31037
rect 49870 31020 50353 31033
rect 31563 30672 31658 30696
rect 41129 30694 41862 30758
rect 52167 30713 52268 30722
rect 31563 30608 31578 30672
rect 31642 30608 31658 30672
rect 31563 30592 31658 30608
rect 31563 30528 31578 30592
rect 31642 30528 31658 30592
rect 31563 30512 31658 30528
rect 31563 30448 31578 30512
rect 31642 30448 31658 30512
rect 31563 30425 31658 30448
rect 52167 30657 52189 30713
rect 52245 30671 52268 30713
rect 52245 30657 53910 30671
rect 52167 30633 53910 30657
rect 52167 30577 52189 30633
rect 52245 30607 53910 30633
rect 53974 30607 53984 30671
rect 52245 30577 52268 30607
rect 52167 30553 52268 30577
rect 52167 30497 52189 30553
rect 52245 30497 52268 30553
rect 52167 30473 52268 30497
rect 52167 30417 52189 30473
rect 52245 30417 52268 30473
rect 52167 30409 52268 30417
rect 38823 30325 38923 30350
rect 44009 30335 44093 30340
rect 38823 30261 38843 30325
rect 38907 30261 38923 30325
rect 43768 30331 44093 30335
rect 43768 30275 44023 30331
rect 44079 30275 44093 30331
rect 43768 30271 44093 30275
rect 44009 30266 44093 30271
rect 38823 30239 38923 30261
rect 31562 30185 31657 30201
rect 31562 30121 31577 30185
rect 31641 30121 31657 30185
rect 31562 30105 31657 30121
rect 31562 30041 31577 30105
rect 31641 30041 31657 30105
rect 31562 30025 31657 30041
rect 31562 29961 31577 30025
rect 31641 29961 31657 30025
rect 52177 30150 52263 30190
rect 52177 30086 52188 30150
rect 52252 30086 52263 30150
rect 52177 30070 52263 30086
rect 52177 30006 52188 30070
rect 52252 30006 52263 30070
rect 54034 30064 54118 30069
rect 52177 29967 52263 30006
rect 53156 30000 53166 30064
rect 53230 30060 54118 30064
rect 53230 30004 54048 30060
rect 54104 30004 54118 30060
rect 53230 30000 54118 30004
rect 54034 29995 54118 30000
rect 31562 29946 31657 29961
rect 53891 29570 53994 29604
rect 38023 28502 38087 29522
rect 44897 28495 44961 29515
rect 53891 29506 53910 29570
rect 53974 29506 53994 29570
rect 53891 29490 53994 29506
rect 53891 29426 53910 29490
rect 53974 29426 53994 29490
rect 53891 29410 53994 29426
rect 53891 29346 53910 29410
rect 53974 29346 53994 29410
rect 46328 29074 46392 29336
rect 53891 29313 53994 29346
rect 53575 29191 53585 29255
rect 53649 29191 53659 29255
rect 54056 29251 54140 29260
rect 54056 29195 54070 29251
rect 54126 29195 54140 29251
rect 46318 29065 46402 29074
rect 46318 29009 46332 29065
rect 46388 29009 46402 29065
rect 46318 29000 46402 29009
rect 53585 29000 53649 29191
rect 54056 29186 54140 29195
rect 54063 29000 54127 29186
rect 53585 28936 54127 29000
rect 38372 28159 39392 28223
rect 40972 28159 41992 28223
rect 43572 28159 44592 28223
rect 54209 19043 54273 31480
rect 54496 19506 54560 32288
rect 54882 20041 54946 33082
rect 55168 20513 55232 33890
rect 55325 33881 55335 33945
rect 55399 33881 55409 33945
rect 55325 33865 55409 33881
rect 55325 33801 55335 33865
rect 55399 33801 55409 33865
rect 55325 33785 55409 33801
rect 55325 33721 55335 33785
rect 55399 33721 55409 33785
rect 55325 33705 55409 33721
rect 55325 33641 55335 33705
rect 55399 33641 55409 33705
rect 55325 33625 55409 33641
rect 55325 33561 55335 33625
rect 55399 33561 55409 33625
rect 55325 33549 55409 33561
rect 55596 33152 55660 34736
rect 57112 34688 57133 37854
rect 57269 34688 57291 40184
rect 68323 40195 68503 40211
rect 68323 38459 68345 40195
rect 68481 39291 68503 40195
rect 80738 39810 80880 39842
rect 71749 39733 71875 39760
rect 71749 39669 71780 39733
rect 71844 39669 71875 39733
rect 80738 39746 80780 39810
rect 80844 39746 80880 39810
rect 80738 39707 80880 39746
rect 71749 39643 71875 39669
rect 77991 39518 78112 39548
rect 77991 39454 78022 39518
rect 78086 39454 78112 39518
rect 77991 39422 78112 39454
rect 68481 39250 70178 39291
rect 71774 39250 71858 39255
rect 68481 39186 70067 39250
rect 70131 39246 71858 39250
rect 70131 39190 71788 39246
rect 71844 39190 71858 39246
rect 70131 39186 71858 39190
rect 68481 39135 70178 39186
rect 71774 39181 71858 39186
rect 68481 38459 68503 39135
rect 68323 38443 68503 38459
rect 80758 38019 80863 38040
rect 71744 37987 71872 38019
rect 68341 37962 68488 37981
rect 68341 37906 68386 37962
rect 68442 37906 68488 37962
rect 68341 37882 68488 37906
rect 71744 37923 71779 37987
rect 71843 37923 71872 37987
rect 80758 37955 80780 38019
rect 80844 37955 80863 38019
rect 80758 37931 80863 37955
rect 71744 37882 71872 37923
rect 68341 37826 68386 37882
rect 68442 37826 68488 37882
rect 68341 37802 68488 37826
rect 68341 37746 68386 37802
rect 68442 37746 68488 37802
rect 68341 37722 68488 37746
rect 68341 37666 68386 37722
rect 68442 37666 68488 37722
rect 68341 37642 68488 37666
rect 68341 37594 68386 37642
rect 68340 37586 68386 37594
rect 68442 37594 68488 37642
rect 68442 37586 70169 37594
rect 68340 37562 70169 37586
rect 68340 37506 68386 37562
rect 68442 37550 70169 37562
rect 70720 37550 70804 37555
rect 68442 37506 70097 37550
rect 68340 37486 70097 37506
rect 70161 37546 70804 37550
rect 70161 37490 70734 37546
rect 70790 37490 70804 37546
rect 70161 37486 70804 37490
rect 68340 37482 70169 37486
rect 68340 37448 68386 37482
rect 68341 37426 68386 37448
rect 68442 37448 70169 37482
rect 70720 37481 70804 37486
rect 68442 37426 68488 37448
rect 68341 37402 68488 37426
rect 68341 37346 68386 37402
rect 68442 37346 68488 37402
rect 68341 37322 68488 37346
rect 68341 37266 68386 37322
rect 68442 37266 68488 37322
rect 68341 37242 68488 37266
rect 68341 37186 68386 37242
rect 68442 37186 68488 37242
rect 68341 37162 68488 37186
rect 68341 37106 68386 37162
rect 68442 37106 68488 37162
rect 71199 37129 71209 37193
rect 71273 37129 71283 37193
rect 68341 37082 68488 37106
rect 68341 37026 68386 37082
rect 68442 37026 68488 37082
rect 68341 37007 68488 37026
rect 71452 36321 71462 36385
rect 71526 36321 71536 36385
rect 71769 36202 71883 36224
rect 68327 36132 68502 36156
rect 68327 35356 68346 36132
rect 68482 35746 68502 36132
rect 71769 36138 71796 36202
rect 71860 36138 71883 36202
rect 71769 36109 71883 36138
rect 80761 36212 80873 36236
rect 80761 36148 80785 36212
rect 80849 36148 80873 36212
rect 80761 36120 80873 36148
rect 78039 35928 78174 35969
rect 78039 35864 78079 35928
rect 78143 35864 78174 35928
rect 78039 35826 78174 35864
rect 68482 35698 70218 35746
rect 70783 35698 70867 35703
rect 68482 35634 70095 35698
rect 70159 35694 70867 35698
rect 70159 35638 70797 35694
rect 70853 35638 70867 35694
rect 70159 35634 70867 35638
rect 68482 35582 70218 35634
rect 70783 35629 70867 35634
rect 68482 35356 68502 35582
rect 68327 35333 68502 35356
rect 57112 34657 57291 34688
rect 63567 34540 68322 34564
rect 63567 34396 63592 34540
rect 68296 34396 68322 34540
rect 63567 34373 68322 34396
rect 71760 34405 71874 34428
rect 71760 34341 71785 34405
rect 71849 34341 71874 34405
rect 71760 34312 71874 34341
rect 80758 34402 80877 34432
rect 80758 34338 80785 34402
rect 80849 34338 80877 34402
rect 80758 34308 80877 34338
rect 93137 33176 93245 33198
rect 55586 33143 55670 33152
rect 55586 33087 55600 33143
rect 55656 33087 55670 33143
rect 55586 33078 55670 33087
rect 93137 33112 93160 33176
rect 93224 33112 93245 33176
rect 93137 33086 93245 33112
rect 55326 32344 55414 32357
rect 55326 32280 55338 32344
rect 55402 32280 55414 32344
rect 55326 32264 55414 32280
rect 55326 32200 55338 32264
rect 55402 32200 55414 32264
rect 55326 32184 55414 32200
rect 55326 32120 55338 32184
rect 55402 32120 55414 32184
rect 55326 32104 55414 32120
rect 55326 32040 55338 32104
rect 55402 32040 55414 32104
rect 55326 32024 55414 32040
rect 55326 31960 55338 32024
rect 55402 31960 55414 32024
rect 55326 31947 55414 31960
rect 55596 31613 55660 33078
rect 93982 32808 94244 32814
rect 93982 32727 94001 32808
rect 91738 32663 94001 32727
rect 91738 32358 91802 32663
rect 92553 32553 92677 32585
rect 93982 32584 94001 32663
rect 94225 32584 94244 32808
rect 93982 32578 94244 32584
rect 92553 32489 92583 32553
rect 92647 32489 92677 32553
rect 92553 32458 92677 32489
rect 93698 32491 93814 32520
rect 93698 32427 93725 32491
rect 93789 32427 93814 32491
rect 93698 32399 93814 32427
rect 91738 32310 92182 32358
rect 91738 32301 92192 32310
rect 91738 32294 92122 32301
rect 55586 31604 55670 31613
rect 55586 31548 55600 31604
rect 55656 31548 55670 31604
rect 55586 31539 55670 31548
rect 55596 31285 55660 31539
rect 55586 31246 55670 31285
rect 55586 31190 55600 31246
rect 55656 31190 55670 31246
rect 55586 31166 55670 31190
rect 55586 31110 55600 31166
rect 55656 31110 55670 31166
rect 55586 31086 55670 31110
rect 55586 31030 55600 31086
rect 55656 31030 55670 31086
rect 55586 30991 55670 31030
rect 91738 31035 91802 32294
rect 92108 32245 92122 32294
rect 92178 32245 92192 32301
rect 92108 32236 92192 32245
rect 97105 32117 97363 32157
rect 95652 32055 96236 32105
rect 95652 31999 95676 32055
rect 95732 31999 96236 32055
rect 95652 31975 96236 31999
rect 95652 31919 95676 31975
rect 95732 31935 96236 31975
rect 97105 32061 97206 32117
rect 97262 32061 97363 32117
rect 97105 32037 97363 32061
rect 97105 31981 97206 32037
rect 97262 31981 97363 32037
rect 97105 31935 97363 31981
rect 95732 31919 97815 31935
rect 93101 31897 93675 31918
rect 93101 31841 93402 31897
rect 93458 31841 93482 31897
rect 93538 31841 93562 31897
rect 93618 31841 93675 31897
rect 95652 31865 97815 31919
rect 93101 31822 93675 31841
rect 92102 31245 92221 31275
rect 92102 31181 92122 31245
rect 92186 31210 92221 31245
rect 93101 31210 93197 31822
rect 95996 31695 97815 31865
rect 95652 31563 95753 31590
rect 95652 31499 95670 31563
rect 95734 31499 95753 31563
rect 95652 31483 95753 31499
rect 95652 31419 95670 31483
rect 95734 31419 95753 31483
rect 95652 31392 95753 31419
rect 93432 31356 94171 31371
rect 93432 31300 93472 31356
rect 93528 31300 93552 31356
rect 93608 31355 94171 31356
rect 93608 31300 94081 31355
rect 93432 31291 94081 31300
rect 94145 31291 94171 31355
rect 93432 31275 94171 31291
rect 92186 31181 93197 31210
rect 92102 31146 93197 31181
rect 92102 31145 92221 31146
rect 55596 30478 55660 30991
rect 91738 30981 92185 31035
rect 91738 30972 92195 30981
rect 91738 30971 92125 30972
rect 55586 30469 55670 30478
rect 55586 30413 55600 30469
rect 55656 30413 55670 30469
rect 55586 30404 55670 30413
rect 91738 29645 91802 30971
rect 92111 30916 92125 30971
rect 92181 30916 92195 30972
rect 92111 30907 92195 30916
rect 93101 30838 93197 31146
rect 93101 30822 93536 30838
rect 93101 30808 93541 30822
rect 93101 30752 93460 30808
rect 93516 30752 93541 30808
rect 95996 30787 96236 31695
rect 97171 31576 97272 31603
rect 97171 31512 97189 31576
rect 97253 31512 97272 31576
rect 97171 31496 97272 31512
rect 97171 31432 97189 31496
rect 97253 31432 97272 31496
rect 97171 31405 97272 31432
rect 97575 31192 97815 31695
rect 99686 31241 103027 31259
rect 97575 31184 98368 31192
rect 97575 30960 97934 31184
rect 98318 30960 98368 31184
rect 99686 31177 99724 31241
rect 99788 31177 99804 31241
rect 99868 31177 99884 31241
rect 99948 31177 99964 31241
rect 100028 31177 100044 31241
rect 100108 31177 100124 31241
rect 100188 31177 100204 31241
rect 100268 31177 100284 31241
rect 100348 31177 100364 31241
rect 100428 31177 100444 31241
rect 100508 31177 100524 31241
rect 100588 31177 100604 31241
rect 100668 31177 100684 31241
rect 100748 31177 100764 31241
rect 100828 31177 100844 31241
rect 100908 31177 100924 31241
rect 100988 31177 101004 31241
rect 101068 31177 101084 31241
rect 101148 31177 101164 31241
rect 101228 31177 101244 31241
rect 101308 31177 101324 31241
rect 101388 31177 101404 31241
rect 101468 31177 101484 31241
rect 101548 31177 101564 31241
rect 101628 31177 101644 31241
rect 101708 31177 101724 31241
rect 101788 31177 101804 31241
rect 101868 31177 101884 31241
rect 101948 31177 101964 31241
rect 102028 31177 102044 31241
rect 102108 31177 102124 31241
rect 102188 31177 102204 31241
rect 102268 31177 102284 31241
rect 102348 31177 102364 31241
rect 102428 31177 102444 31241
rect 102508 31177 102524 31241
rect 102588 31177 102604 31241
rect 102668 31177 102684 31241
rect 102748 31177 102764 31241
rect 102828 31177 102844 31241
rect 102908 31177 102924 31241
rect 102988 31177 103027 31241
rect 99686 31160 103027 31177
rect 97575 30952 98368 30960
rect 97575 30819 97815 30952
rect 93101 30742 93541 30752
rect 93436 30738 93541 30742
rect 92094 29907 92202 29930
rect 92094 29843 92121 29907
rect 92185 29888 92202 29907
rect 92185 29843 92738 29888
rect 92094 29824 92738 29843
rect 92094 29818 92202 29824
rect 92674 29736 92738 29824
rect 93440 29749 93536 30738
rect 95635 30694 96236 30787
rect 95635 30638 95676 30694
rect 95732 30638 96236 30694
rect 95635 30547 96236 30638
rect 97170 30781 97815 30819
rect 97170 30725 97198 30781
rect 97254 30725 97815 30781
rect 97170 30701 97815 30725
rect 97170 30645 97198 30701
rect 97254 30645 97815 30701
rect 97170 30579 97815 30645
rect 94055 30271 94171 30292
rect 94055 30207 94081 30271
rect 94145 30207 94171 30271
rect 94055 30186 94171 30207
rect 95647 30232 95748 30259
rect 95647 30168 95665 30232
rect 95729 30168 95748 30232
rect 95647 30152 95748 30168
rect 95647 30088 95665 30152
rect 95729 30088 95748 30152
rect 95647 30061 95748 30088
rect 93028 29736 93536 29749
rect 92674 29725 93536 29736
rect 92674 29672 93085 29725
rect 93028 29669 93085 29672
rect 93141 29669 93165 29725
rect 93221 29669 93536 29725
rect 93028 29653 93536 29669
rect 91738 29589 92182 29645
rect 91738 29581 92192 29589
rect 91738 28310 91802 29581
rect 92108 29580 92192 29581
rect 92108 29524 92122 29580
rect 92178 29524 92192 29580
rect 92108 29515 92192 29524
rect 93028 28749 93124 29653
rect 95996 29417 96236 30547
rect 97176 30229 97277 30256
rect 97176 30165 97194 30229
rect 97258 30165 97277 30229
rect 97176 30149 97277 30165
rect 97176 30085 97194 30149
rect 97258 30085 97277 30149
rect 97176 30058 97277 30085
rect 97575 29438 97815 30579
rect 104557 29822 104813 29827
rect 104557 29812 120001 29822
rect 104557 29596 104577 29812
rect 104793 29596 120001 29812
rect 104557 29586 120001 29596
rect 104557 29581 104813 29586
rect 95655 29304 96236 29417
rect 95655 29248 95677 29304
rect 95733 29248 96236 29304
rect 93592 29183 94171 29199
rect 93592 29177 94081 29183
rect 93592 29121 93610 29177
rect 93666 29121 93690 29177
rect 93746 29121 93770 29177
rect 93826 29121 94081 29177
rect 93592 29119 94081 29121
rect 94145 29119 94171 29183
rect 95655 29177 96236 29248
rect 97182 29401 97815 29438
rect 97182 29345 97215 29401
rect 97271 29345 97815 29401
rect 97182 29321 97815 29345
rect 97182 29265 97215 29321
rect 97271 29265 97815 29321
rect 97182 29198 97815 29265
rect 93592 29103 94171 29119
rect 95646 28879 95747 28906
rect 95646 28815 95664 28879
rect 95728 28815 95747 28879
rect 95646 28799 95747 28815
rect 93028 28655 93539 28749
rect 95646 28735 95664 28799
rect 95728 28735 95747 28799
rect 95646 28708 95747 28735
rect 93028 28653 93631 28655
rect 93443 28634 93631 28653
rect 93443 28578 93462 28634
rect 93518 28578 93542 28634
rect 93598 28578 93631 28634
rect 93443 28559 93631 28578
rect 92108 28514 92213 28538
rect 92108 28450 92129 28514
rect 92193 28502 92213 28514
rect 93443 28502 93539 28559
rect 92193 28450 93539 28502
rect 92108 28438 93539 28450
rect 92108 28425 92213 28438
rect 91738 28246 92182 28310
rect 92108 28214 92182 28246
rect 92108 28205 92192 28214
rect 92108 28149 92122 28205
rect 92178 28149 92192 28205
rect 92108 28140 92192 28149
rect 93443 27649 93539 28438
rect 94056 28095 94172 28116
rect 94056 28031 94082 28095
rect 94146 28031 94172 28095
rect 94056 28010 94172 28031
rect 95996 28008 96236 29177
rect 97176 28857 97277 28884
rect 97176 28793 97194 28857
rect 97258 28793 97277 28857
rect 97176 28777 97277 28793
rect 97176 28713 97194 28777
rect 97258 28713 97277 28777
rect 97176 28686 97277 28713
rect 97575 28289 97815 29198
rect 97575 28281 98366 28289
rect 95642 27947 96236 28008
rect 95642 27891 95677 27947
rect 95733 27891 96236 27947
rect 95642 27867 96236 27891
rect 95642 27811 95677 27867
rect 95733 27840 96236 27867
rect 97109 28022 97349 28059
rect 97109 27966 97205 28022
rect 97261 27966 97349 28022
rect 97109 27942 97349 27966
rect 97109 27886 97205 27942
rect 97261 27886 97349 27942
rect 97109 27840 97349 27886
rect 97575 28057 97932 28281
rect 98316 28057 98366 28281
rect 99683 28242 103063 28260
rect 99683 28178 99701 28242
rect 99765 28178 99781 28242
rect 99845 28178 99861 28242
rect 99925 28178 99941 28242
rect 100005 28178 100021 28242
rect 100085 28178 100101 28242
rect 100165 28178 100181 28242
rect 100245 28178 100261 28242
rect 100325 28178 100341 28242
rect 100405 28178 100421 28242
rect 100485 28178 100501 28242
rect 100565 28178 100581 28242
rect 100645 28178 100661 28242
rect 100725 28178 100741 28242
rect 100805 28178 100821 28242
rect 100885 28178 100901 28242
rect 100965 28178 100981 28242
rect 101045 28178 101061 28242
rect 101125 28178 101141 28242
rect 101205 28178 101221 28242
rect 101285 28178 101301 28242
rect 101365 28178 101381 28242
rect 101445 28178 101461 28242
rect 101525 28178 101541 28242
rect 101605 28178 101621 28242
rect 101685 28178 101701 28242
rect 101765 28178 101781 28242
rect 101845 28178 101861 28242
rect 101925 28178 101941 28242
rect 102005 28178 102021 28242
rect 102085 28178 102101 28242
rect 102165 28178 102181 28242
rect 102245 28178 102261 28242
rect 102325 28178 102341 28242
rect 102405 28178 102421 28242
rect 102485 28178 102501 28242
rect 102565 28178 102581 28242
rect 102645 28178 102661 28242
rect 102725 28178 102741 28242
rect 102805 28178 102821 28242
rect 102885 28178 102901 28242
rect 102965 28178 102981 28242
rect 103045 28178 103063 28242
rect 99683 28161 103063 28178
rect 97575 28049 98366 28057
rect 97575 27840 97815 28049
rect 95733 27811 97815 27840
rect 95642 27768 97815 27811
rect 93443 27558 93542 27649
rect 95996 27600 97815 27768
rect 93443 27545 93590 27558
rect 93443 27489 93488 27545
rect 93544 27489 93590 27545
rect 93443 27476 93590 27489
rect 95649 27479 95750 27506
rect 92099 27144 92210 27166
rect 92099 27080 92125 27144
rect 92189 27135 92210 27144
rect 93453 27135 93517 27476
rect 95649 27415 95667 27479
rect 95731 27415 95750 27479
rect 95649 27399 95750 27415
rect 95649 27335 95667 27399
rect 95731 27335 95750 27399
rect 95649 27308 95750 27335
rect 97173 27473 97274 27500
rect 97173 27409 97191 27473
rect 97255 27409 97274 27473
rect 97173 27393 97274 27409
rect 97173 27329 97191 27393
rect 97255 27329 97274 27393
rect 97173 27302 97274 27329
rect 92189 27080 93517 27135
rect 92099 27071 93517 27080
rect 92099 27051 92210 27071
rect 97575 27067 97815 27600
rect 93137 26236 93245 26258
rect 93137 26172 93160 26236
rect 93224 26172 93245 26236
rect 93137 26146 93245 26172
rect 93982 25868 94244 25874
rect 93982 25787 94001 25868
rect 91738 25723 94001 25787
rect 91738 25418 91802 25723
rect 92553 25613 92677 25645
rect 93982 25644 94001 25723
rect 94225 25644 94244 25868
rect 93982 25638 94244 25644
rect 92553 25549 92583 25613
rect 92647 25549 92677 25613
rect 92553 25518 92677 25549
rect 93698 25551 93814 25580
rect 93698 25487 93725 25551
rect 93789 25487 93814 25551
rect 93698 25459 93814 25487
rect 91738 25370 92182 25418
rect 91738 25361 92192 25370
rect 91738 25354 92122 25361
rect 57406 24243 78211 24259
rect 57406 24099 57416 24243
rect 78200 24099 78211 24243
rect 57406 24084 78211 24099
rect 91738 24095 91802 25354
rect 92108 25305 92122 25354
rect 92178 25305 92192 25361
rect 92108 25296 92192 25305
rect 97105 25177 97363 25217
rect 95652 25115 96236 25165
rect 95652 25059 95676 25115
rect 95732 25059 96236 25115
rect 95652 25035 96236 25059
rect 95652 24979 95676 25035
rect 95732 24995 96236 25035
rect 97105 25121 97206 25177
rect 97262 25121 97363 25177
rect 97105 25097 97363 25121
rect 97105 25041 97206 25097
rect 97262 25041 97363 25097
rect 97105 24995 97363 25041
rect 95732 24979 97815 24995
rect 93101 24957 93675 24978
rect 93101 24901 93402 24957
rect 93458 24901 93482 24957
rect 93538 24901 93562 24957
rect 93618 24901 93675 24957
rect 95652 24925 97815 24979
rect 93101 24882 93675 24901
rect 92102 24305 92221 24335
rect 92102 24241 92122 24305
rect 92186 24270 92221 24305
rect 93101 24270 93197 24882
rect 95996 24755 97815 24925
rect 95652 24623 95753 24650
rect 95652 24559 95670 24623
rect 95734 24559 95753 24623
rect 95652 24543 95753 24559
rect 95652 24479 95670 24543
rect 95734 24479 95753 24543
rect 95652 24452 95753 24479
rect 93432 24416 94171 24431
rect 93432 24360 93472 24416
rect 93528 24360 93552 24416
rect 93608 24415 94171 24416
rect 93608 24360 94081 24415
rect 93432 24351 94081 24360
rect 94145 24351 94171 24415
rect 93432 24335 94171 24351
rect 92186 24241 93197 24270
rect 92102 24206 93197 24241
rect 92102 24205 92221 24206
rect 91738 24041 92185 24095
rect 91738 24032 92195 24041
rect 91738 24031 92125 24032
rect 91738 22705 91802 24031
rect 92111 23976 92125 24031
rect 92181 23976 92195 24032
rect 92111 23967 92195 23976
rect 93101 23898 93197 24206
rect 93101 23882 93536 23898
rect 93101 23868 93541 23882
rect 93101 23812 93460 23868
rect 93516 23812 93541 23868
rect 95996 23847 96236 24755
rect 97171 24636 97272 24663
rect 97171 24572 97189 24636
rect 97253 24572 97272 24636
rect 97171 24556 97272 24572
rect 97171 24492 97189 24556
rect 97253 24492 97272 24556
rect 97171 24465 97272 24492
rect 97575 24252 97815 24755
rect 99683 24308 103034 24336
rect 97575 24244 98368 24252
rect 97575 24020 97934 24244
rect 98318 24020 98368 24244
rect 99683 24244 99726 24308
rect 99790 24244 99806 24308
rect 99870 24244 99886 24308
rect 99950 24244 99966 24308
rect 100030 24244 100046 24308
rect 100110 24244 100126 24308
rect 100190 24244 100206 24308
rect 100270 24244 100286 24308
rect 100350 24244 100366 24308
rect 100430 24244 100446 24308
rect 100510 24244 100526 24308
rect 100590 24244 100606 24308
rect 100670 24244 100686 24308
rect 100750 24244 100766 24308
rect 100830 24244 100846 24308
rect 100910 24244 100926 24308
rect 100990 24244 101006 24308
rect 101070 24244 101086 24308
rect 101150 24244 101166 24308
rect 101230 24244 101246 24308
rect 101310 24244 101326 24308
rect 101390 24244 101406 24308
rect 101470 24244 101486 24308
rect 101550 24244 101566 24308
rect 101630 24244 101646 24308
rect 101710 24244 101726 24308
rect 101790 24244 101806 24308
rect 101870 24244 101886 24308
rect 101950 24244 101966 24308
rect 102030 24244 102046 24308
rect 102110 24244 102126 24308
rect 102190 24244 102206 24308
rect 102270 24244 102286 24308
rect 102350 24244 102366 24308
rect 102430 24244 102446 24308
rect 102510 24244 102526 24308
rect 102590 24244 102606 24308
rect 102670 24244 102686 24308
rect 102750 24244 102766 24308
rect 102830 24244 102846 24308
rect 102910 24244 102926 24308
rect 102990 24244 103034 24308
rect 99683 24216 103034 24244
rect 97575 24012 98368 24020
rect 97575 23879 97815 24012
rect 93101 23802 93541 23812
rect 93436 23798 93541 23802
rect 92094 22967 92202 22990
rect 92094 22903 92121 22967
rect 92185 22948 92202 22967
rect 92185 22903 92738 22948
rect 92094 22884 92738 22903
rect 92094 22878 92202 22884
rect 92674 22796 92738 22884
rect 93440 22809 93536 23798
rect 95635 23754 96236 23847
rect 95635 23698 95676 23754
rect 95732 23698 96236 23754
rect 95635 23607 96236 23698
rect 97170 23841 97815 23879
rect 97170 23785 97198 23841
rect 97254 23785 97815 23841
rect 97170 23761 97815 23785
rect 97170 23705 97198 23761
rect 97254 23705 97815 23761
rect 97170 23639 97815 23705
rect 94055 23331 94171 23352
rect 94055 23267 94081 23331
rect 94145 23267 94171 23331
rect 94055 23246 94171 23267
rect 95647 23292 95748 23319
rect 95647 23228 95665 23292
rect 95729 23228 95748 23292
rect 95647 23212 95748 23228
rect 95647 23148 95665 23212
rect 95729 23148 95748 23212
rect 95647 23121 95748 23148
rect 93028 22796 93536 22809
rect 92674 22785 93536 22796
rect 92674 22732 93085 22785
rect 93028 22729 93085 22732
rect 93141 22729 93165 22785
rect 93221 22729 93536 22785
rect 93028 22713 93536 22729
rect 91738 22649 92182 22705
rect 91738 22641 92192 22649
rect 91738 21370 91802 22641
rect 92108 22640 92192 22641
rect 92108 22584 92122 22640
rect 92178 22584 92192 22640
rect 92108 22575 92192 22584
rect 93028 21809 93124 22713
rect 95996 22477 96236 23607
rect 97176 23289 97277 23316
rect 97176 23225 97194 23289
rect 97258 23225 97277 23289
rect 97176 23209 97277 23225
rect 97176 23145 97194 23209
rect 97258 23145 97277 23209
rect 97176 23118 97277 23145
rect 97575 22498 97815 23639
rect 104573 22882 104829 22887
rect 104573 22872 120001 22882
rect 104573 22656 104593 22872
rect 104809 22656 120001 22872
rect 104573 22646 120001 22656
rect 104573 22641 104829 22646
rect 95655 22364 96236 22477
rect 95655 22308 95677 22364
rect 95733 22308 96236 22364
rect 93592 22243 94171 22259
rect 93592 22237 94081 22243
rect 93592 22181 93610 22237
rect 93666 22181 93690 22237
rect 93746 22181 93770 22237
rect 93826 22181 94081 22237
rect 93592 22179 94081 22181
rect 94145 22179 94171 22243
rect 95655 22237 96236 22308
rect 97182 22461 97815 22498
rect 97182 22405 97215 22461
rect 97271 22405 97815 22461
rect 97182 22381 97815 22405
rect 97182 22325 97215 22381
rect 97271 22325 97815 22381
rect 97182 22258 97815 22325
rect 93592 22163 94171 22179
rect 95646 21939 95747 21966
rect 95646 21875 95664 21939
rect 95728 21875 95747 21939
rect 95646 21859 95747 21875
rect 93028 21715 93539 21809
rect 95646 21795 95664 21859
rect 95728 21795 95747 21859
rect 95646 21768 95747 21795
rect 93028 21713 93631 21715
rect 93443 21694 93631 21713
rect 93443 21638 93462 21694
rect 93518 21638 93542 21694
rect 93598 21638 93631 21694
rect 93443 21619 93631 21638
rect 92108 21574 92213 21598
rect 92108 21510 92129 21574
rect 92193 21562 92213 21574
rect 93443 21562 93539 21619
rect 92193 21510 93539 21562
rect 92108 21498 93539 21510
rect 92108 21485 92213 21498
rect 91738 21306 92182 21370
rect 92108 21274 92182 21306
rect 92108 21265 92192 21274
rect 92108 21209 92122 21265
rect 92178 21209 92192 21265
rect 92108 21200 92192 21209
rect 93443 20709 93539 21498
rect 94056 21155 94172 21176
rect 94056 21091 94082 21155
rect 94146 21091 94172 21155
rect 94056 21070 94172 21091
rect 95996 21068 96236 22237
rect 97176 21917 97277 21944
rect 97176 21853 97194 21917
rect 97258 21853 97277 21917
rect 97176 21837 97277 21853
rect 97176 21773 97194 21837
rect 97258 21773 97277 21837
rect 97176 21746 97277 21773
rect 97575 21349 97815 22258
rect 97575 21341 98366 21349
rect 95642 21007 96236 21068
rect 95642 20951 95677 21007
rect 95733 20951 96236 21007
rect 95642 20927 96236 20951
rect 95642 20871 95677 20927
rect 95733 20900 96236 20927
rect 97109 21082 97349 21119
rect 97109 21026 97205 21082
rect 97261 21026 97349 21082
rect 97109 21002 97349 21026
rect 97109 20946 97205 21002
rect 97261 20946 97349 21002
rect 97109 20900 97349 20946
rect 97575 21117 97932 21341
rect 98316 21117 98366 21341
rect 99671 21302 103037 21319
rect 99671 21238 99682 21302
rect 99746 21238 99762 21302
rect 99826 21238 99842 21302
rect 99906 21238 99922 21302
rect 99986 21238 100002 21302
rect 100066 21238 100082 21302
rect 100146 21238 100162 21302
rect 100226 21238 100242 21302
rect 100306 21238 100322 21302
rect 100386 21238 100402 21302
rect 100466 21238 100482 21302
rect 100546 21238 100562 21302
rect 100626 21238 100642 21302
rect 100706 21238 100722 21302
rect 100786 21238 100802 21302
rect 100866 21238 100882 21302
rect 100946 21238 100962 21302
rect 101026 21238 101042 21302
rect 101106 21238 101122 21302
rect 101186 21238 101202 21302
rect 101266 21238 101282 21302
rect 101346 21238 101362 21302
rect 101426 21238 101442 21302
rect 101506 21238 101522 21302
rect 101586 21238 101602 21302
rect 101666 21238 101682 21302
rect 101746 21238 101762 21302
rect 101826 21238 101842 21302
rect 101906 21238 101922 21302
rect 101986 21238 102002 21302
rect 102066 21238 102082 21302
rect 102146 21238 102162 21302
rect 102226 21238 102242 21302
rect 102306 21238 102322 21302
rect 102386 21238 102402 21302
rect 102466 21238 102482 21302
rect 102546 21238 102562 21302
rect 102626 21238 102642 21302
rect 102706 21238 102722 21302
rect 102786 21238 102802 21302
rect 102866 21238 102882 21302
rect 102946 21238 102962 21302
rect 103026 21238 103037 21302
rect 99671 21221 103037 21238
rect 97575 21109 98366 21117
rect 97575 20900 97815 21109
rect 95733 20871 97815 20900
rect 95642 20828 97815 20871
rect 93443 20618 93542 20709
rect 95996 20660 97815 20828
rect 93443 20605 93590 20618
rect 93443 20549 93488 20605
rect 93544 20549 93590 20605
rect 93443 20536 93590 20549
rect 95649 20539 95750 20566
rect 55168 20449 78296 20513
rect 78360 20449 78370 20513
rect 92099 20204 92210 20226
rect 92099 20140 92125 20204
rect 92189 20195 92210 20204
rect 93453 20195 93517 20536
rect 95649 20475 95667 20539
rect 95731 20475 95750 20539
rect 95649 20459 95750 20475
rect 95649 20395 95667 20459
rect 95731 20395 95750 20459
rect 95649 20368 95750 20395
rect 97173 20533 97274 20560
rect 97173 20469 97191 20533
rect 97255 20469 97274 20533
rect 97173 20453 97274 20469
rect 97173 20389 97191 20453
rect 97255 20389 97274 20453
rect 97173 20362 97274 20389
rect 92189 20140 93517 20195
rect 92099 20131 93517 20140
rect 92099 20111 92210 20131
rect 97575 20127 97815 20660
rect 54882 19977 78296 20041
rect 78360 19977 78370 20041
rect 54496 19442 78296 19506
rect 78360 19442 78370 19506
rect 54209 18979 78296 19043
rect 78360 18979 78370 19043
rect 53489 17178 53601 17205
rect 53489 17114 53513 17178
rect 53577 17114 53601 17178
rect 53489 17098 53601 17114
rect 53489 17034 53513 17098
rect 53577 17034 53601 17098
rect 53489 17018 53601 17034
rect 53489 16954 53513 17018
rect 53577 16954 53601 17018
rect 53489 16938 53601 16954
rect 53489 16874 53513 16938
rect 53577 16874 53601 16938
rect 53489 16858 53601 16874
rect 53489 16794 53513 16858
rect 53577 16794 53601 16858
rect 53489 16778 53601 16794
rect 53489 16714 53513 16778
rect 53577 16714 53601 16778
rect 53489 16698 53601 16714
rect 53489 16634 53513 16698
rect 53577 16634 53601 16698
rect 53489 16618 53601 16634
rect 53489 16554 53513 16618
rect 53577 16554 53601 16618
rect 53489 16538 53601 16554
rect 53489 16474 53513 16538
rect 53577 16474 53601 16538
rect 53489 16458 53601 16474
rect 53489 16394 53513 16458
rect 53577 16394 53601 16458
rect 53489 16378 53601 16394
rect 53489 16314 53513 16378
rect 53577 16314 53601 16378
rect 53489 16298 53601 16314
rect 53489 16234 53513 16298
rect 53577 16234 53601 16298
rect 53489 16218 53601 16234
rect 53489 16154 53513 16218
rect 53577 16154 53601 16218
rect 53489 16138 53601 16154
rect 53489 16074 53513 16138
rect 53577 16074 53601 16138
rect 53489 16058 53601 16074
rect 53489 15994 53513 16058
rect 53577 15994 53601 16058
rect 53489 15978 53601 15994
rect 53489 15914 53513 15978
rect 53577 15914 53601 15978
rect 53489 15898 53601 15914
rect 53489 15834 53513 15898
rect 53577 15834 53601 15898
rect 53489 15818 53601 15834
rect 53489 15754 53513 15818
rect 53577 15754 53601 15818
rect 53489 15738 53601 15754
rect 53489 15674 53513 15738
rect 53577 15674 53601 15738
rect 53489 15658 53601 15674
rect 53489 15594 53513 15658
rect 53577 15594 53601 15658
rect 53489 15578 53601 15594
rect 53489 15514 53513 15578
rect 53577 15514 53601 15578
rect 53489 15498 53601 15514
rect 53489 15434 53513 15498
rect 53577 15434 53601 15498
rect 53489 15418 53601 15434
rect 53489 15354 53513 15418
rect 53577 15354 53601 15418
rect 53489 15338 53601 15354
rect 53489 15274 53513 15338
rect 53577 15274 53601 15338
rect 53489 15258 53601 15274
rect 53489 15194 53513 15258
rect 53577 15194 53601 15258
rect 53489 15178 53601 15194
rect 53489 15114 53513 15178
rect 53577 15114 53601 15178
rect 53489 15098 53601 15114
rect 53489 15034 53513 15098
rect 53577 15034 53601 15098
rect 53489 15018 53601 15034
rect 53489 14954 53513 15018
rect 53577 14954 53601 15018
rect 53489 14938 53601 14954
rect 53489 14874 53513 14938
rect 53577 14874 53601 14938
rect 53489 14858 53601 14874
rect 53489 14794 53513 14858
rect 53577 14794 53601 14858
rect 53489 14778 53601 14794
rect 53489 14714 53513 14778
rect 53577 14714 53601 14778
rect 53489 14698 53601 14714
rect 53489 14634 53513 14698
rect 53577 14634 53601 14698
rect 53489 14618 53601 14634
rect 53489 14554 53513 14618
rect 53577 14554 53601 14618
rect 53489 14538 53601 14554
rect 53489 14474 53513 14538
rect 53577 14474 53601 14538
rect 53489 14458 53601 14474
rect 53489 14394 53513 14458
rect 53577 14394 53601 14458
rect 53489 14378 53601 14394
rect 53489 14314 53513 14378
rect 53577 14314 53601 14378
rect 53489 14298 53601 14314
rect 53489 14234 53513 14298
rect 53577 14234 53601 14298
rect 53489 14218 53601 14234
rect 53489 14154 53513 14218
rect 53577 14154 53601 14218
rect 53489 14138 53601 14154
rect 53489 14074 53513 14138
rect 53577 14074 53601 14138
rect 53489 14058 53601 14074
rect 53489 13994 53513 14058
rect 53577 13994 53601 14058
rect 53489 13978 53601 13994
rect 53489 13914 53513 13978
rect 53577 13914 53601 13978
rect 53489 13887 53601 13914
rect 56484 17171 56618 17202
rect 56484 17107 56519 17171
rect 56583 17107 56618 17171
rect 56484 17091 56618 17107
rect 56484 17027 56519 17091
rect 56583 17027 56618 17091
rect 56484 17011 56618 17027
rect 56484 16947 56519 17011
rect 56583 16947 56618 17011
rect 56484 16931 56618 16947
rect 56484 16867 56519 16931
rect 56583 16867 56618 16931
rect 56484 16851 56618 16867
rect 56484 16787 56519 16851
rect 56583 16787 56618 16851
rect 56484 16771 56618 16787
rect 56484 16707 56519 16771
rect 56583 16707 56618 16771
rect 56484 16691 56618 16707
rect 56484 16627 56519 16691
rect 56583 16627 56618 16691
rect 56484 16611 56618 16627
rect 56484 16547 56519 16611
rect 56583 16547 56618 16611
rect 56484 16531 56618 16547
rect 56484 16467 56519 16531
rect 56583 16467 56618 16531
rect 56484 16451 56618 16467
rect 56484 16387 56519 16451
rect 56583 16387 56618 16451
rect 56484 16371 56618 16387
rect 56484 16307 56519 16371
rect 56583 16307 56618 16371
rect 56484 16291 56618 16307
rect 56484 16227 56519 16291
rect 56583 16227 56618 16291
rect 56484 16211 56618 16227
rect 56484 16147 56519 16211
rect 56583 16147 56618 16211
rect 56484 16131 56618 16147
rect 56484 16067 56519 16131
rect 56583 16067 56618 16131
rect 56484 16051 56618 16067
rect 56484 15987 56519 16051
rect 56583 15987 56618 16051
rect 56484 15971 56618 15987
rect 56484 15907 56519 15971
rect 56583 15907 56618 15971
rect 56484 15891 56618 15907
rect 56484 15827 56519 15891
rect 56583 15827 56618 15891
rect 56484 15811 56618 15827
rect 56484 15747 56519 15811
rect 56583 15747 56618 15811
rect 56484 15731 56618 15747
rect 56484 15667 56519 15731
rect 56583 15667 56618 15731
rect 56484 15651 56618 15667
rect 56484 15587 56519 15651
rect 56583 15587 56618 15651
rect 56484 15571 56618 15587
rect 56484 15507 56519 15571
rect 56583 15507 56618 15571
rect 56484 15491 56618 15507
rect 56484 15427 56519 15491
rect 56583 15427 56618 15491
rect 56484 15411 56618 15427
rect 56484 15347 56519 15411
rect 56583 15347 56618 15411
rect 56484 15331 56618 15347
rect 56484 15267 56519 15331
rect 56583 15267 56618 15331
rect 56484 15251 56618 15267
rect 56484 15187 56519 15251
rect 56583 15187 56618 15251
rect 56484 15171 56618 15187
rect 56484 15107 56519 15171
rect 56583 15107 56618 15171
rect 56484 15091 56618 15107
rect 56484 15027 56519 15091
rect 56583 15027 56618 15091
rect 56484 15011 56618 15027
rect 56484 14947 56519 15011
rect 56583 14947 56618 15011
rect 56484 14931 56618 14947
rect 56484 14867 56519 14931
rect 56583 14867 56618 14931
rect 56484 14851 56618 14867
rect 56484 14787 56519 14851
rect 56583 14787 56618 14851
rect 56484 14771 56618 14787
rect 56484 14707 56519 14771
rect 56583 14707 56618 14771
rect 56484 14691 56618 14707
rect 56484 14627 56519 14691
rect 56583 14627 56618 14691
rect 56484 14611 56618 14627
rect 56484 14547 56519 14611
rect 56583 14547 56618 14611
rect 56484 14531 56618 14547
rect 56484 14467 56519 14531
rect 56583 14467 56618 14531
rect 56484 14451 56618 14467
rect 56484 14387 56519 14451
rect 56583 14387 56618 14451
rect 56484 14371 56618 14387
rect 56484 14307 56519 14371
rect 56583 14307 56618 14371
rect 56484 14291 56618 14307
rect 56484 14227 56519 14291
rect 56583 14227 56618 14291
rect 56484 14211 56618 14227
rect 56484 14147 56519 14211
rect 56583 14147 56618 14211
rect 56484 14131 56618 14147
rect 56484 14067 56519 14131
rect 56583 14067 56618 14131
rect 56484 14051 56618 14067
rect 56484 13987 56519 14051
rect 56583 13987 56618 14051
rect 56484 13971 56618 13987
rect 56484 13907 56519 13971
rect 56583 13907 56618 13971
rect 56484 13877 56618 13907
rect 54905 11930 55161 11945
rect 54905 11714 54925 11930
rect 55141 11714 55161 11930
rect 54905 11699 55161 11714
rect 54915 5157 55151 11699
rect 54915 4921 56209 5157
rect 55973 0 56209 4921
<< via3 >>
rect 40263 100710 40327 100714
rect 40263 100654 40267 100710
rect 40267 100654 40323 100710
rect 40323 100654 40327 100710
rect 40263 100650 40327 100654
rect 40263 100630 40327 100634
rect 40263 100574 40267 100630
rect 40267 100574 40323 100630
rect 40323 100574 40327 100630
rect 40263 100570 40327 100574
rect 40263 100550 40327 100554
rect 40263 100494 40267 100550
rect 40267 100494 40323 100550
rect 40323 100494 40327 100550
rect 40263 100490 40327 100494
rect 40263 100470 40327 100474
rect 40263 100414 40267 100470
rect 40267 100414 40323 100470
rect 40323 100414 40327 100470
rect 40263 100410 40327 100414
rect 40263 100390 40327 100394
rect 40263 100334 40267 100390
rect 40267 100334 40323 100390
rect 40323 100334 40327 100390
rect 40263 100330 40327 100334
rect 40263 100310 40327 100314
rect 40263 100254 40267 100310
rect 40267 100254 40323 100310
rect 40323 100254 40327 100310
rect 40263 100250 40327 100254
rect 40263 100230 40327 100234
rect 40263 100174 40267 100230
rect 40267 100174 40323 100230
rect 40323 100174 40327 100230
rect 40263 100170 40327 100174
rect 40263 100150 40327 100154
rect 40263 100094 40267 100150
rect 40267 100094 40323 100150
rect 40323 100094 40327 100150
rect 40263 100090 40327 100094
rect 40263 100070 40327 100074
rect 40263 100014 40267 100070
rect 40267 100014 40323 100070
rect 40323 100014 40327 100070
rect 40263 100010 40327 100014
rect 40263 99990 40327 99994
rect 40263 99934 40267 99990
rect 40267 99934 40323 99990
rect 40323 99934 40327 99990
rect 40263 99930 40327 99934
rect 40263 99910 40327 99914
rect 40263 99854 40267 99910
rect 40267 99854 40323 99910
rect 40323 99854 40327 99910
rect 40263 99850 40327 99854
rect 40263 99830 40327 99834
rect 40263 99774 40267 99830
rect 40267 99774 40323 99830
rect 40323 99774 40327 99830
rect 40263 99770 40327 99774
rect 40263 99750 40327 99754
rect 40263 99694 40267 99750
rect 40267 99694 40323 99750
rect 40323 99694 40327 99750
rect 40263 99690 40327 99694
rect 40263 99670 40327 99674
rect 40263 99614 40267 99670
rect 40267 99614 40323 99670
rect 40323 99614 40327 99670
rect 40263 99610 40327 99614
rect 40263 99590 40327 99594
rect 40263 99534 40267 99590
rect 40267 99534 40323 99590
rect 40323 99534 40327 99590
rect 40263 99530 40327 99534
rect 40263 99510 40327 99514
rect 40263 99454 40267 99510
rect 40267 99454 40323 99510
rect 40323 99454 40327 99510
rect 40263 99450 40327 99454
rect 40263 99430 40327 99434
rect 40263 99374 40267 99430
rect 40267 99374 40323 99430
rect 40323 99374 40327 99430
rect 40263 99370 40327 99374
rect 40263 99350 40327 99354
rect 40263 99294 40267 99350
rect 40267 99294 40323 99350
rect 40323 99294 40327 99350
rect 40263 99290 40327 99294
rect 40263 99270 40327 99274
rect 40263 99214 40267 99270
rect 40267 99214 40323 99270
rect 40323 99214 40327 99270
rect 40263 99210 40327 99214
rect 40263 99190 40327 99194
rect 40263 99134 40267 99190
rect 40267 99134 40323 99190
rect 40323 99134 40327 99190
rect 40263 99130 40327 99134
rect 40263 99110 40327 99114
rect 40263 99054 40267 99110
rect 40267 99054 40323 99110
rect 40323 99054 40327 99110
rect 40263 99050 40327 99054
rect 40263 99030 40327 99034
rect 40263 98974 40267 99030
rect 40267 98974 40323 99030
rect 40323 98974 40327 99030
rect 40263 98970 40327 98974
rect 40263 98950 40327 98954
rect 40263 98894 40267 98950
rect 40267 98894 40323 98950
rect 40323 98894 40327 98950
rect 40263 98890 40327 98894
rect 40263 98870 40327 98874
rect 40263 98814 40267 98870
rect 40267 98814 40323 98870
rect 40323 98814 40327 98870
rect 40263 98810 40327 98814
rect 40263 98790 40327 98794
rect 40263 98734 40267 98790
rect 40267 98734 40323 98790
rect 40323 98734 40327 98790
rect 40263 98730 40327 98734
rect 40263 98710 40327 98714
rect 40263 98654 40267 98710
rect 40267 98654 40323 98710
rect 40323 98654 40327 98710
rect 40263 98650 40327 98654
rect 40263 98630 40327 98634
rect 40263 98574 40267 98630
rect 40267 98574 40323 98630
rect 40323 98574 40327 98630
rect 40263 98570 40327 98574
rect 40263 98550 40327 98554
rect 40263 98494 40267 98550
rect 40267 98494 40323 98550
rect 40323 98494 40327 98550
rect 40263 98490 40327 98494
rect 40263 98470 40327 98474
rect 40263 98414 40267 98470
rect 40267 98414 40323 98470
rect 40323 98414 40327 98470
rect 40263 98410 40327 98414
rect 40263 98390 40327 98394
rect 40263 98334 40267 98390
rect 40267 98334 40323 98390
rect 40323 98334 40327 98390
rect 40263 98330 40327 98334
rect 40263 98310 40327 98314
rect 40263 98254 40267 98310
rect 40267 98254 40323 98310
rect 40323 98254 40327 98310
rect 40263 98250 40327 98254
rect 40263 98230 40327 98234
rect 40263 98174 40267 98230
rect 40267 98174 40323 98230
rect 40323 98174 40327 98230
rect 40263 98170 40327 98174
rect 40263 98150 40327 98154
rect 40263 98094 40267 98150
rect 40267 98094 40323 98150
rect 40323 98094 40327 98150
rect 40263 98090 40327 98094
rect 40263 98070 40327 98074
rect 40263 98014 40267 98070
rect 40267 98014 40323 98070
rect 40323 98014 40327 98070
rect 40263 98010 40327 98014
rect 40263 97990 40327 97994
rect 40263 97934 40267 97990
rect 40267 97934 40323 97990
rect 40323 97934 40327 97990
rect 40263 97930 40327 97934
rect 40263 97910 40327 97914
rect 40263 97854 40267 97910
rect 40267 97854 40323 97910
rect 40323 97854 40327 97910
rect 40263 97850 40327 97854
rect 40263 97830 40327 97834
rect 40263 97774 40267 97830
rect 40267 97774 40323 97830
rect 40323 97774 40327 97830
rect 40263 97770 40327 97774
rect 40263 97750 40327 97754
rect 40263 97694 40267 97750
rect 40267 97694 40323 97750
rect 40323 97694 40327 97750
rect 40263 97690 40327 97694
rect 40263 97670 40327 97674
rect 40263 97614 40267 97670
rect 40267 97614 40323 97670
rect 40323 97614 40327 97670
rect 40263 97610 40327 97614
rect 40263 97590 40327 97594
rect 40263 97534 40267 97590
rect 40267 97534 40323 97590
rect 40323 97534 40327 97590
rect 40263 97530 40327 97534
rect 40263 97510 40327 97514
rect 40263 97454 40267 97510
rect 40267 97454 40323 97510
rect 40323 97454 40327 97510
rect 40263 97450 40327 97454
rect 43264 100716 43328 100720
rect 43264 100660 43268 100716
rect 43268 100660 43324 100716
rect 43324 100660 43328 100716
rect 43264 100656 43328 100660
rect 43264 100636 43328 100640
rect 43264 100580 43268 100636
rect 43268 100580 43324 100636
rect 43324 100580 43328 100636
rect 43264 100576 43328 100580
rect 43264 100556 43328 100560
rect 43264 100500 43268 100556
rect 43268 100500 43324 100556
rect 43324 100500 43328 100556
rect 43264 100496 43328 100500
rect 43264 100476 43328 100480
rect 43264 100420 43268 100476
rect 43268 100420 43324 100476
rect 43324 100420 43328 100476
rect 43264 100416 43328 100420
rect 43264 100396 43328 100400
rect 43264 100340 43268 100396
rect 43268 100340 43324 100396
rect 43324 100340 43328 100396
rect 43264 100336 43328 100340
rect 43264 100316 43328 100320
rect 43264 100260 43268 100316
rect 43268 100260 43324 100316
rect 43324 100260 43328 100316
rect 43264 100256 43328 100260
rect 43264 100236 43328 100240
rect 43264 100180 43268 100236
rect 43268 100180 43324 100236
rect 43324 100180 43328 100236
rect 43264 100176 43328 100180
rect 43264 100156 43328 100160
rect 43264 100100 43268 100156
rect 43268 100100 43324 100156
rect 43324 100100 43328 100156
rect 43264 100096 43328 100100
rect 43264 100076 43328 100080
rect 43264 100020 43268 100076
rect 43268 100020 43324 100076
rect 43324 100020 43328 100076
rect 43264 100016 43328 100020
rect 43264 99996 43328 100000
rect 43264 99940 43268 99996
rect 43268 99940 43324 99996
rect 43324 99940 43328 99996
rect 43264 99936 43328 99940
rect 43264 99916 43328 99920
rect 43264 99860 43268 99916
rect 43268 99860 43324 99916
rect 43324 99860 43328 99916
rect 43264 99856 43328 99860
rect 43264 99836 43328 99840
rect 43264 99780 43268 99836
rect 43268 99780 43324 99836
rect 43324 99780 43328 99836
rect 43264 99776 43328 99780
rect 43264 99756 43328 99760
rect 43264 99700 43268 99756
rect 43268 99700 43324 99756
rect 43324 99700 43328 99756
rect 43264 99696 43328 99700
rect 43264 99676 43328 99680
rect 43264 99620 43268 99676
rect 43268 99620 43324 99676
rect 43324 99620 43328 99676
rect 43264 99616 43328 99620
rect 43264 99596 43328 99600
rect 43264 99540 43268 99596
rect 43268 99540 43324 99596
rect 43324 99540 43328 99596
rect 43264 99536 43328 99540
rect 43264 99516 43328 99520
rect 43264 99460 43268 99516
rect 43268 99460 43324 99516
rect 43324 99460 43328 99516
rect 43264 99456 43328 99460
rect 43264 99436 43328 99440
rect 43264 99380 43268 99436
rect 43268 99380 43324 99436
rect 43324 99380 43328 99436
rect 43264 99376 43328 99380
rect 43264 99356 43328 99360
rect 43264 99300 43268 99356
rect 43268 99300 43324 99356
rect 43324 99300 43328 99356
rect 43264 99296 43328 99300
rect 43264 99276 43328 99280
rect 43264 99220 43268 99276
rect 43268 99220 43324 99276
rect 43324 99220 43328 99276
rect 43264 99216 43328 99220
rect 43264 99196 43328 99200
rect 43264 99140 43268 99196
rect 43268 99140 43324 99196
rect 43324 99140 43328 99196
rect 43264 99136 43328 99140
rect 43264 99116 43328 99120
rect 43264 99060 43268 99116
rect 43268 99060 43324 99116
rect 43324 99060 43328 99116
rect 43264 99056 43328 99060
rect 43264 99036 43328 99040
rect 43264 98980 43268 99036
rect 43268 98980 43324 99036
rect 43324 98980 43328 99036
rect 43264 98976 43328 98980
rect 43264 98956 43328 98960
rect 43264 98900 43268 98956
rect 43268 98900 43324 98956
rect 43324 98900 43328 98956
rect 43264 98896 43328 98900
rect 43264 98876 43328 98880
rect 43264 98820 43268 98876
rect 43268 98820 43324 98876
rect 43324 98820 43328 98876
rect 43264 98816 43328 98820
rect 43264 98796 43328 98800
rect 43264 98740 43268 98796
rect 43268 98740 43324 98796
rect 43324 98740 43328 98796
rect 43264 98736 43328 98740
rect 43264 98716 43328 98720
rect 43264 98660 43268 98716
rect 43268 98660 43324 98716
rect 43324 98660 43328 98716
rect 43264 98656 43328 98660
rect 43264 98636 43328 98640
rect 43264 98580 43268 98636
rect 43268 98580 43324 98636
rect 43324 98580 43328 98636
rect 43264 98576 43328 98580
rect 43264 98556 43328 98560
rect 43264 98500 43268 98556
rect 43268 98500 43324 98556
rect 43324 98500 43328 98556
rect 43264 98496 43328 98500
rect 43264 98476 43328 98480
rect 43264 98420 43268 98476
rect 43268 98420 43324 98476
rect 43324 98420 43328 98476
rect 43264 98416 43328 98420
rect 43264 98396 43328 98400
rect 43264 98340 43268 98396
rect 43268 98340 43324 98396
rect 43324 98340 43328 98396
rect 43264 98336 43328 98340
rect 43264 98316 43328 98320
rect 43264 98260 43268 98316
rect 43268 98260 43324 98316
rect 43324 98260 43328 98316
rect 43264 98256 43328 98260
rect 43264 98236 43328 98240
rect 43264 98180 43268 98236
rect 43268 98180 43324 98236
rect 43324 98180 43328 98236
rect 43264 98176 43328 98180
rect 43264 98156 43328 98160
rect 43264 98100 43268 98156
rect 43268 98100 43324 98156
rect 43324 98100 43328 98156
rect 43264 98096 43328 98100
rect 43264 98076 43328 98080
rect 43264 98020 43268 98076
rect 43268 98020 43324 98076
rect 43324 98020 43328 98076
rect 43264 98016 43328 98020
rect 43264 97996 43328 98000
rect 43264 97940 43268 97996
rect 43268 97940 43324 97996
rect 43324 97940 43328 97996
rect 43264 97936 43328 97940
rect 43264 97916 43328 97920
rect 43264 97860 43268 97916
rect 43268 97860 43324 97916
rect 43324 97860 43328 97916
rect 43264 97856 43328 97860
rect 43264 97836 43328 97840
rect 43264 97780 43268 97836
rect 43268 97780 43324 97836
rect 43324 97780 43328 97836
rect 43264 97776 43328 97780
rect 43264 97756 43328 97760
rect 43264 97700 43268 97756
rect 43268 97700 43324 97756
rect 43324 97700 43328 97756
rect 43264 97696 43328 97700
rect 43264 97676 43328 97680
rect 43264 97620 43268 97676
rect 43268 97620 43324 97676
rect 43324 97620 43328 97676
rect 43264 97616 43328 97620
rect 43264 97596 43328 97600
rect 43264 97540 43268 97596
rect 43268 97540 43324 97596
rect 43324 97540 43328 97596
rect 43264 97536 43328 97540
rect 43264 97516 43328 97520
rect 43264 97460 43268 97516
rect 43268 97460 43324 97516
rect 43324 97460 43328 97516
rect 43264 97456 43328 97460
rect 68269 100696 68273 100716
rect 68273 100696 68329 100716
rect 68329 100696 68333 100716
rect 68269 100672 68333 100696
rect 68269 100652 68273 100672
rect 68273 100652 68329 100672
rect 68329 100652 68333 100672
rect 68269 100616 68273 100636
rect 68273 100616 68329 100636
rect 68329 100616 68333 100636
rect 68269 100592 68333 100616
rect 68269 100572 68273 100592
rect 68273 100572 68329 100592
rect 68329 100572 68333 100592
rect 68269 100536 68273 100556
rect 68273 100536 68329 100556
rect 68329 100536 68333 100556
rect 68269 100512 68333 100536
rect 68269 100492 68273 100512
rect 68273 100492 68329 100512
rect 68329 100492 68333 100512
rect 68269 100456 68273 100476
rect 68273 100456 68329 100476
rect 68329 100456 68333 100476
rect 68269 100432 68333 100456
rect 68269 100412 68273 100432
rect 68273 100412 68329 100432
rect 68329 100412 68333 100432
rect 68269 100376 68273 100396
rect 68273 100376 68329 100396
rect 68329 100376 68333 100396
rect 68269 100352 68333 100376
rect 68269 100332 68273 100352
rect 68273 100332 68329 100352
rect 68329 100332 68333 100352
rect 68269 100296 68273 100316
rect 68273 100296 68329 100316
rect 68329 100296 68333 100316
rect 68269 100272 68333 100296
rect 68269 100252 68273 100272
rect 68273 100252 68329 100272
rect 68329 100252 68333 100272
rect 68269 100216 68273 100236
rect 68273 100216 68329 100236
rect 68329 100216 68333 100236
rect 68269 100192 68333 100216
rect 68269 100172 68273 100192
rect 68273 100172 68329 100192
rect 68329 100172 68333 100192
rect 68269 100136 68273 100156
rect 68273 100136 68329 100156
rect 68329 100136 68333 100156
rect 68269 100112 68333 100136
rect 68269 100092 68273 100112
rect 68273 100092 68329 100112
rect 68329 100092 68333 100112
rect 68269 100056 68273 100076
rect 68273 100056 68329 100076
rect 68329 100056 68333 100076
rect 68269 100032 68333 100056
rect 68269 100012 68273 100032
rect 68273 100012 68329 100032
rect 68329 100012 68333 100032
rect 68269 99976 68273 99996
rect 68273 99976 68329 99996
rect 68329 99976 68333 99996
rect 68269 99952 68333 99976
rect 68269 99932 68273 99952
rect 68273 99932 68329 99952
rect 68329 99932 68333 99952
rect 68269 99896 68273 99916
rect 68273 99896 68329 99916
rect 68329 99896 68333 99916
rect 68269 99872 68333 99896
rect 68269 99852 68273 99872
rect 68273 99852 68329 99872
rect 68329 99852 68333 99872
rect 68269 99816 68273 99836
rect 68273 99816 68329 99836
rect 68329 99816 68333 99836
rect 68269 99792 68333 99816
rect 68269 99772 68273 99792
rect 68273 99772 68329 99792
rect 68329 99772 68333 99792
rect 68269 99736 68273 99756
rect 68273 99736 68329 99756
rect 68329 99736 68333 99756
rect 68269 99712 68333 99736
rect 68269 99692 68273 99712
rect 68273 99692 68329 99712
rect 68329 99692 68333 99712
rect 68269 99656 68273 99676
rect 68273 99656 68329 99676
rect 68329 99656 68333 99676
rect 68269 99632 68333 99656
rect 68269 99612 68273 99632
rect 68273 99612 68329 99632
rect 68329 99612 68333 99632
rect 68269 99576 68273 99596
rect 68273 99576 68329 99596
rect 68329 99576 68333 99596
rect 68269 99552 68333 99576
rect 68269 99532 68273 99552
rect 68273 99532 68329 99552
rect 68329 99532 68333 99552
rect 68269 99496 68273 99516
rect 68273 99496 68329 99516
rect 68329 99496 68333 99516
rect 68269 99472 68333 99496
rect 68269 99452 68273 99472
rect 68273 99452 68329 99472
rect 68329 99452 68333 99472
rect 68269 99416 68273 99436
rect 68273 99416 68329 99436
rect 68329 99416 68333 99436
rect 68269 99392 68333 99416
rect 68269 99372 68273 99392
rect 68273 99372 68329 99392
rect 68329 99372 68333 99392
rect 68269 99336 68273 99356
rect 68273 99336 68329 99356
rect 68329 99336 68333 99356
rect 68269 99312 68333 99336
rect 68269 99292 68273 99312
rect 68273 99292 68329 99312
rect 68329 99292 68333 99312
rect 68269 99256 68273 99276
rect 68273 99256 68329 99276
rect 68329 99256 68333 99276
rect 68269 99232 68333 99256
rect 68269 99212 68273 99232
rect 68273 99212 68329 99232
rect 68329 99212 68333 99232
rect 68269 99176 68273 99196
rect 68273 99176 68329 99196
rect 68329 99176 68333 99196
rect 68269 99152 68333 99176
rect 68269 99132 68273 99152
rect 68273 99132 68329 99152
rect 68329 99132 68333 99152
rect 68269 99096 68273 99116
rect 68273 99096 68329 99116
rect 68329 99096 68333 99116
rect 68269 99072 68333 99096
rect 68269 99052 68273 99072
rect 68273 99052 68329 99072
rect 68329 99052 68333 99072
rect 68269 99016 68273 99036
rect 68273 99016 68329 99036
rect 68329 99016 68333 99036
rect 68269 98992 68333 99016
rect 68269 98972 68273 98992
rect 68273 98972 68329 98992
rect 68329 98972 68333 98992
rect 68269 98936 68273 98956
rect 68273 98936 68329 98956
rect 68329 98936 68333 98956
rect 68269 98912 68333 98936
rect 68269 98892 68273 98912
rect 68273 98892 68329 98912
rect 68329 98892 68333 98912
rect 68269 98856 68273 98876
rect 68273 98856 68329 98876
rect 68329 98856 68333 98876
rect 68269 98832 68333 98856
rect 68269 98812 68273 98832
rect 68273 98812 68329 98832
rect 68329 98812 68333 98832
rect 68269 98776 68273 98796
rect 68273 98776 68329 98796
rect 68329 98776 68333 98796
rect 68269 98752 68333 98776
rect 68269 98732 68273 98752
rect 68273 98732 68329 98752
rect 68329 98732 68333 98752
rect 68269 98696 68273 98716
rect 68273 98696 68329 98716
rect 68329 98696 68333 98716
rect 68269 98672 68333 98696
rect 68269 98652 68273 98672
rect 68273 98652 68329 98672
rect 68329 98652 68333 98672
rect 68269 98616 68273 98636
rect 68273 98616 68329 98636
rect 68329 98616 68333 98636
rect 68269 98592 68333 98616
rect 68269 98572 68273 98592
rect 68273 98572 68329 98592
rect 68329 98572 68333 98592
rect 68269 98536 68273 98556
rect 68273 98536 68329 98556
rect 68329 98536 68333 98556
rect 68269 98512 68333 98536
rect 68269 98492 68273 98512
rect 68273 98492 68329 98512
rect 68329 98492 68333 98512
rect 68269 98456 68273 98476
rect 68273 98456 68329 98476
rect 68329 98456 68333 98476
rect 68269 98432 68333 98456
rect 68269 98412 68273 98432
rect 68273 98412 68329 98432
rect 68329 98412 68333 98432
rect 68269 98376 68273 98396
rect 68273 98376 68329 98396
rect 68329 98376 68333 98396
rect 68269 98352 68333 98376
rect 68269 98332 68273 98352
rect 68273 98332 68329 98352
rect 68329 98332 68333 98352
rect 68269 98296 68273 98316
rect 68273 98296 68329 98316
rect 68329 98296 68333 98316
rect 68269 98272 68333 98296
rect 68269 98252 68273 98272
rect 68273 98252 68329 98272
rect 68329 98252 68333 98272
rect 68269 98216 68273 98236
rect 68273 98216 68329 98236
rect 68329 98216 68333 98236
rect 68269 98192 68333 98216
rect 68269 98172 68273 98192
rect 68273 98172 68329 98192
rect 68329 98172 68333 98192
rect 68269 98136 68273 98156
rect 68273 98136 68329 98156
rect 68329 98136 68333 98156
rect 68269 98112 68333 98136
rect 68269 98092 68273 98112
rect 68273 98092 68329 98112
rect 68329 98092 68333 98112
rect 68269 98056 68273 98076
rect 68273 98056 68329 98076
rect 68329 98056 68333 98076
rect 68269 98032 68333 98056
rect 68269 98012 68273 98032
rect 68273 98012 68329 98032
rect 68329 98012 68333 98032
rect 68269 97976 68273 97996
rect 68273 97976 68329 97996
rect 68329 97976 68333 97996
rect 68269 97952 68333 97976
rect 68269 97932 68273 97952
rect 68273 97932 68329 97952
rect 68329 97932 68333 97952
rect 68269 97896 68273 97916
rect 68273 97896 68329 97916
rect 68329 97896 68333 97916
rect 68269 97872 68333 97896
rect 68269 97852 68273 97872
rect 68273 97852 68329 97872
rect 68329 97852 68333 97872
rect 68269 97816 68273 97836
rect 68273 97816 68329 97836
rect 68329 97816 68333 97836
rect 68269 97792 68333 97816
rect 68269 97772 68273 97792
rect 68273 97772 68329 97792
rect 68329 97772 68333 97792
rect 68269 97736 68273 97756
rect 68273 97736 68329 97756
rect 68329 97736 68333 97756
rect 68269 97712 68333 97736
rect 68269 97692 68273 97712
rect 68273 97692 68329 97712
rect 68329 97692 68333 97712
rect 68269 97656 68273 97676
rect 68273 97656 68329 97676
rect 68329 97656 68333 97676
rect 68269 97632 68333 97656
rect 68269 97612 68273 97632
rect 68273 97612 68329 97632
rect 68329 97612 68333 97632
rect 68269 97576 68273 97596
rect 68273 97576 68329 97596
rect 68329 97576 68333 97596
rect 68269 97552 68333 97576
rect 68269 97532 68273 97552
rect 68273 97532 68329 97552
rect 68329 97532 68333 97552
rect 68269 97496 68273 97516
rect 68273 97496 68329 97516
rect 68329 97496 68333 97516
rect 68269 97472 68333 97496
rect 68269 97452 68273 97472
rect 68273 97452 68329 97472
rect 68329 97452 68333 97472
rect 71270 100709 71274 100729
rect 71274 100709 71330 100729
rect 71330 100709 71334 100729
rect 71270 100685 71334 100709
rect 71270 100665 71274 100685
rect 71274 100665 71330 100685
rect 71330 100665 71334 100685
rect 71270 100629 71274 100649
rect 71274 100629 71330 100649
rect 71330 100629 71334 100649
rect 71270 100605 71334 100629
rect 71270 100585 71274 100605
rect 71274 100585 71330 100605
rect 71330 100585 71334 100605
rect 71270 100549 71274 100569
rect 71274 100549 71330 100569
rect 71330 100549 71334 100569
rect 71270 100525 71334 100549
rect 71270 100505 71274 100525
rect 71274 100505 71330 100525
rect 71330 100505 71334 100525
rect 71270 100469 71274 100489
rect 71274 100469 71330 100489
rect 71330 100469 71334 100489
rect 71270 100445 71334 100469
rect 71270 100425 71274 100445
rect 71274 100425 71330 100445
rect 71330 100425 71334 100445
rect 71270 100389 71274 100409
rect 71274 100389 71330 100409
rect 71330 100389 71334 100409
rect 71270 100365 71334 100389
rect 71270 100345 71274 100365
rect 71274 100345 71330 100365
rect 71330 100345 71334 100365
rect 71270 100309 71274 100329
rect 71274 100309 71330 100329
rect 71330 100309 71334 100329
rect 71270 100285 71334 100309
rect 71270 100265 71274 100285
rect 71274 100265 71330 100285
rect 71330 100265 71334 100285
rect 71270 100229 71274 100249
rect 71274 100229 71330 100249
rect 71330 100229 71334 100249
rect 71270 100205 71334 100229
rect 71270 100185 71274 100205
rect 71274 100185 71330 100205
rect 71330 100185 71334 100205
rect 71270 100149 71274 100169
rect 71274 100149 71330 100169
rect 71330 100149 71334 100169
rect 71270 100125 71334 100149
rect 71270 100105 71274 100125
rect 71274 100105 71330 100125
rect 71330 100105 71334 100125
rect 71270 100069 71274 100089
rect 71274 100069 71330 100089
rect 71330 100069 71334 100089
rect 71270 100045 71334 100069
rect 71270 100025 71274 100045
rect 71274 100025 71330 100045
rect 71330 100025 71334 100045
rect 71270 99989 71274 100009
rect 71274 99989 71330 100009
rect 71330 99989 71334 100009
rect 71270 99965 71334 99989
rect 71270 99945 71274 99965
rect 71274 99945 71330 99965
rect 71330 99945 71334 99965
rect 71270 99909 71274 99929
rect 71274 99909 71330 99929
rect 71330 99909 71334 99929
rect 71270 99885 71334 99909
rect 71270 99865 71274 99885
rect 71274 99865 71330 99885
rect 71330 99865 71334 99885
rect 71270 99829 71274 99849
rect 71274 99829 71330 99849
rect 71330 99829 71334 99849
rect 71270 99805 71334 99829
rect 71270 99785 71274 99805
rect 71274 99785 71330 99805
rect 71330 99785 71334 99805
rect 71270 99749 71274 99769
rect 71274 99749 71330 99769
rect 71330 99749 71334 99769
rect 71270 99725 71334 99749
rect 71270 99705 71274 99725
rect 71274 99705 71330 99725
rect 71330 99705 71334 99725
rect 71270 99669 71274 99689
rect 71274 99669 71330 99689
rect 71330 99669 71334 99689
rect 71270 99645 71334 99669
rect 71270 99625 71274 99645
rect 71274 99625 71330 99645
rect 71330 99625 71334 99645
rect 71270 99589 71274 99609
rect 71274 99589 71330 99609
rect 71330 99589 71334 99609
rect 71270 99565 71334 99589
rect 71270 99545 71274 99565
rect 71274 99545 71330 99565
rect 71330 99545 71334 99565
rect 71270 99509 71274 99529
rect 71274 99509 71330 99529
rect 71330 99509 71334 99529
rect 71270 99485 71334 99509
rect 71270 99465 71274 99485
rect 71274 99465 71330 99485
rect 71330 99465 71334 99485
rect 71270 99429 71274 99449
rect 71274 99429 71330 99449
rect 71330 99429 71334 99449
rect 71270 99405 71334 99429
rect 71270 99385 71274 99405
rect 71274 99385 71330 99405
rect 71330 99385 71334 99405
rect 71270 99349 71274 99369
rect 71274 99349 71330 99369
rect 71330 99349 71334 99369
rect 71270 99325 71334 99349
rect 71270 99305 71274 99325
rect 71274 99305 71330 99325
rect 71330 99305 71334 99325
rect 71270 99269 71274 99289
rect 71274 99269 71330 99289
rect 71330 99269 71334 99289
rect 71270 99245 71334 99269
rect 71270 99225 71274 99245
rect 71274 99225 71330 99245
rect 71330 99225 71334 99245
rect 71270 99189 71274 99209
rect 71274 99189 71330 99209
rect 71330 99189 71334 99209
rect 71270 99165 71334 99189
rect 71270 99145 71274 99165
rect 71274 99145 71330 99165
rect 71330 99145 71334 99165
rect 71270 99109 71274 99129
rect 71274 99109 71330 99129
rect 71330 99109 71334 99129
rect 71270 99085 71334 99109
rect 71270 99065 71274 99085
rect 71274 99065 71330 99085
rect 71330 99065 71334 99085
rect 71270 99029 71274 99049
rect 71274 99029 71330 99049
rect 71330 99029 71334 99049
rect 71270 99005 71334 99029
rect 71270 98985 71274 99005
rect 71274 98985 71330 99005
rect 71330 98985 71334 99005
rect 71270 98949 71274 98969
rect 71274 98949 71330 98969
rect 71330 98949 71334 98969
rect 71270 98925 71334 98949
rect 71270 98905 71274 98925
rect 71274 98905 71330 98925
rect 71330 98905 71334 98925
rect 71270 98869 71274 98889
rect 71274 98869 71330 98889
rect 71330 98869 71334 98889
rect 71270 98845 71334 98869
rect 71270 98825 71274 98845
rect 71274 98825 71330 98845
rect 71330 98825 71334 98845
rect 71270 98789 71274 98809
rect 71274 98789 71330 98809
rect 71330 98789 71334 98809
rect 71270 98765 71334 98789
rect 71270 98745 71274 98765
rect 71274 98745 71330 98765
rect 71330 98745 71334 98765
rect 71270 98709 71274 98729
rect 71274 98709 71330 98729
rect 71330 98709 71334 98729
rect 71270 98685 71334 98709
rect 71270 98665 71274 98685
rect 71274 98665 71330 98685
rect 71330 98665 71334 98685
rect 71270 98629 71274 98649
rect 71274 98629 71330 98649
rect 71330 98629 71334 98649
rect 71270 98605 71334 98629
rect 71270 98585 71274 98605
rect 71274 98585 71330 98605
rect 71330 98585 71334 98605
rect 71270 98549 71274 98569
rect 71274 98549 71330 98569
rect 71330 98549 71334 98569
rect 71270 98525 71334 98549
rect 71270 98505 71274 98525
rect 71274 98505 71330 98525
rect 71330 98505 71334 98525
rect 71270 98469 71274 98489
rect 71274 98469 71330 98489
rect 71330 98469 71334 98489
rect 71270 98445 71334 98469
rect 71270 98425 71274 98445
rect 71274 98425 71330 98445
rect 71330 98425 71334 98445
rect 71270 98389 71274 98409
rect 71274 98389 71330 98409
rect 71330 98389 71334 98409
rect 71270 98365 71334 98389
rect 71270 98345 71274 98365
rect 71274 98345 71330 98365
rect 71330 98345 71334 98365
rect 71270 98309 71274 98329
rect 71274 98309 71330 98329
rect 71330 98309 71334 98329
rect 71270 98285 71334 98309
rect 71270 98265 71274 98285
rect 71274 98265 71330 98285
rect 71330 98265 71334 98285
rect 71270 98229 71274 98249
rect 71274 98229 71330 98249
rect 71330 98229 71334 98249
rect 71270 98205 71334 98229
rect 71270 98185 71274 98205
rect 71274 98185 71330 98205
rect 71330 98185 71334 98205
rect 71270 98149 71274 98169
rect 71274 98149 71330 98169
rect 71330 98149 71334 98169
rect 71270 98125 71334 98149
rect 71270 98105 71274 98125
rect 71274 98105 71330 98125
rect 71330 98105 71334 98125
rect 71270 98069 71274 98089
rect 71274 98069 71330 98089
rect 71330 98069 71334 98089
rect 71270 98045 71334 98069
rect 71270 98025 71274 98045
rect 71274 98025 71330 98045
rect 71330 98025 71334 98045
rect 71270 97989 71274 98009
rect 71274 97989 71330 98009
rect 71330 97989 71334 98009
rect 71270 97965 71334 97989
rect 71270 97945 71274 97965
rect 71274 97945 71330 97965
rect 71330 97945 71334 97965
rect 71270 97909 71274 97929
rect 71274 97909 71330 97929
rect 71330 97909 71334 97929
rect 71270 97885 71334 97909
rect 71270 97865 71274 97885
rect 71274 97865 71330 97885
rect 71330 97865 71334 97885
rect 71270 97829 71274 97849
rect 71274 97829 71330 97849
rect 71330 97829 71334 97849
rect 71270 97805 71334 97829
rect 71270 97785 71274 97805
rect 71274 97785 71330 97805
rect 71330 97785 71334 97805
rect 71270 97749 71274 97769
rect 71274 97749 71330 97769
rect 71330 97749 71334 97769
rect 71270 97725 71334 97749
rect 71270 97705 71274 97725
rect 71274 97705 71330 97725
rect 71330 97705 71334 97725
rect 71270 97669 71274 97689
rect 71274 97669 71330 97689
rect 71330 97669 71334 97689
rect 71270 97645 71334 97669
rect 71270 97625 71274 97645
rect 71274 97625 71330 97645
rect 71330 97625 71334 97645
rect 71270 97589 71274 97609
rect 71274 97589 71330 97609
rect 71330 97589 71334 97609
rect 71270 97565 71334 97589
rect 71270 97545 71274 97565
rect 71274 97545 71330 97565
rect 71330 97545 71334 97565
rect 71270 97509 71274 97529
rect 71274 97509 71330 97529
rect 71330 97509 71334 97529
rect 71270 97485 71334 97509
rect 71270 97465 71274 97485
rect 71274 97465 71330 97485
rect 71330 97465 71334 97485
rect 40430 95820 40494 95824
rect 40430 95764 40434 95820
rect 40434 95764 40490 95820
rect 40490 95764 40494 95820
rect 40430 95760 40494 95764
rect 41608 95816 41672 95820
rect 41608 95760 41612 95816
rect 41612 95760 41668 95816
rect 41668 95760 41672 95816
rect 41608 95756 41672 95760
rect 41825 95823 41889 95827
rect 41825 95767 41829 95823
rect 41829 95767 41885 95823
rect 41885 95767 41889 95823
rect 41825 95763 41889 95767
rect 42959 95820 43023 95824
rect 42959 95764 42963 95820
rect 42963 95764 43019 95820
rect 43019 95764 43023 95820
rect 42959 95760 43023 95764
rect 40540 94316 40604 94320
rect 40540 94260 40544 94316
rect 40544 94260 40600 94316
rect 40600 94260 40604 94316
rect 40540 94256 40604 94260
rect 41654 94302 41718 94306
rect 41654 94246 41658 94302
rect 41658 94246 41714 94302
rect 41714 94246 41718 94302
rect 41654 94242 41718 94246
rect 41867 94303 41931 94307
rect 41867 94247 41871 94303
rect 41871 94247 41927 94303
rect 41927 94247 41931 94303
rect 41867 94243 41931 94247
rect 43031 94303 43095 94307
rect 43031 94247 43035 94303
rect 43035 94247 43091 94303
rect 43091 94247 43095 94303
rect 43031 94243 43095 94247
rect 93725 93292 93789 93356
rect 93160 92699 93224 92763
rect 41672 92510 41736 92514
rect 41672 92454 41676 92510
rect 41676 92454 41732 92510
rect 41732 92454 41736 92510
rect 41672 92450 41736 92454
rect 41672 92430 41736 92434
rect 41672 92374 41676 92430
rect 41676 92374 41732 92430
rect 41732 92374 41736 92430
rect 41672 92370 41736 92374
rect 41672 92350 41736 92354
rect 41672 92294 41676 92350
rect 41676 92294 41732 92350
rect 41732 92294 41736 92350
rect 41672 92290 41736 92294
rect 41135 92273 41199 92277
rect 41135 92217 41139 92273
rect 41139 92217 41195 92273
rect 41195 92217 41199 92273
rect 41135 92213 41199 92217
rect 41135 92193 41199 92197
rect 41135 92137 41139 92193
rect 41139 92137 41195 92193
rect 41195 92137 41199 92193
rect 41135 92133 41199 92137
rect 41672 92270 41736 92274
rect 41672 92214 41676 92270
rect 41676 92214 41732 92270
rect 41732 92214 41736 92270
rect 41672 92210 41736 92214
rect 42219 92276 42283 92280
rect 42219 92220 42223 92276
rect 42223 92220 42279 92276
rect 42279 92220 42283 92276
rect 42219 92216 42283 92220
rect 42219 92196 42283 92200
rect 42219 92140 42223 92196
rect 42223 92140 42279 92196
rect 42279 92140 42283 92196
rect 42219 92136 42283 92140
rect 92571 92039 92635 92103
rect 40517 91631 40581 91635
rect 40517 91575 40521 91631
rect 40521 91575 40577 91631
rect 40577 91575 40581 91631
rect 40517 91571 40581 91575
rect 41672 91625 41736 91629
rect 41672 91569 41676 91625
rect 41676 91569 41732 91625
rect 41732 91569 41736 91625
rect 41672 91565 41736 91569
rect 42790 91636 42854 91640
rect 42790 91580 42794 91636
rect 42794 91580 42850 91636
rect 42850 91580 42854 91636
rect 42790 91576 42854 91580
rect 43998 90727 44062 90791
rect 49021 90727 49085 90791
rect 44779 90404 44843 90468
rect 49828 90404 49892 90468
rect 45789 89971 45853 90035
rect 54421 89971 54485 90035
rect 46558 89718 46622 89782
rect 55228 89718 55292 89782
rect 49021 89287 49085 89351
rect 54421 89287 54485 89351
rect 49828 89034 49892 89098
rect 55228 89034 55292 89098
rect 74525 88746 74589 88750
rect 74525 88690 74529 88746
rect 74529 88690 74585 88746
rect 74585 88690 74589 88746
rect 74525 88686 74589 88690
rect 74525 88666 74589 88670
rect 74525 88610 74529 88666
rect 74529 88610 74585 88666
rect 74585 88610 74589 88666
rect 74525 88606 74589 88610
rect 74525 88586 74589 88590
rect 74525 88530 74529 88586
rect 74529 88530 74585 88586
rect 74585 88530 74589 88586
rect 74525 88526 74589 88530
rect 74525 88506 74589 88510
rect 74525 88450 74529 88506
rect 74529 88450 74585 88506
rect 74585 88450 74589 88506
rect 74525 88446 74589 88450
rect 74525 88426 74589 88430
rect 74525 88370 74529 88426
rect 74529 88370 74585 88426
rect 74585 88370 74589 88426
rect 74525 88366 74589 88370
rect 74525 88346 74589 88350
rect 74525 88290 74529 88346
rect 74529 88290 74585 88346
rect 74585 88290 74589 88346
rect 74525 88286 74589 88290
rect 74525 88266 74589 88270
rect 74525 88210 74529 88266
rect 74529 88210 74585 88266
rect 74585 88210 74589 88266
rect 74525 88206 74589 88210
rect 81053 88746 81117 88750
rect 81053 88690 81057 88746
rect 81057 88690 81113 88746
rect 81113 88690 81117 88746
rect 81053 88686 81117 88690
rect 81053 88666 81117 88670
rect 81053 88610 81057 88666
rect 81057 88610 81113 88666
rect 81113 88610 81117 88666
rect 81053 88606 81117 88610
rect 81053 88586 81117 88590
rect 81053 88530 81057 88586
rect 81057 88530 81113 88586
rect 81113 88530 81117 88586
rect 81053 88526 81117 88530
rect 81053 88506 81117 88510
rect 81053 88450 81057 88506
rect 81057 88450 81113 88506
rect 81113 88450 81117 88506
rect 81053 88446 81117 88450
rect 81053 88426 81117 88430
rect 81053 88370 81057 88426
rect 81057 88370 81113 88426
rect 81113 88370 81117 88426
rect 81053 88366 81117 88370
rect 81053 88346 81117 88350
rect 81053 88290 81057 88346
rect 81057 88290 81113 88346
rect 81113 88290 81117 88346
rect 81053 88286 81117 88290
rect 81053 88266 81117 88270
rect 81053 88210 81057 88266
rect 81057 88210 81113 88266
rect 81113 88210 81117 88266
rect 81053 88206 81117 88210
rect 88669 88746 88733 88750
rect 88669 88690 88673 88746
rect 88673 88690 88729 88746
rect 88729 88690 88733 88746
rect 88669 88686 88733 88690
rect 88669 88666 88733 88670
rect 88669 88610 88673 88666
rect 88673 88610 88729 88666
rect 88729 88610 88733 88666
rect 88669 88606 88733 88610
rect 88669 88586 88733 88590
rect 88669 88530 88673 88586
rect 88673 88530 88729 88586
rect 88729 88530 88733 88586
rect 88669 88526 88733 88530
rect 88669 88506 88733 88510
rect 88669 88450 88673 88506
rect 88673 88450 88729 88506
rect 88729 88450 88733 88506
rect 88669 88446 88733 88450
rect 88669 88426 88733 88430
rect 88669 88370 88673 88426
rect 88673 88370 88729 88426
rect 88729 88370 88733 88426
rect 88669 88366 88733 88370
rect 88669 88346 88733 88350
rect 88669 88290 88673 88346
rect 88673 88290 88729 88346
rect 88729 88290 88733 88346
rect 88669 88286 88733 88290
rect 88669 88266 88733 88270
rect 88669 88210 88673 88266
rect 88673 88210 88729 88266
rect 88729 88210 88733 88266
rect 88669 88206 88733 88210
rect 46038 87251 46342 87555
rect 46907 87360 46971 87424
rect 47239 87420 47303 87424
rect 47239 87364 47243 87420
rect 47243 87364 47299 87420
rect 47299 87364 47303 87420
rect 47239 87360 47303 87364
rect 47319 87420 47383 87424
rect 47319 87364 47323 87420
rect 47323 87364 47379 87420
rect 47379 87364 47383 87420
rect 47319 87360 47383 87364
rect 47399 87420 47463 87424
rect 47399 87364 47403 87420
rect 47403 87364 47459 87420
rect 47459 87364 47463 87420
rect 47399 87360 47463 87364
rect 47479 87420 47543 87424
rect 47479 87364 47483 87420
rect 47483 87364 47539 87420
rect 47539 87364 47543 87420
rect 47479 87360 47543 87364
rect 47559 87420 47623 87424
rect 47559 87364 47563 87420
rect 47563 87364 47619 87420
rect 47619 87364 47623 87420
rect 47559 87360 47623 87364
rect 49050 87422 49114 87426
rect 49050 87366 49054 87422
rect 49054 87366 49110 87422
rect 49110 87366 49114 87422
rect 49050 87362 49114 87366
rect 49130 87422 49194 87426
rect 49130 87366 49134 87422
rect 49134 87366 49190 87422
rect 49190 87366 49194 87422
rect 49130 87362 49194 87366
rect 49210 87422 49274 87426
rect 49210 87366 49214 87422
rect 49214 87366 49270 87422
rect 49270 87366 49274 87422
rect 49210 87362 49274 87366
rect 49290 87422 49354 87426
rect 49290 87366 49294 87422
rect 49294 87366 49350 87422
rect 49350 87366 49354 87422
rect 49290 87362 49354 87366
rect 49370 87422 49434 87426
rect 49370 87366 49374 87422
rect 49374 87366 49430 87422
rect 49430 87366 49434 87422
rect 49370 87362 49434 87366
rect 50845 87418 50909 87422
rect 50845 87362 50849 87418
rect 50849 87362 50905 87418
rect 50905 87362 50909 87418
rect 50845 87358 50909 87362
rect 50925 87418 50989 87422
rect 50925 87362 50929 87418
rect 50929 87362 50985 87418
rect 50985 87362 50989 87418
rect 50925 87358 50989 87362
rect 51005 87418 51069 87422
rect 51005 87362 51009 87418
rect 51009 87362 51065 87418
rect 51065 87362 51069 87418
rect 51005 87358 51069 87362
rect 51085 87418 51149 87422
rect 51085 87362 51089 87418
rect 51089 87362 51145 87418
rect 51145 87362 51149 87418
rect 51085 87358 51149 87362
rect 51165 87418 51229 87422
rect 51165 87362 51169 87418
rect 51169 87362 51225 87418
rect 51225 87362 51229 87418
rect 51165 87358 51229 87362
rect 52644 87416 52708 87420
rect 52644 87360 52648 87416
rect 52648 87360 52704 87416
rect 52704 87360 52708 87416
rect 52644 87356 52708 87360
rect 52724 87416 52788 87420
rect 52724 87360 52728 87416
rect 52728 87360 52784 87416
rect 52784 87360 52788 87416
rect 52724 87356 52788 87360
rect 52804 87416 52868 87420
rect 52804 87360 52808 87416
rect 52808 87360 52864 87416
rect 52864 87360 52868 87416
rect 52804 87356 52868 87360
rect 52884 87416 52948 87420
rect 52884 87360 52888 87416
rect 52888 87360 52944 87416
rect 52944 87360 52948 87416
rect 52884 87356 52948 87360
rect 52964 87416 53028 87420
rect 52964 87360 52968 87416
rect 52968 87360 53024 87416
rect 53024 87360 53028 87416
rect 52964 87356 53028 87360
rect 54435 87420 54499 87424
rect 54435 87364 54439 87420
rect 54439 87364 54495 87420
rect 54495 87364 54499 87420
rect 54435 87360 54499 87364
rect 54515 87420 54579 87424
rect 54515 87364 54519 87420
rect 54519 87364 54575 87420
rect 54575 87364 54579 87420
rect 54515 87360 54579 87364
rect 54595 87420 54659 87424
rect 54595 87364 54599 87420
rect 54599 87364 54655 87420
rect 54655 87364 54659 87420
rect 54595 87360 54659 87364
rect 54675 87420 54739 87424
rect 54675 87364 54679 87420
rect 54679 87364 54735 87420
rect 54735 87364 54739 87420
rect 54675 87360 54739 87364
rect 54755 87420 54819 87424
rect 54755 87364 54759 87420
rect 54759 87364 54815 87420
rect 54815 87364 54819 87420
rect 54755 87360 54819 87364
rect 56237 87416 56301 87420
rect 56237 87360 56241 87416
rect 56241 87360 56297 87416
rect 56297 87360 56301 87416
rect 56237 87356 56301 87360
rect 56317 87416 56381 87420
rect 56317 87360 56321 87416
rect 56321 87360 56377 87416
rect 56377 87360 56381 87416
rect 56317 87356 56381 87360
rect 56397 87416 56461 87420
rect 56397 87360 56401 87416
rect 56401 87360 56457 87416
rect 56457 87360 56461 87416
rect 56397 87356 56461 87360
rect 56477 87416 56541 87420
rect 56477 87360 56481 87416
rect 56481 87360 56537 87416
rect 56537 87360 56541 87416
rect 56477 87356 56541 87360
rect 56557 87416 56621 87420
rect 56557 87360 56561 87416
rect 56561 87360 56617 87416
rect 56617 87360 56621 87416
rect 56557 87356 56621 87360
rect 50163 87216 50387 87220
rect 50163 87000 50167 87216
rect 50167 87000 50383 87216
rect 50383 87000 50387 87216
rect 50163 86996 50387 87000
rect 57884 87242 58348 87246
rect 57884 87026 57888 87242
rect 57888 87026 58344 87242
rect 58344 87026 58348 87242
rect 57884 87022 58348 87026
rect 75070 86743 75134 86747
rect 75070 86687 75074 86743
rect 75074 86687 75130 86743
rect 75130 86687 75134 86743
rect 75070 86683 75134 86687
rect 75070 86663 75134 86667
rect 75070 86607 75074 86663
rect 75074 86607 75130 86663
rect 75130 86607 75134 86663
rect 75070 86603 75134 86607
rect 75070 86583 75134 86587
rect 75070 86527 75074 86583
rect 75074 86527 75130 86583
rect 75130 86527 75134 86583
rect 75070 86523 75134 86527
rect 75070 86503 75134 86507
rect 75070 86447 75074 86503
rect 75074 86447 75130 86503
rect 75130 86447 75134 86503
rect 75070 86443 75134 86447
rect 75070 86423 75134 86427
rect 75070 86367 75074 86423
rect 75074 86367 75130 86423
rect 75130 86367 75134 86423
rect 75070 86363 75134 86367
rect 75070 86343 75134 86347
rect 75070 86287 75074 86343
rect 75074 86287 75130 86343
rect 75130 86287 75134 86343
rect 75070 86283 75134 86287
rect 75070 86263 75134 86267
rect 75070 86207 75074 86263
rect 75074 86207 75130 86263
rect 75130 86207 75134 86263
rect 75070 86203 75134 86207
rect 76158 86743 76222 86747
rect 76158 86687 76162 86743
rect 76162 86687 76218 86743
rect 76218 86687 76222 86743
rect 76158 86683 76222 86687
rect 76158 86663 76222 86667
rect 76158 86607 76162 86663
rect 76162 86607 76218 86663
rect 76218 86607 76222 86663
rect 76158 86603 76222 86607
rect 76158 86583 76222 86587
rect 76158 86527 76162 86583
rect 76162 86527 76218 86583
rect 76218 86527 76222 86583
rect 76158 86523 76222 86527
rect 76158 86503 76222 86507
rect 76158 86447 76162 86503
rect 76162 86447 76218 86503
rect 76218 86447 76222 86503
rect 76158 86443 76222 86447
rect 76158 86423 76222 86427
rect 76158 86367 76162 86423
rect 76162 86367 76218 86423
rect 76218 86367 76222 86423
rect 76158 86363 76222 86367
rect 76158 86343 76222 86347
rect 76158 86287 76162 86343
rect 76162 86287 76218 86343
rect 76218 86287 76222 86343
rect 76158 86283 76222 86287
rect 76158 86263 76222 86267
rect 76158 86207 76162 86263
rect 76162 86207 76218 86263
rect 76218 86207 76222 86263
rect 76158 86203 76222 86207
rect 78334 86743 78398 86747
rect 78334 86687 78338 86743
rect 78338 86687 78394 86743
rect 78394 86687 78398 86743
rect 78334 86683 78398 86687
rect 78334 86663 78398 86667
rect 78334 86607 78338 86663
rect 78338 86607 78394 86663
rect 78394 86607 78398 86663
rect 78334 86603 78398 86607
rect 78334 86583 78398 86587
rect 78334 86527 78338 86583
rect 78338 86527 78394 86583
rect 78394 86527 78398 86583
rect 78334 86523 78398 86527
rect 78334 86503 78398 86507
rect 78334 86447 78338 86503
rect 78338 86447 78394 86503
rect 78394 86447 78398 86503
rect 78334 86443 78398 86447
rect 78334 86423 78398 86427
rect 78334 86367 78338 86423
rect 78338 86367 78394 86423
rect 78394 86367 78398 86423
rect 78334 86363 78398 86367
rect 78334 86343 78398 86347
rect 78334 86287 78338 86343
rect 78338 86287 78394 86343
rect 78394 86287 78398 86343
rect 78334 86283 78398 86287
rect 78334 86263 78398 86267
rect 78334 86207 78338 86263
rect 78338 86207 78394 86263
rect 78394 86207 78398 86263
rect 78334 86203 78398 86207
rect 79422 86743 79486 86747
rect 79422 86687 79426 86743
rect 79426 86687 79482 86743
rect 79482 86687 79486 86743
rect 79422 86683 79486 86687
rect 79422 86663 79486 86667
rect 79422 86607 79426 86663
rect 79426 86607 79482 86663
rect 79482 86607 79486 86663
rect 79422 86603 79486 86607
rect 79422 86583 79486 86587
rect 79422 86527 79426 86583
rect 79426 86527 79482 86583
rect 79482 86527 79486 86583
rect 79422 86523 79486 86527
rect 79422 86503 79486 86507
rect 79422 86447 79426 86503
rect 79426 86447 79482 86503
rect 79482 86447 79486 86503
rect 79422 86443 79486 86447
rect 79422 86423 79486 86427
rect 79422 86367 79426 86423
rect 79426 86367 79482 86423
rect 79482 86367 79486 86423
rect 79422 86363 79486 86367
rect 79422 86343 79486 86347
rect 79422 86287 79426 86343
rect 79426 86287 79482 86343
rect 79482 86287 79486 86343
rect 79422 86283 79486 86287
rect 79422 86263 79486 86267
rect 79422 86207 79426 86263
rect 79426 86207 79482 86263
rect 79482 86207 79486 86263
rect 79422 86203 79486 86207
rect 80510 86743 80574 86747
rect 80510 86687 80514 86743
rect 80514 86687 80570 86743
rect 80570 86687 80574 86743
rect 80510 86683 80574 86687
rect 80510 86663 80574 86667
rect 80510 86607 80514 86663
rect 80514 86607 80570 86663
rect 80570 86607 80574 86663
rect 80510 86603 80574 86607
rect 80510 86583 80574 86587
rect 80510 86527 80514 86583
rect 80514 86527 80570 86583
rect 80570 86527 80574 86583
rect 80510 86523 80574 86527
rect 80510 86503 80574 86507
rect 80510 86447 80514 86503
rect 80514 86447 80570 86503
rect 80570 86447 80574 86503
rect 80510 86443 80574 86447
rect 80510 86423 80574 86427
rect 80510 86367 80514 86423
rect 80514 86367 80570 86423
rect 80570 86367 80574 86423
rect 80510 86363 80574 86367
rect 80510 86343 80574 86347
rect 80510 86287 80514 86343
rect 80514 86287 80570 86343
rect 80570 86287 80574 86343
rect 80510 86283 80574 86287
rect 80510 86263 80574 86267
rect 80510 86207 80514 86263
rect 80514 86207 80570 86263
rect 80570 86207 80574 86263
rect 80510 86203 80574 86207
rect 81598 86743 81662 86747
rect 81598 86687 81602 86743
rect 81602 86687 81658 86743
rect 81658 86687 81662 86743
rect 81598 86683 81662 86687
rect 81598 86663 81662 86667
rect 81598 86607 81602 86663
rect 81602 86607 81658 86663
rect 81658 86607 81662 86663
rect 81598 86603 81662 86607
rect 81598 86583 81662 86587
rect 81598 86527 81602 86583
rect 81602 86527 81658 86583
rect 81658 86527 81662 86583
rect 81598 86523 81662 86527
rect 81598 86503 81662 86507
rect 81598 86447 81602 86503
rect 81602 86447 81658 86503
rect 81658 86447 81662 86503
rect 81598 86443 81662 86447
rect 81598 86423 81662 86427
rect 81598 86367 81602 86423
rect 81602 86367 81658 86423
rect 81658 86367 81662 86423
rect 81598 86363 81662 86367
rect 81598 86343 81662 86347
rect 81598 86287 81602 86343
rect 81602 86287 81658 86343
rect 81658 86287 81662 86343
rect 81598 86283 81662 86287
rect 81598 86263 81662 86267
rect 81598 86207 81602 86263
rect 81602 86207 81658 86263
rect 81658 86207 81662 86263
rect 81598 86203 81662 86207
rect 82686 86743 82750 86747
rect 82686 86687 82690 86743
rect 82690 86687 82746 86743
rect 82746 86687 82750 86743
rect 82686 86683 82750 86687
rect 82686 86663 82750 86667
rect 82686 86607 82690 86663
rect 82690 86607 82746 86663
rect 82746 86607 82750 86663
rect 82686 86603 82750 86607
rect 82686 86583 82750 86587
rect 82686 86527 82690 86583
rect 82690 86527 82746 86583
rect 82746 86527 82750 86583
rect 82686 86523 82750 86527
rect 82686 86503 82750 86507
rect 82686 86447 82690 86503
rect 82690 86447 82746 86503
rect 82746 86447 82750 86503
rect 82686 86443 82750 86447
rect 82686 86423 82750 86427
rect 82686 86367 82690 86423
rect 82690 86367 82746 86423
rect 82746 86367 82750 86423
rect 82686 86363 82750 86367
rect 82686 86343 82750 86347
rect 82686 86287 82690 86343
rect 82690 86287 82746 86343
rect 82746 86287 82750 86343
rect 82686 86283 82750 86287
rect 82686 86263 82750 86267
rect 82686 86207 82690 86263
rect 82690 86207 82746 86263
rect 82746 86207 82750 86263
rect 82686 86203 82750 86207
rect 83774 86743 83838 86747
rect 83774 86687 83778 86743
rect 83778 86687 83834 86743
rect 83834 86687 83838 86743
rect 83774 86683 83838 86687
rect 83774 86663 83838 86667
rect 83774 86607 83778 86663
rect 83778 86607 83834 86663
rect 83834 86607 83838 86663
rect 83774 86603 83838 86607
rect 83774 86583 83838 86587
rect 83774 86527 83778 86583
rect 83778 86527 83834 86583
rect 83834 86527 83838 86583
rect 83774 86523 83838 86527
rect 83774 86503 83838 86507
rect 83774 86447 83778 86503
rect 83778 86447 83834 86503
rect 83834 86447 83838 86503
rect 83774 86443 83838 86447
rect 83774 86423 83838 86427
rect 83774 86367 83778 86423
rect 83778 86367 83834 86423
rect 83834 86367 83838 86423
rect 83774 86363 83838 86367
rect 83774 86343 83838 86347
rect 83774 86287 83778 86343
rect 83778 86287 83834 86343
rect 83834 86287 83838 86343
rect 83774 86283 83838 86287
rect 83774 86263 83838 86267
rect 83774 86207 83778 86263
rect 83778 86207 83834 86263
rect 83834 86207 83838 86263
rect 83774 86203 83838 86207
rect 85950 86743 86014 86747
rect 85950 86687 85954 86743
rect 85954 86687 86010 86743
rect 86010 86687 86014 86743
rect 85950 86683 86014 86687
rect 85950 86663 86014 86667
rect 85950 86607 85954 86663
rect 85954 86607 86010 86663
rect 86010 86607 86014 86663
rect 85950 86603 86014 86607
rect 85950 86583 86014 86587
rect 85950 86527 85954 86583
rect 85954 86527 86010 86583
rect 86010 86527 86014 86583
rect 85950 86523 86014 86527
rect 85950 86503 86014 86507
rect 85950 86447 85954 86503
rect 85954 86447 86010 86503
rect 86010 86447 86014 86503
rect 85950 86443 86014 86447
rect 85950 86423 86014 86427
rect 85950 86367 85954 86423
rect 85954 86367 86010 86423
rect 86010 86367 86014 86423
rect 85950 86363 86014 86367
rect 85950 86343 86014 86347
rect 85950 86287 85954 86343
rect 85954 86287 86010 86343
rect 86010 86287 86014 86343
rect 85950 86283 86014 86287
rect 85950 86263 86014 86267
rect 85950 86207 85954 86263
rect 85954 86207 86010 86263
rect 86010 86207 86014 86263
rect 85950 86203 86014 86207
rect 87038 86743 87102 86747
rect 87038 86687 87042 86743
rect 87042 86687 87098 86743
rect 87098 86687 87102 86743
rect 87038 86683 87102 86687
rect 87038 86663 87102 86667
rect 87038 86607 87042 86663
rect 87042 86607 87098 86663
rect 87098 86607 87102 86663
rect 87038 86603 87102 86607
rect 87038 86583 87102 86587
rect 87038 86527 87042 86583
rect 87042 86527 87098 86583
rect 87098 86527 87102 86583
rect 87038 86523 87102 86527
rect 87038 86503 87102 86507
rect 87038 86447 87042 86503
rect 87042 86447 87098 86503
rect 87098 86447 87102 86503
rect 87038 86443 87102 86447
rect 87038 86423 87102 86427
rect 87038 86367 87042 86423
rect 87042 86367 87098 86423
rect 87098 86367 87102 86423
rect 87038 86363 87102 86367
rect 87038 86343 87102 86347
rect 87038 86287 87042 86343
rect 87042 86287 87098 86343
rect 87098 86287 87102 86343
rect 87038 86283 87102 86287
rect 87038 86263 87102 86267
rect 87038 86207 87042 86263
rect 87042 86207 87098 86263
rect 87098 86207 87102 86263
rect 87038 86203 87102 86207
rect 88126 86743 88190 86747
rect 88126 86687 88130 86743
rect 88130 86687 88186 86743
rect 88186 86687 88190 86743
rect 88126 86683 88190 86687
rect 88126 86663 88190 86667
rect 88126 86607 88130 86663
rect 88130 86607 88186 86663
rect 88186 86607 88190 86663
rect 88126 86603 88190 86607
rect 88126 86583 88190 86587
rect 88126 86527 88130 86583
rect 88130 86527 88186 86583
rect 88186 86527 88190 86583
rect 88126 86523 88190 86527
rect 88126 86503 88190 86507
rect 88126 86447 88130 86503
rect 88130 86447 88186 86503
rect 88186 86447 88190 86503
rect 88126 86443 88190 86447
rect 88126 86423 88190 86427
rect 88126 86367 88130 86423
rect 88130 86367 88186 86423
rect 88186 86367 88190 86423
rect 88126 86363 88190 86367
rect 88126 86343 88190 86347
rect 88126 86287 88130 86343
rect 88130 86287 88186 86343
rect 88186 86287 88190 86343
rect 88126 86283 88190 86287
rect 88126 86263 88190 86267
rect 88126 86207 88130 86263
rect 88130 86207 88186 86263
rect 88186 86207 88190 86263
rect 88126 86203 88190 86207
rect 48537 78613 48601 78617
rect 48537 78557 48541 78613
rect 48541 78557 48597 78613
rect 48597 78557 48601 78613
rect 48537 78553 48601 78557
rect 50228 78614 50292 78618
rect 50228 78558 50232 78614
rect 50232 78558 50288 78614
rect 50288 78558 50292 78614
rect 50228 78554 50292 78558
rect 51933 78613 51997 78617
rect 51933 78557 51937 78613
rect 51937 78557 51993 78613
rect 51993 78557 51997 78613
rect 51933 78553 51997 78557
rect 53729 78613 53793 78617
rect 53729 78557 53733 78613
rect 53733 78557 53789 78613
rect 53789 78557 53793 78613
rect 53729 78553 53793 78557
rect 55558 78613 55622 78617
rect 55558 78557 55562 78613
rect 55562 78557 55618 78613
rect 55618 78557 55622 78613
rect 55558 78553 55622 78557
rect 47399 78421 47463 78425
rect 47399 78365 47403 78421
rect 47403 78365 47459 78421
rect 47459 78365 47463 78421
rect 47399 78361 47463 78365
rect 47479 78421 47543 78425
rect 47479 78365 47483 78421
rect 47483 78365 47539 78421
rect 47539 78365 47543 78421
rect 47479 78361 47543 78365
rect 47559 78421 47623 78425
rect 47559 78365 47563 78421
rect 47563 78365 47619 78421
rect 47619 78365 47623 78421
rect 47559 78361 47623 78365
rect 49194 78420 49258 78424
rect 49194 78364 49198 78420
rect 49198 78364 49254 78420
rect 49254 78364 49258 78420
rect 49194 78360 49258 78364
rect 49274 78420 49338 78424
rect 49274 78364 49278 78420
rect 49278 78364 49334 78420
rect 49334 78364 49338 78420
rect 49274 78360 49338 78364
rect 49354 78420 49418 78424
rect 49354 78364 49358 78420
rect 49358 78364 49414 78420
rect 49414 78364 49418 78420
rect 49354 78360 49418 78364
rect 50994 78422 51058 78426
rect 50994 78366 50998 78422
rect 50998 78366 51054 78422
rect 51054 78366 51058 78422
rect 50994 78362 51058 78366
rect 51074 78422 51138 78426
rect 51074 78366 51078 78422
rect 51078 78366 51134 78422
rect 51134 78366 51138 78422
rect 51074 78362 51138 78366
rect 51154 78422 51218 78426
rect 51154 78366 51158 78422
rect 51158 78366 51214 78422
rect 51214 78366 51218 78422
rect 51154 78362 51218 78366
rect 52792 78421 52856 78425
rect 52792 78365 52796 78421
rect 52796 78365 52852 78421
rect 52852 78365 52856 78421
rect 52792 78361 52856 78365
rect 52872 78421 52936 78425
rect 52872 78365 52876 78421
rect 52876 78365 52932 78421
rect 52932 78365 52936 78421
rect 52872 78361 52936 78365
rect 52952 78421 53016 78425
rect 52952 78365 52956 78421
rect 52956 78365 53012 78421
rect 53012 78365 53016 78421
rect 52952 78361 53016 78365
rect 54590 78422 54654 78426
rect 54590 78366 54594 78422
rect 54594 78366 54650 78422
rect 54650 78366 54654 78422
rect 54590 78362 54654 78366
rect 54670 78422 54734 78426
rect 54670 78366 54674 78422
rect 54674 78366 54730 78422
rect 54730 78366 54734 78422
rect 54670 78362 54734 78366
rect 54750 78422 54814 78426
rect 54750 78366 54754 78422
rect 54754 78366 54810 78422
rect 54810 78366 54814 78422
rect 54750 78362 54814 78366
rect 56393 78421 56457 78425
rect 56393 78365 56397 78421
rect 56397 78365 56453 78421
rect 56453 78365 56457 78421
rect 56393 78361 56457 78365
rect 56473 78421 56537 78425
rect 56473 78365 56477 78421
rect 56477 78365 56533 78421
rect 56533 78365 56537 78421
rect 56473 78361 56537 78365
rect 56553 78421 56617 78425
rect 56553 78365 56557 78421
rect 56557 78365 56613 78421
rect 56613 78365 56617 78421
rect 56553 78361 56617 78365
rect 57270 78422 57334 78426
rect 57270 78366 57274 78422
rect 57274 78366 57330 78422
rect 57330 78366 57334 78422
rect 57270 78362 57334 78366
rect 49829 78041 49893 78105
rect 55229 78041 55293 78105
rect 49021 77788 49085 77852
rect 54421 77788 54485 77852
rect 46558 77360 46622 77424
rect 55229 77360 55293 77424
rect 45789 77104 45853 77168
rect 54421 77104 54485 77168
rect 57455 84824 57599 84828
rect 57455 77168 57459 84824
rect 57459 77168 57595 84824
rect 57595 77168 57599 84824
rect 57455 77164 57599 77168
rect 44779 76671 44843 76735
rect 49829 76671 49893 76735
rect 43998 76348 44062 76412
rect 49021 76348 49085 76412
rect 48250 75261 48314 75265
rect 48250 75205 48254 75261
rect 48254 75205 48310 75261
rect 48310 75205 48314 75261
rect 48250 75201 48314 75205
rect 48250 75181 48314 75185
rect 48250 75125 48254 75181
rect 48254 75125 48310 75181
rect 48310 75125 48314 75181
rect 48250 75121 48314 75125
rect 49372 75265 49436 75269
rect 49372 75209 49376 75265
rect 49376 75209 49432 75265
rect 49432 75209 49436 75265
rect 49372 75205 49436 75209
rect 48250 75101 48314 75105
rect 48250 75045 48254 75101
rect 48254 75045 48310 75101
rect 48310 75045 48314 75101
rect 48250 75041 48314 75045
rect 51434 75064 53178 75068
rect 51434 74928 51438 75064
rect 51438 74928 53174 75064
rect 53174 74928 53178 75064
rect 51434 74924 53178 74928
rect 53753 75075 54537 75079
rect 53753 74939 53757 75075
rect 53757 74939 54533 75075
rect 54533 74939 54537 75075
rect 53753 74935 54537 74939
rect 55452 75065 56316 75069
rect 55452 74929 55456 75065
rect 55456 74929 56312 75065
rect 56312 74929 56316 75065
rect 55452 74925 56316 74929
rect 48235 74794 48299 74798
rect 48235 74738 48239 74794
rect 48239 74738 48295 74794
rect 48295 74738 48299 74794
rect 48235 74734 48299 74738
rect 48235 74714 48299 74718
rect 48235 74658 48239 74714
rect 48239 74658 48295 74714
rect 48295 74658 48299 74714
rect 48235 74654 48299 74658
rect 48235 74634 48299 74638
rect 38089 74554 38153 74618
rect 48235 74578 48239 74634
rect 48239 74578 48295 74634
rect 48295 74578 48299 74634
rect 48235 74574 48299 74578
rect 48235 74554 48299 74558
rect 48235 74498 48239 74554
rect 48239 74498 48295 74554
rect 48295 74498 48299 74554
rect 48235 74494 48299 74498
rect 48235 74474 48299 74478
rect 48235 74418 48239 74474
rect 48239 74418 48295 74474
rect 48295 74418 48299 74474
rect 48235 74414 48299 74418
rect 48614 74459 48678 74463
rect 48614 74403 48618 74459
rect 48618 74403 48674 74459
rect 48674 74403 48678 74459
rect 48614 74399 48678 74403
rect 48614 74030 48678 74094
rect 30044 73738 30108 73742
rect 30044 73682 30048 73738
rect 30048 73682 30104 73738
rect 30104 73682 30108 73738
rect 30044 73678 30108 73682
rect 30124 73738 30188 73742
rect 30124 73682 30128 73738
rect 30128 73682 30184 73738
rect 30184 73682 30188 73738
rect 30124 73678 30188 73682
rect 30204 73738 30268 73742
rect 30204 73682 30208 73738
rect 30208 73682 30264 73738
rect 30264 73682 30268 73738
rect 30204 73678 30268 73682
rect 30284 73738 30348 73742
rect 30284 73682 30288 73738
rect 30288 73682 30344 73738
rect 30344 73682 30348 73738
rect 30284 73678 30348 73682
rect 49372 73382 49436 73446
rect 31130 73196 31194 73200
rect 31130 73140 31134 73196
rect 31134 73140 31190 73196
rect 31190 73140 31194 73196
rect 31130 73136 31194 73140
rect 31210 73196 31274 73200
rect 31210 73140 31214 73196
rect 31214 73140 31270 73196
rect 31270 73140 31274 73196
rect 31210 73136 31274 73140
rect 31290 73196 31354 73200
rect 31290 73140 31294 73196
rect 31294 73140 31350 73196
rect 31350 73140 31354 73196
rect 31290 73136 31354 73140
rect 31370 73196 31434 73200
rect 31370 73140 31374 73196
rect 31374 73140 31430 73196
rect 31430 73140 31434 73196
rect 31370 73136 31434 73140
rect 51182 74738 51326 74742
rect 51182 71802 51186 74738
rect 51186 71802 51322 74738
rect 51322 71802 51326 74738
rect 51182 71798 51326 71802
rect 57043 71813 57047 74757
rect 57047 71813 57183 74757
rect 57183 71813 57187 74757
rect 67306 84836 67610 84840
rect 67306 71660 67310 84836
rect 67310 71660 67606 84836
rect 67606 71660 67610 84836
rect 67306 71656 67610 71660
rect 74525 84746 74589 84750
rect 74525 84690 74529 84746
rect 74529 84690 74585 84746
rect 74585 84690 74589 84746
rect 74525 84686 74589 84690
rect 74525 84666 74589 84670
rect 74525 84610 74529 84666
rect 74529 84610 74585 84666
rect 74585 84610 74589 84666
rect 74525 84606 74589 84610
rect 74525 84586 74589 84590
rect 74525 84530 74529 84586
rect 74529 84530 74585 84586
rect 74585 84530 74589 84586
rect 74525 84526 74589 84530
rect 74525 84506 74589 84510
rect 74525 84450 74529 84506
rect 74529 84450 74585 84506
rect 74585 84450 74589 84506
rect 74525 84446 74589 84450
rect 74525 84426 74589 84430
rect 74525 84370 74529 84426
rect 74529 84370 74585 84426
rect 74585 84370 74589 84426
rect 74525 84366 74589 84370
rect 74525 84346 74589 84350
rect 74525 84290 74529 84346
rect 74529 84290 74585 84346
rect 74585 84290 74589 84346
rect 74525 84286 74589 84290
rect 74525 84266 74589 84270
rect 74525 84210 74529 84266
rect 74529 84210 74585 84266
rect 74585 84210 74589 84266
rect 74525 84206 74589 84210
rect 75613 84746 75677 84750
rect 75613 84690 75617 84746
rect 75617 84690 75673 84746
rect 75673 84690 75677 84746
rect 75613 84686 75677 84690
rect 75613 84666 75677 84670
rect 75613 84610 75617 84666
rect 75617 84610 75673 84666
rect 75673 84610 75677 84666
rect 75613 84606 75677 84610
rect 75613 84586 75677 84590
rect 75613 84530 75617 84586
rect 75617 84530 75673 84586
rect 75673 84530 75677 84586
rect 75613 84526 75677 84530
rect 75613 84506 75677 84510
rect 75613 84450 75617 84506
rect 75617 84450 75673 84506
rect 75673 84450 75677 84506
rect 75613 84446 75677 84450
rect 75613 84426 75677 84430
rect 75613 84370 75617 84426
rect 75617 84370 75673 84426
rect 75673 84370 75677 84426
rect 75613 84366 75677 84370
rect 75613 84346 75677 84350
rect 75613 84290 75617 84346
rect 75617 84290 75673 84346
rect 75673 84290 75677 84346
rect 75613 84286 75677 84290
rect 75613 84266 75677 84270
rect 75613 84210 75617 84266
rect 75617 84210 75673 84266
rect 75673 84210 75677 84266
rect 75613 84206 75677 84210
rect 76701 84746 76765 84750
rect 76701 84690 76705 84746
rect 76705 84690 76761 84746
rect 76761 84690 76765 84746
rect 76701 84686 76765 84690
rect 76701 84666 76765 84670
rect 76701 84610 76705 84666
rect 76705 84610 76761 84666
rect 76761 84610 76765 84666
rect 76701 84606 76765 84610
rect 76701 84586 76765 84590
rect 76701 84530 76705 84586
rect 76705 84530 76761 84586
rect 76761 84530 76765 84586
rect 76701 84526 76765 84530
rect 76701 84506 76765 84510
rect 76701 84450 76705 84506
rect 76705 84450 76761 84506
rect 76761 84450 76765 84506
rect 76701 84446 76765 84450
rect 76701 84426 76765 84430
rect 76701 84370 76705 84426
rect 76705 84370 76761 84426
rect 76761 84370 76765 84426
rect 76701 84366 76765 84370
rect 76701 84346 76765 84350
rect 76701 84290 76705 84346
rect 76705 84290 76761 84346
rect 76761 84290 76765 84346
rect 76701 84286 76765 84290
rect 76701 84266 76765 84270
rect 76701 84210 76705 84266
rect 76705 84210 76761 84266
rect 76761 84210 76765 84266
rect 76701 84206 76765 84210
rect 77789 84746 77853 84750
rect 77789 84690 77793 84746
rect 77793 84690 77849 84746
rect 77849 84690 77853 84746
rect 77789 84686 77853 84690
rect 77789 84666 77853 84670
rect 77789 84610 77793 84666
rect 77793 84610 77849 84666
rect 77849 84610 77853 84666
rect 77789 84606 77853 84610
rect 77789 84586 77853 84590
rect 77789 84530 77793 84586
rect 77793 84530 77849 84586
rect 77849 84530 77853 84586
rect 77789 84526 77853 84530
rect 77789 84506 77853 84510
rect 77789 84450 77793 84506
rect 77793 84450 77849 84506
rect 77849 84450 77853 84506
rect 77789 84446 77853 84450
rect 77789 84426 77853 84430
rect 77789 84370 77793 84426
rect 77793 84370 77849 84426
rect 77849 84370 77853 84426
rect 77789 84366 77853 84370
rect 77789 84346 77853 84350
rect 77789 84290 77793 84346
rect 77793 84290 77849 84346
rect 77849 84290 77853 84346
rect 77789 84286 77853 84290
rect 77789 84266 77853 84270
rect 77789 84210 77793 84266
rect 77793 84210 77849 84266
rect 77849 84210 77853 84266
rect 77789 84206 77853 84210
rect 78877 84746 78941 84750
rect 78877 84690 78881 84746
rect 78881 84690 78937 84746
rect 78937 84690 78941 84746
rect 78877 84686 78941 84690
rect 78877 84666 78941 84670
rect 78877 84610 78881 84666
rect 78881 84610 78937 84666
rect 78937 84610 78941 84666
rect 78877 84606 78941 84610
rect 78877 84586 78941 84590
rect 78877 84530 78881 84586
rect 78881 84530 78937 84586
rect 78937 84530 78941 84586
rect 78877 84526 78941 84530
rect 78877 84506 78941 84510
rect 78877 84450 78881 84506
rect 78881 84450 78937 84506
rect 78937 84450 78941 84506
rect 78877 84446 78941 84450
rect 78877 84426 78941 84430
rect 78877 84370 78881 84426
rect 78881 84370 78937 84426
rect 78937 84370 78941 84426
rect 78877 84366 78941 84370
rect 78877 84346 78941 84350
rect 78877 84290 78881 84346
rect 78881 84290 78937 84346
rect 78937 84290 78941 84346
rect 78877 84286 78941 84290
rect 78877 84266 78941 84270
rect 78877 84210 78881 84266
rect 78881 84210 78937 84266
rect 78937 84210 78941 84266
rect 78877 84206 78941 84210
rect 79965 84746 80029 84750
rect 79965 84690 79969 84746
rect 79969 84690 80025 84746
rect 80025 84690 80029 84746
rect 79965 84686 80029 84690
rect 79965 84666 80029 84670
rect 79965 84610 79969 84666
rect 79969 84610 80025 84666
rect 80025 84610 80029 84666
rect 79965 84606 80029 84610
rect 79965 84586 80029 84590
rect 79965 84530 79969 84586
rect 79969 84530 80025 84586
rect 80025 84530 80029 84586
rect 79965 84526 80029 84530
rect 79965 84506 80029 84510
rect 79965 84450 79969 84506
rect 79969 84450 80025 84506
rect 80025 84450 80029 84506
rect 79965 84446 80029 84450
rect 79965 84426 80029 84430
rect 79965 84370 79969 84426
rect 79969 84370 80025 84426
rect 80025 84370 80029 84426
rect 79965 84366 80029 84370
rect 79965 84346 80029 84350
rect 79965 84290 79969 84346
rect 79969 84290 80025 84346
rect 80025 84290 80029 84346
rect 79965 84286 80029 84290
rect 79965 84266 80029 84270
rect 79965 84210 79969 84266
rect 79969 84210 80025 84266
rect 80025 84210 80029 84266
rect 79965 84206 80029 84210
rect 81053 84746 81117 84750
rect 81053 84690 81057 84746
rect 81057 84690 81113 84746
rect 81113 84690 81117 84746
rect 81053 84686 81117 84690
rect 81053 84666 81117 84670
rect 81053 84610 81057 84666
rect 81057 84610 81113 84666
rect 81113 84610 81117 84666
rect 81053 84606 81117 84610
rect 81053 84586 81117 84590
rect 81053 84530 81057 84586
rect 81057 84530 81113 84586
rect 81113 84530 81117 84586
rect 81053 84526 81117 84530
rect 81053 84506 81117 84510
rect 81053 84450 81057 84506
rect 81057 84450 81113 84506
rect 81113 84450 81117 84506
rect 81053 84446 81117 84450
rect 81053 84426 81117 84430
rect 81053 84370 81057 84426
rect 81057 84370 81113 84426
rect 81113 84370 81117 84426
rect 81053 84366 81117 84370
rect 81053 84346 81117 84350
rect 81053 84290 81057 84346
rect 81057 84290 81113 84346
rect 81113 84290 81117 84346
rect 81053 84286 81117 84290
rect 81053 84266 81117 84270
rect 81053 84210 81057 84266
rect 81057 84210 81113 84266
rect 81113 84210 81117 84266
rect 81053 84206 81117 84210
rect 82141 84746 82205 84750
rect 82141 84690 82145 84746
rect 82145 84690 82201 84746
rect 82201 84690 82205 84746
rect 82141 84686 82205 84690
rect 82141 84666 82205 84670
rect 82141 84610 82145 84666
rect 82145 84610 82201 84666
rect 82201 84610 82205 84666
rect 82141 84606 82205 84610
rect 82141 84586 82205 84590
rect 82141 84530 82145 84586
rect 82145 84530 82201 84586
rect 82201 84530 82205 84586
rect 82141 84526 82205 84530
rect 82141 84506 82205 84510
rect 82141 84450 82145 84506
rect 82145 84450 82201 84506
rect 82201 84450 82205 84506
rect 82141 84446 82205 84450
rect 82141 84426 82205 84430
rect 82141 84370 82145 84426
rect 82145 84370 82201 84426
rect 82201 84370 82205 84426
rect 82141 84366 82205 84370
rect 82141 84346 82205 84350
rect 82141 84290 82145 84346
rect 82145 84290 82201 84346
rect 82201 84290 82205 84346
rect 82141 84286 82205 84290
rect 82141 84266 82205 84270
rect 82141 84210 82145 84266
rect 82145 84210 82201 84266
rect 82201 84210 82205 84266
rect 82141 84206 82205 84210
rect 83229 84746 83293 84750
rect 83229 84690 83233 84746
rect 83233 84690 83289 84746
rect 83289 84690 83293 84746
rect 83229 84686 83293 84690
rect 83229 84666 83293 84670
rect 83229 84610 83233 84666
rect 83233 84610 83289 84666
rect 83289 84610 83293 84666
rect 83229 84606 83293 84610
rect 83229 84586 83293 84590
rect 83229 84530 83233 84586
rect 83233 84530 83289 84586
rect 83289 84530 83293 84586
rect 83229 84526 83293 84530
rect 83229 84506 83293 84510
rect 83229 84450 83233 84506
rect 83233 84450 83289 84506
rect 83289 84450 83293 84506
rect 83229 84446 83293 84450
rect 83229 84426 83293 84430
rect 83229 84370 83233 84426
rect 83233 84370 83289 84426
rect 83289 84370 83293 84426
rect 83229 84366 83293 84370
rect 83229 84346 83293 84350
rect 83229 84290 83233 84346
rect 83233 84290 83289 84346
rect 83289 84290 83293 84346
rect 83229 84286 83293 84290
rect 83229 84266 83293 84270
rect 83229 84210 83233 84266
rect 83233 84210 83289 84266
rect 83289 84210 83293 84266
rect 83229 84206 83293 84210
rect 84317 84746 84381 84750
rect 84317 84690 84321 84746
rect 84321 84690 84377 84746
rect 84377 84690 84381 84746
rect 84317 84686 84381 84690
rect 84317 84666 84381 84670
rect 84317 84610 84321 84666
rect 84321 84610 84377 84666
rect 84377 84610 84381 84666
rect 84317 84606 84381 84610
rect 84317 84586 84381 84590
rect 84317 84530 84321 84586
rect 84321 84530 84377 84586
rect 84377 84530 84381 84586
rect 84317 84526 84381 84530
rect 84317 84506 84381 84510
rect 84317 84450 84321 84506
rect 84321 84450 84377 84506
rect 84377 84450 84381 84506
rect 84317 84446 84381 84450
rect 84317 84426 84381 84430
rect 84317 84370 84321 84426
rect 84321 84370 84377 84426
rect 84377 84370 84381 84426
rect 84317 84366 84381 84370
rect 84317 84346 84381 84350
rect 84317 84290 84321 84346
rect 84321 84290 84377 84346
rect 84377 84290 84381 84346
rect 84317 84286 84381 84290
rect 84317 84266 84381 84270
rect 84317 84210 84321 84266
rect 84321 84210 84377 84266
rect 84377 84210 84381 84266
rect 84317 84206 84381 84210
rect 85405 84746 85469 84750
rect 85405 84690 85409 84746
rect 85409 84690 85465 84746
rect 85465 84690 85469 84746
rect 85405 84686 85469 84690
rect 85405 84666 85469 84670
rect 85405 84610 85409 84666
rect 85409 84610 85465 84666
rect 85465 84610 85469 84666
rect 85405 84606 85469 84610
rect 85405 84586 85469 84590
rect 85405 84530 85409 84586
rect 85409 84530 85465 84586
rect 85465 84530 85469 84586
rect 85405 84526 85469 84530
rect 85405 84506 85469 84510
rect 85405 84450 85409 84506
rect 85409 84450 85465 84506
rect 85465 84450 85469 84506
rect 85405 84446 85469 84450
rect 85405 84426 85469 84430
rect 85405 84370 85409 84426
rect 85409 84370 85465 84426
rect 85465 84370 85469 84426
rect 85405 84366 85469 84370
rect 85405 84346 85469 84350
rect 85405 84290 85409 84346
rect 85409 84290 85465 84346
rect 85465 84290 85469 84346
rect 85405 84286 85469 84290
rect 85405 84266 85469 84270
rect 85405 84210 85409 84266
rect 85409 84210 85465 84266
rect 85465 84210 85469 84266
rect 85405 84206 85469 84210
rect 86493 84746 86557 84750
rect 86493 84690 86497 84746
rect 86497 84690 86553 84746
rect 86553 84690 86557 84746
rect 86493 84686 86557 84690
rect 86493 84666 86557 84670
rect 86493 84610 86497 84666
rect 86497 84610 86553 84666
rect 86553 84610 86557 84666
rect 86493 84606 86557 84610
rect 86493 84586 86557 84590
rect 86493 84530 86497 84586
rect 86497 84530 86553 84586
rect 86553 84530 86557 84586
rect 86493 84526 86557 84530
rect 86493 84506 86557 84510
rect 86493 84450 86497 84506
rect 86497 84450 86553 84506
rect 86553 84450 86557 84506
rect 86493 84446 86557 84450
rect 86493 84426 86557 84430
rect 86493 84370 86497 84426
rect 86497 84370 86553 84426
rect 86553 84370 86557 84426
rect 86493 84366 86557 84370
rect 86493 84346 86557 84350
rect 86493 84290 86497 84346
rect 86497 84290 86553 84346
rect 86553 84290 86557 84346
rect 86493 84286 86557 84290
rect 86493 84266 86557 84270
rect 86493 84210 86497 84266
rect 86497 84210 86553 84266
rect 86553 84210 86557 84266
rect 86493 84206 86557 84210
rect 87581 84746 87645 84750
rect 87581 84690 87585 84746
rect 87585 84690 87641 84746
rect 87641 84690 87645 84746
rect 87581 84686 87645 84690
rect 87581 84666 87645 84670
rect 87581 84610 87585 84666
rect 87585 84610 87641 84666
rect 87641 84610 87645 84666
rect 87581 84606 87645 84610
rect 87581 84586 87645 84590
rect 87581 84530 87585 84586
rect 87585 84530 87641 84586
rect 87641 84530 87645 84586
rect 87581 84526 87645 84530
rect 87581 84506 87645 84510
rect 87581 84450 87585 84506
rect 87585 84450 87641 84506
rect 87641 84450 87645 84506
rect 87581 84446 87645 84450
rect 87581 84426 87645 84430
rect 87581 84370 87585 84426
rect 87585 84370 87641 84426
rect 87641 84370 87645 84426
rect 87581 84366 87645 84370
rect 87581 84346 87645 84350
rect 87581 84290 87585 84346
rect 87585 84290 87641 84346
rect 87641 84290 87645 84346
rect 87581 84286 87645 84290
rect 87581 84266 87645 84270
rect 87581 84210 87585 84266
rect 87585 84210 87641 84266
rect 87641 84210 87645 84266
rect 87581 84206 87645 84210
rect 88669 84746 88733 84750
rect 88669 84690 88673 84746
rect 88673 84690 88729 84746
rect 88729 84690 88733 84746
rect 88669 84686 88733 84690
rect 88669 84666 88733 84670
rect 88669 84610 88673 84666
rect 88673 84610 88729 84666
rect 88729 84610 88733 84666
rect 88669 84606 88733 84610
rect 88669 84586 88733 84590
rect 88669 84530 88673 84586
rect 88673 84530 88729 84586
rect 88729 84530 88733 84586
rect 88669 84526 88733 84530
rect 88669 84506 88733 84510
rect 88669 84450 88673 84506
rect 88673 84450 88729 84506
rect 88729 84450 88733 84506
rect 88669 84446 88733 84450
rect 88669 84426 88733 84430
rect 88669 84370 88673 84426
rect 88673 84370 88729 84426
rect 88729 84370 88733 84426
rect 88669 84366 88733 84370
rect 88669 84346 88733 84350
rect 88669 84290 88673 84346
rect 88673 84290 88729 84346
rect 88729 84290 88733 84346
rect 88669 84286 88733 84290
rect 88669 84266 88733 84270
rect 88669 84210 88673 84266
rect 88673 84210 88729 84266
rect 88729 84210 88733 84266
rect 88669 84206 88733 84210
rect 75070 82743 75134 82747
rect 75070 82687 75074 82743
rect 75074 82687 75130 82743
rect 75130 82687 75134 82743
rect 75070 82683 75134 82687
rect 75070 82663 75134 82667
rect 75070 82607 75074 82663
rect 75074 82607 75130 82663
rect 75130 82607 75134 82663
rect 75070 82603 75134 82607
rect 75070 82583 75134 82587
rect 75070 82527 75074 82583
rect 75074 82527 75130 82583
rect 75130 82527 75134 82583
rect 75070 82523 75134 82527
rect 75070 82503 75134 82507
rect 75070 82447 75074 82503
rect 75074 82447 75130 82503
rect 75130 82447 75134 82503
rect 75070 82443 75134 82447
rect 75070 82423 75134 82427
rect 75070 82367 75074 82423
rect 75074 82367 75130 82423
rect 75130 82367 75134 82423
rect 75070 82363 75134 82367
rect 75070 82343 75134 82347
rect 75070 82287 75074 82343
rect 75074 82287 75130 82343
rect 75130 82287 75134 82343
rect 75070 82283 75134 82287
rect 75070 82263 75134 82267
rect 75070 82207 75074 82263
rect 75074 82207 75130 82263
rect 75130 82207 75134 82263
rect 75070 82203 75134 82207
rect 76158 82743 76222 82747
rect 76158 82687 76162 82743
rect 76162 82687 76218 82743
rect 76218 82687 76222 82743
rect 76158 82683 76222 82687
rect 76158 82663 76222 82667
rect 76158 82607 76162 82663
rect 76162 82607 76218 82663
rect 76218 82607 76222 82663
rect 76158 82603 76222 82607
rect 76158 82583 76222 82587
rect 76158 82527 76162 82583
rect 76162 82527 76218 82583
rect 76218 82527 76222 82583
rect 76158 82523 76222 82527
rect 76158 82503 76222 82507
rect 76158 82447 76162 82503
rect 76162 82447 76218 82503
rect 76218 82447 76222 82503
rect 76158 82443 76222 82447
rect 76158 82423 76222 82427
rect 76158 82367 76162 82423
rect 76162 82367 76218 82423
rect 76218 82367 76222 82423
rect 76158 82363 76222 82367
rect 76158 82343 76222 82347
rect 76158 82287 76162 82343
rect 76162 82287 76218 82343
rect 76218 82287 76222 82343
rect 76158 82283 76222 82287
rect 76158 82263 76222 82267
rect 76158 82207 76162 82263
rect 76162 82207 76218 82263
rect 76218 82207 76222 82263
rect 76158 82203 76222 82207
rect 77246 82743 77310 82747
rect 77246 82687 77250 82743
rect 77250 82687 77306 82743
rect 77306 82687 77310 82743
rect 77246 82683 77310 82687
rect 77246 82663 77310 82667
rect 77246 82607 77250 82663
rect 77250 82607 77306 82663
rect 77306 82607 77310 82663
rect 77246 82603 77310 82607
rect 77246 82583 77310 82587
rect 77246 82527 77250 82583
rect 77250 82527 77306 82583
rect 77306 82527 77310 82583
rect 77246 82523 77310 82527
rect 77246 82503 77310 82507
rect 77246 82447 77250 82503
rect 77250 82447 77306 82503
rect 77306 82447 77310 82503
rect 77246 82443 77310 82447
rect 77246 82423 77310 82427
rect 77246 82367 77250 82423
rect 77250 82367 77306 82423
rect 77306 82367 77310 82423
rect 77246 82363 77310 82367
rect 77246 82343 77310 82347
rect 77246 82287 77250 82343
rect 77250 82287 77306 82343
rect 77306 82287 77310 82343
rect 77246 82283 77310 82287
rect 77246 82263 77310 82267
rect 77246 82207 77250 82263
rect 77250 82207 77306 82263
rect 77306 82207 77310 82263
rect 77246 82203 77310 82207
rect 78334 82743 78398 82747
rect 78334 82687 78338 82743
rect 78338 82687 78394 82743
rect 78394 82687 78398 82743
rect 78334 82683 78398 82687
rect 78334 82663 78398 82667
rect 78334 82607 78338 82663
rect 78338 82607 78394 82663
rect 78394 82607 78398 82663
rect 78334 82603 78398 82607
rect 78334 82583 78398 82587
rect 78334 82527 78338 82583
rect 78338 82527 78394 82583
rect 78394 82527 78398 82583
rect 78334 82523 78398 82527
rect 78334 82503 78398 82507
rect 78334 82447 78338 82503
rect 78338 82447 78394 82503
rect 78394 82447 78398 82503
rect 78334 82443 78398 82447
rect 78334 82423 78398 82427
rect 78334 82367 78338 82423
rect 78338 82367 78394 82423
rect 78394 82367 78398 82423
rect 78334 82363 78398 82367
rect 78334 82343 78398 82347
rect 78334 82287 78338 82343
rect 78338 82287 78394 82343
rect 78394 82287 78398 82343
rect 78334 82283 78398 82287
rect 78334 82263 78398 82267
rect 78334 82207 78338 82263
rect 78338 82207 78394 82263
rect 78394 82207 78398 82263
rect 78334 82203 78398 82207
rect 79422 82743 79486 82747
rect 79422 82687 79426 82743
rect 79426 82687 79482 82743
rect 79482 82687 79486 82743
rect 79422 82683 79486 82687
rect 79422 82663 79486 82667
rect 79422 82607 79426 82663
rect 79426 82607 79482 82663
rect 79482 82607 79486 82663
rect 79422 82603 79486 82607
rect 79422 82583 79486 82587
rect 79422 82527 79426 82583
rect 79426 82527 79482 82583
rect 79482 82527 79486 82583
rect 79422 82523 79486 82527
rect 79422 82503 79486 82507
rect 79422 82447 79426 82503
rect 79426 82447 79482 82503
rect 79482 82447 79486 82503
rect 79422 82443 79486 82447
rect 79422 82423 79486 82427
rect 79422 82367 79426 82423
rect 79426 82367 79482 82423
rect 79482 82367 79486 82423
rect 79422 82363 79486 82367
rect 79422 82343 79486 82347
rect 79422 82287 79426 82343
rect 79426 82287 79482 82343
rect 79482 82287 79486 82343
rect 79422 82283 79486 82287
rect 79422 82263 79486 82267
rect 79422 82207 79426 82263
rect 79426 82207 79482 82263
rect 79482 82207 79486 82263
rect 79422 82203 79486 82207
rect 80510 82743 80574 82747
rect 80510 82687 80514 82743
rect 80514 82687 80570 82743
rect 80570 82687 80574 82743
rect 80510 82683 80574 82687
rect 80510 82663 80574 82667
rect 80510 82607 80514 82663
rect 80514 82607 80570 82663
rect 80570 82607 80574 82663
rect 80510 82603 80574 82607
rect 80510 82583 80574 82587
rect 80510 82527 80514 82583
rect 80514 82527 80570 82583
rect 80570 82527 80574 82583
rect 80510 82523 80574 82527
rect 80510 82503 80574 82507
rect 80510 82447 80514 82503
rect 80514 82447 80570 82503
rect 80570 82447 80574 82503
rect 80510 82443 80574 82447
rect 80510 82423 80574 82427
rect 80510 82367 80514 82423
rect 80514 82367 80570 82423
rect 80570 82367 80574 82423
rect 80510 82363 80574 82367
rect 80510 82343 80574 82347
rect 80510 82287 80514 82343
rect 80514 82287 80570 82343
rect 80570 82287 80574 82343
rect 80510 82283 80574 82287
rect 80510 82263 80574 82267
rect 80510 82207 80514 82263
rect 80514 82207 80570 82263
rect 80570 82207 80574 82263
rect 80510 82203 80574 82207
rect 81598 82743 81662 82747
rect 81598 82687 81602 82743
rect 81602 82687 81658 82743
rect 81658 82687 81662 82743
rect 81598 82683 81662 82687
rect 81598 82663 81662 82667
rect 81598 82607 81602 82663
rect 81602 82607 81658 82663
rect 81658 82607 81662 82663
rect 81598 82603 81662 82607
rect 81598 82583 81662 82587
rect 81598 82527 81602 82583
rect 81602 82527 81658 82583
rect 81658 82527 81662 82583
rect 81598 82523 81662 82527
rect 81598 82503 81662 82507
rect 81598 82447 81602 82503
rect 81602 82447 81658 82503
rect 81658 82447 81662 82503
rect 81598 82443 81662 82447
rect 81598 82423 81662 82427
rect 81598 82367 81602 82423
rect 81602 82367 81658 82423
rect 81658 82367 81662 82423
rect 81598 82363 81662 82367
rect 81598 82343 81662 82347
rect 81598 82287 81602 82343
rect 81602 82287 81658 82343
rect 81658 82287 81662 82343
rect 81598 82283 81662 82287
rect 81598 82263 81662 82267
rect 81598 82207 81602 82263
rect 81602 82207 81658 82263
rect 81658 82207 81662 82263
rect 81598 82203 81662 82207
rect 82686 82743 82750 82747
rect 82686 82687 82690 82743
rect 82690 82687 82746 82743
rect 82746 82687 82750 82743
rect 82686 82683 82750 82687
rect 82686 82663 82750 82667
rect 82686 82607 82690 82663
rect 82690 82607 82746 82663
rect 82746 82607 82750 82663
rect 82686 82603 82750 82607
rect 82686 82583 82750 82587
rect 82686 82527 82690 82583
rect 82690 82527 82746 82583
rect 82746 82527 82750 82583
rect 82686 82523 82750 82527
rect 82686 82503 82750 82507
rect 82686 82447 82690 82503
rect 82690 82447 82746 82503
rect 82746 82447 82750 82503
rect 82686 82443 82750 82447
rect 82686 82423 82750 82427
rect 82686 82367 82690 82423
rect 82690 82367 82746 82423
rect 82746 82367 82750 82423
rect 82686 82363 82750 82367
rect 82686 82343 82750 82347
rect 82686 82287 82690 82343
rect 82690 82287 82746 82343
rect 82746 82287 82750 82343
rect 82686 82283 82750 82287
rect 82686 82263 82750 82267
rect 82686 82207 82690 82263
rect 82690 82207 82746 82263
rect 82746 82207 82750 82263
rect 82686 82203 82750 82207
rect 83774 82743 83838 82747
rect 83774 82687 83778 82743
rect 83778 82687 83834 82743
rect 83834 82687 83838 82743
rect 83774 82683 83838 82687
rect 83774 82663 83838 82667
rect 83774 82607 83778 82663
rect 83778 82607 83834 82663
rect 83834 82607 83838 82663
rect 83774 82603 83838 82607
rect 83774 82583 83838 82587
rect 83774 82527 83778 82583
rect 83778 82527 83834 82583
rect 83834 82527 83838 82583
rect 83774 82523 83838 82527
rect 83774 82503 83838 82507
rect 83774 82447 83778 82503
rect 83778 82447 83834 82503
rect 83834 82447 83838 82503
rect 83774 82443 83838 82447
rect 83774 82423 83838 82427
rect 83774 82367 83778 82423
rect 83778 82367 83834 82423
rect 83834 82367 83838 82423
rect 83774 82363 83838 82367
rect 83774 82343 83838 82347
rect 83774 82287 83778 82343
rect 83778 82287 83834 82343
rect 83834 82287 83838 82343
rect 83774 82283 83838 82287
rect 83774 82263 83838 82267
rect 83774 82207 83778 82263
rect 83778 82207 83834 82263
rect 83834 82207 83838 82263
rect 83774 82203 83838 82207
rect 84862 82743 84926 82747
rect 84862 82687 84866 82743
rect 84866 82687 84922 82743
rect 84922 82687 84926 82743
rect 84862 82683 84926 82687
rect 84862 82663 84926 82667
rect 84862 82607 84866 82663
rect 84866 82607 84922 82663
rect 84922 82607 84926 82663
rect 84862 82603 84926 82607
rect 84862 82583 84926 82587
rect 84862 82527 84866 82583
rect 84866 82527 84922 82583
rect 84922 82527 84926 82583
rect 84862 82523 84926 82527
rect 84862 82503 84926 82507
rect 84862 82447 84866 82503
rect 84866 82447 84922 82503
rect 84922 82447 84926 82503
rect 84862 82443 84926 82447
rect 84862 82423 84926 82427
rect 84862 82367 84866 82423
rect 84866 82367 84922 82423
rect 84922 82367 84926 82423
rect 84862 82363 84926 82367
rect 84862 82343 84926 82347
rect 84862 82287 84866 82343
rect 84866 82287 84922 82343
rect 84922 82287 84926 82343
rect 84862 82283 84926 82287
rect 84862 82263 84926 82267
rect 84862 82207 84866 82263
rect 84866 82207 84922 82263
rect 84922 82207 84926 82263
rect 84862 82203 84926 82207
rect 85950 82743 86014 82747
rect 85950 82687 85954 82743
rect 85954 82687 86010 82743
rect 86010 82687 86014 82743
rect 85950 82683 86014 82687
rect 85950 82663 86014 82667
rect 85950 82607 85954 82663
rect 85954 82607 86010 82663
rect 86010 82607 86014 82663
rect 85950 82603 86014 82607
rect 85950 82583 86014 82587
rect 85950 82527 85954 82583
rect 85954 82527 86010 82583
rect 86010 82527 86014 82583
rect 85950 82523 86014 82527
rect 85950 82503 86014 82507
rect 85950 82447 85954 82503
rect 85954 82447 86010 82503
rect 86010 82447 86014 82503
rect 85950 82443 86014 82447
rect 85950 82423 86014 82427
rect 85950 82367 85954 82423
rect 85954 82367 86010 82423
rect 86010 82367 86014 82423
rect 85950 82363 86014 82367
rect 85950 82343 86014 82347
rect 85950 82287 85954 82343
rect 85954 82287 86010 82343
rect 86010 82287 86014 82343
rect 85950 82283 86014 82287
rect 85950 82263 86014 82267
rect 85950 82207 85954 82263
rect 85954 82207 86010 82263
rect 86010 82207 86014 82263
rect 85950 82203 86014 82207
rect 87038 82743 87102 82747
rect 87038 82687 87042 82743
rect 87042 82687 87098 82743
rect 87098 82687 87102 82743
rect 87038 82683 87102 82687
rect 87038 82663 87102 82667
rect 87038 82607 87042 82663
rect 87042 82607 87098 82663
rect 87098 82607 87102 82663
rect 87038 82603 87102 82607
rect 87038 82583 87102 82587
rect 87038 82527 87042 82583
rect 87042 82527 87098 82583
rect 87098 82527 87102 82583
rect 87038 82523 87102 82527
rect 87038 82503 87102 82507
rect 87038 82447 87042 82503
rect 87042 82447 87098 82503
rect 87098 82447 87102 82503
rect 87038 82443 87102 82447
rect 87038 82423 87102 82427
rect 87038 82367 87042 82423
rect 87042 82367 87098 82423
rect 87098 82367 87102 82423
rect 87038 82363 87102 82367
rect 87038 82343 87102 82347
rect 87038 82287 87042 82343
rect 87042 82287 87098 82343
rect 87098 82287 87102 82343
rect 87038 82283 87102 82287
rect 87038 82263 87102 82267
rect 87038 82207 87042 82263
rect 87042 82207 87098 82263
rect 87098 82207 87102 82263
rect 87038 82203 87102 82207
rect 88126 82743 88190 82747
rect 88126 82687 88130 82743
rect 88130 82687 88186 82743
rect 88186 82687 88190 82743
rect 88126 82683 88190 82687
rect 88126 82663 88190 82667
rect 88126 82607 88130 82663
rect 88130 82607 88186 82663
rect 88186 82607 88190 82663
rect 88126 82603 88190 82607
rect 88126 82583 88190 82587
rect 88126 82527 88130 82583
rect 88130 82527 88186 82583
rect 88186 82527 88190 82583
rect 88126 82523 88190 82527
rect 88126 82503 88190 82507
rect 88126 82447 88130 82503
rect 88130 82447 88186 82503
rect 88186 82447 88190 82503
rect 88126 82443 88190 82447
rect 88126 82423 88190 82427
rect 88126 82367 88130 82423
rect 88130 82367 88186 82423
rect 88186 82367 88190 82423
rect 88126 82363 88190 82367
rect 88126 82343 88190 82347
rect 88126 82287 88130 82343
rect 88130 82287 88186 82343
rect 88186 82287 88190 82343
rect 88126 82283 88190 82287
rect 88126 82263 88190 82267
rect 88126 82207 88130 82263
rect 88130 82207 88186 82263
rect 88186 82207 88190 82263
rect 88126 82203 88190 82207
rect 74525 80746 74589 80750
rect 74525 80690 74529 80746
rect 74529 80690 74585 80746
rect 74585 80690 74589 80746
rect 74525 80686 74589 80690
rect 74525 80666 74589 80670
rect 74525 80610 74529 80666
rect 74529 80610 74585 80666
rect 74585 80610 74589 80666
rect 74525 80606 74589 80610
rect 74525 80586 74589 80590
rect 74525 80530 74529 80586
rect 74529 80530 74585 80586
rect 74585 80530 74589 80586
rect 74525 80526 74589 80530
rect 74525 80506 74589 80510
rect 74525 80450 74529 80506
rect 74529 80450 74585 80506
rect 74585 80450 74589 80506
rect 74525 80446 74589 80450
rect 74525 80426 74589 80430
rect 74525 80370 74529 80426
rect 74529 80370 74585 80426
rect 74585 80370 74589 80426
rect 74525 80366 74589 80370
rect 74525 80346 74589 80350
rect 74525 80290 74529 80346
rect 74529 80290 74585 80346
rect 74585 80290 74589 80346
rect 74525 80286 74589 80290
rect 74525 80266 74589 80270
rect 74525 80210 74529 80266
rect 74529 80210 74585 80266
rect 74585 80210 74589 80266
rect 74525 80206 74589 80210
rect 75613 80746 75677 80750
rect 75613 80690 75617 80746
rect 75617 80690 75673 80746
rect 75673 80690 75677 80746
rect 75613 80686 75677 80690
rect 75613 80666 75677 80670
rect 75613 80610 75617 80666
rect 75617 80610 75673 80666
rect 75673 80610 75677 80666
rect 75613 80606 75677 80610
rect 75613 80586 75677 80590
rect 75613 80530 75617 80586
rect 75617 80530 75673 80586
rect 75673 80530 75677 80586
rect 75613 80526 75677 80530
rect 75613 80506 75677 80510
rect 75613 80450 75617 80506
rect 75617 80450 75673 80506
rect 75673 80450 75677 80506
rect 75613 80446 75677 80450
rect 75613 80426 75677 80430
rect 75613 80370 75617 80426
rect 75617 80370 75673 80426
rect 75673 80370 75677 80426
rect 75613 80366 75677 80370
rect 75613 80346 75677 80350
rect 75613 80290 75617 80346
rect 75617 80290 75673 80346
rect 75673 80290 75677 80346
rect 75613 80286 75677 80290
rect 75613 80266 75677 80270
rect 75613 80210 75617 80266
rect 75617 80210 75673 80266
rect 75673 80210 75677 80266
rect 75613 80206 75677 80210
rect 76701 80746 76765 80750
rect 76701 80690 76705 80746
rect 76705 80690 76761 80746
rect 76761 80690 76765 80746
rect 76701 80686 76765 80690
rect 76701 80666 76765 80670
rect 76701 80610 76705 80666
rect 76705 80610 76761 80666
rect 76761 80610 76765 80666
rect 76701 80606 76765 80610
rect 76701 80586 76765 80590
rect 76701 80530 76705 80586
rect 76705 80530 76761 80586
rect 76761 80530 76765 80586
rect 76701 80526 76765 80530
rect 76701 80506 76765 80510
rect 76701 80450 76705 80506
rect 76705 80450 76761 80506
rect 76761 80450 76765 80506
rect 76701 80446 76765 80450
rect 76701 80426 76765 80430
rect 76701 80370 76705 80426
rect 76705 80370 76761 80426
rect 76761 80370 76765 80426
rect 76701 80366 76765 80370
rect 76701 80346 76765 80350
rect 76701 80290 76705 80346
rect 76705 80290 76761 80346
rect 76761 80290 76765 80346
rect 76701 80286 76765 80290
rect 76701 80266 76765 80270
rect 76701 80210 76705 80266
rect 76705 80210 76761 80266
rect 76761 80210 76765 80266
rect 76701 80206 76765 80210
rect 77789 80746 77853 80750
rect 77789 80690 77793 80746
rect 77793 80690 77849 80746
rect 77849 80690 77853 80746
rect 77789 80686 77853 80690
rect 77789 80666 77853 80670
rect 77789 80610 77793 80666
rect 77793 80610 77849 80666
rect 77849 80610 77853 80666
rect 77789 80606 77853 80610
rect 77789 80586 77853 80590
rect 77789 80530 77793 80586
rect 77793 80530 77849 80586
rect 77849 80530 77853 80586
rect 77789 80526 77853 80530
rect 77789 80506 77853 80510
rect 77789 80450 77793 80506
rect 77793 80450 77849 80506
rect 77849 80450 77853 80506
rect 77789 80446 77853 80450
rect 77789 80426 77853 80430
rect 77789 80370 77793 80426
rect 77793 80370 77849 80426
rect 77849 80370 77853 80426
rect 77789 80366 77853 80370
rect 77789 80346 77853 80350
rect 77789 80290 77793 80346
rect 77793 80290 77849 80346
rect 77849 80290 77853 80346
rect 77789 80286 77853 80290
rect 77789 80266 77853 80270
rect 77789 80210 77793 80266
rect 77793 80210 77849 80266
rect 77849 80210 77853 80266
rect 77789 80206 77853 80210
rect 78877 80746 78941 80750
rect 78877 80690 78881 80746
rect 78881 80690 78937 80746
rect 78937 80690 78941 80746
rect 78877 80686 78941 80690
rect 78877 80666 78941 80670
rect 78877 80610 78881 80666
rect 78881 80610 78937 80666
rect 78937 80610 78941 80666
rect 78877 80606 78941 80610
rect 78877 80586 78941 80590
rect 78877 80530 78881 80586
rect 78881 80530 78937 80586
rect 78937 80530 78941 80586
rect 78877 80526 78941 80530
rect 78877 80506 78941 80510
rect 78877 80450 78881 80506
rect 78881 80450 78937 80506
rect 78937 80450 78941 80506
rect 78877 80446 78941 80450
rect 78877 80426 78941 80430
rect 78877 80370 78881 80426
rect 78881 80370 78937 80426
rect 78937 80370 78941 80426
rect 78877 80366 78941 80370
rect 78877 80346 78941 80350
rect 78877 80290 78881 80346
rect 78881 80290 78937 80346
rect 78937 80290 78941 80346
rect 78877 80286 78941 80290
rect 78877 80266 78941 80270
rect 78877 80210 78881 80266
rect 78881 80210 78937 80266
rect 78937 80210 78941 80266
rect 78877 80206 78941 80210
rect 79965 80746 80029 80750
rect 79965 80690 79969 80746
rect 79969 80690 80025 80746
rect 80025 80690 80029 80746
rect 79965 80686 80029 80690
rect 79965 80666 80029 80670
rect 79965 80610 79969 80666
rect 79969 80610 80025 80666
rect 80025 80610 80029 80666
rect 79965 80606 80029 80610
rect 79965 80586 80029 80590
rect 79965 80530 79969 80586
rect 79969 80530 80025 80586
rect 80025 80530 80029 80586
rect 79965 80526 80029 80530
rect 79965 80506 80029 80510
rect 79965 80450 79969 80506
rect 79969 80450 80025 80506
rect 80025 80450 80029 80506
rect 79965 80446 80029 80450
rect 79965 80426 80029 80430
rect 79965 80370 79969 80426
rect 79969 80370 80025 80426
rect 80025 80370 80029 80426
rect 79965 80366 80029 80370
rect 79965 80346 80029 80350
rect 79965 80290 79969 80346
rect 79969 80290 80025 80346
rect 80025 80290 80029 80346
rect 79965 80286 80029 80290
rect 79965 80266 80029 80270
rect 79965 80210 79969 80266
rect 79969 80210 80025 80266
rect 80025 80210 80029 80266
rect 79965 80206 80029 80210
rect 81053 80746 81117 80750
rect 81053 80690 81057 80746
rect 81057 80690 81113 80746
rect 81113 80690 81117 80746
rect 81053 80686 81117 80690
rect 81053 80666 81117 80670
rect 81053 80610 81057 80666
rect 81057 80610 81113 80666
rect 81113 80610 81117 80666
rect 81053 80606 81117 80610
rect 81053 80586 81117 80590
rect 81053 80530 81057 80586
rect 81057 80530 81113 80586
rect 81113 80530 81117 80586
rect 81053 80526 81117 80530
rect 81053 80506 81117 80510
rect 81053 80450 81057 80506
rect 81057 80450 81113 80506
rect 81113 80450 81117 80506
rect 81053 80446 81117 80450
rect 81053 80426 81117 80430
rect 81053 80370 81057 80426
rect 81057 80370 81113 80426
rect 81113 80370 81117 80426
rect 81053 80366 81117 80370
rect 81053 80346 81117 80350
rect 81053 80290 81057 80346
rect 81057 80290 81113 80346
rect 81113 80290 81117 80346
rect 81053 80286 81117 80290
rect 81053 80266 81117 80270
rect 81053 80210 81057 80266
rect 81057 80210 81113 80266
rect 81113 80210 81117 80266
rect 81053 80206 81117 80210
rect 82141 80746 82205 80750
rect 82141 80690 82145 80746
rect 82145 80690 82201 80746
rect 82201 80690 82205 80746
rect 82141 80686 82205 80690
rect 82141 80666 82205 80670
rect 82141 80610 82145 80666
rect 82145 80610 82201 80666
rect 82201 80610 82205 80666
rect 82141 80606 82205 80610
rect 82141 80586 82205 80590
rect 82141 80530 82145 80586
rect 82145 80530 82201 80586
rect 82201 80530 82205 80586
rect 82141 80526 82205 80530
rect 82141 80506 82205 80510
rect 82141 80450 82145 80506
rect 82145 80450 82201 80506
rect 82201 80450 82205 80506
rect 82141 80446 82205 80450
rect 82141 80426 82205 80430
rect 82141 80370 82145 80426
rect 82145 80370 82201 80426
rect 82201 80370 82205 80426
rect 82141 80366 82205 80370
rect 82141 80346 82205 80350
rect 82141 80290 82145 80346
rect 82145 80290 82201 80346
rect 82201 80290 82205 80346
rect 82141 80286 82205 80290
rect 82141 80266 82205 80270
rect 82141 80210 82145 80266
rect 82145 80210 82201 80266
rect 82201 80210 82205 80266
rect 82141 80206 82205 80210
rect 83229 80746 83293 80750
rect 83229 80690 83233 80746
rect 83233 80690 83289 80746
rect 83289 80690 83293 80746
rect 83229 80686 83293 80690
rect 83229 80666 83293 80670
rect 83229 80610 83233 80666
rect 83233 80610 83289 80666
rect 83289 80610 83293 80666
rect 83229 80606 83293 80610
rect 83229 80586 83293 80590
rect 83229 80530 83233 80586
rect 83233 80530 83289 80586
rect 83289 80530 83293 80586
rect 83229 80526 83293 80530
rect 83229 80506 83293 80510
rect 83229 80450 83233 80506
rect 83233 80450 83289 80506
rect 83289 80450 83293 80506
rect 83229 80446 83293 80450
rect 83229 80426 83293 80430
rect 83229 80370 83233 80426
rect 83233 80370 83289 80426
rect 83289 80370 83293 80426
rect 83229 80366 83293 80370
rect 83229 80346 83293 80350
rect 83229 80290 83233 80346
rect 83233 80290 83289 80346
rect 83289 80290 83293 80346
rect 83229 80286 83293 80290
rect 83229 80266 83293 80270
rect 83229 80210 83233 80266
rect 83233 80210 83289 80266
rect 83289 80210 83293 80266
rect 83229 80206 83293 80210
rect 84317 80746 84381 80750
rect 84317 80690 84321 80746
rect 84321 80690 84377 80746
rect 84377 80690 84381 80746
rect 84317 80686 84381 80690
rect 84317 80666 84381 80670
rect 84317 80610 84321 80666
rect 84321 80610 84377 80666
rect 84377 80610 84381 80666
rect 84317 80606 84381 80610
rect 84317 80586 84381 80590
rect 84317 80530 84321 80586
rect 84321 80530 84377 80586
rect 84377 80530 84381 80586
rect 84317 80526 84381 80530
rect 84317 80506 84381 80510
rect 84317 80450 84321 80506
rect 84321 80450 84377 80506
rect 84377 80450 84381 80506
rect 84317 80446 84381 80450
rect 84317 80426 84381 80430
rect 84317 80370 84321 80426
rect 84321 80370 84377 80426
rect 84377 80370 84381 80426
rect 84317 80366 84381 80370
rect 84317 80346 84381 80350
rect 84317 80290 84321 80346
rect 84321 80290 84377 80346
rect 84377 80290 84381 80346
rect 84317 80286 84381 80290
rect 84317 80266 84381 80270
rect 84317 80210 84321 80266
rect 84321 80210 84377 80266
rect 84377 80210 84381 80266
rect 84317 80206 84381 80210
rect 85405 80746 85469 80750
rect 85405 80690 85409 80746
rect 85409 80690 85465 80746
rect 85465 80690 85469 80746
rect 85405 80686 85469 80690
rect 85405 80666 85469 80670
rect 85405 80610 85409 80666
rect 85409 80610 85465 80666
rect 85465 80610 85469 80666
rect 85405 80606 85469 80610
rect 85405 80586 85469 80590
rect 85405 80530 85409 80586
rect 85409 80530 85465 80586
rect 85465 80530 85469 80586
rect 85405 80526 85469 80530
rect 85405 80506 85469 80510
rect 85405 80450 85409 80506
rect 85409 80450 85465 80506
rect 85465 80450 85469 80506
rect 85405 80446 85469 80450
rect 85405 80426 85469 80430
rect 85405 80370 85409 80426
rect 85409 80370 85465 80426
rect 85465 80370 85469 80426
rect 85405 80366 85469 80370
rect 85405 80346 85469 80350
rect 85405 80290 85409 80346
rect 85409 80290 85465 80346
rect 85465 80290 85469 80346
rect 85405 80286 85469 80290
rect 85405 80266 85469 80270
rect 85405 80210 85409 80266
rect 85409 80210 85465 80266
rect 85465 80210 85469 80266
rect 85405 80206 85469 80210
rect 86493 80746 86557 80750
rect 86493 80690 86497 80746
rect 86497 80690 86553 80746
rect 86553 80690 86557 80746
rect 86493 80686 86557 80690
rect 86493 80666 86557 80670
rect 86493 80610 86497 80666
rect 86497 80610 86553 80666
rect 86553 80610 86557 80666
rect 86493 80606 86557 80610
rect 86493 80586 86557 80590
rect 86493 80530 86497 80586
rect 86497 80530 86553 80586
rect 86553 80530 86557 80586
rect 86493 80526 86557 80530
rect 86493 80506 86557 80510
rect 86493 80450 86497 80506
rect 86497 80450 86553 80506
rect 86553 80450 86557 80506
rect 86493 80446 86557 80450
rect 86493 80426 86557 80430
rect 86493 80370 86497 80426
rect 86497 80370 86553 80426
rect 86553 80370 86557 80426
rect 86493 80366 86557 80370
rect 86493 80346 86557 80350
rect 86493 80290 86497 80346
rect 86497 80290 86553 80346
rect 86553 80290 86557 80346
rect 86493 80286 86557 80290
rect 86493 80266 86557 80270
rect 86493 80210 86497 80266
rect 86497 80210 86553 80266
rect 86553 80210 86557 80266
rect 86493 80206 86557 80210
rect 87581 80746 87645 80750
rect 87581 80690 87585 80746
rect 87585 80690 87641 80746
rect 87641 80690 87645 80746
rect 87581 80686 87645 80690
rect 87581 80666 87645 80670
rect 87581 80610 87585 80666
rect 87585 80610 87641 80666
rect 87641 80610 87645 80666
rect 87581 80606 87645 80610
rect 87581 80586 87645 80590
rect 87581 80530 87585 80586
rect 87585 80530 87641 80586
rect 87641 80530 87645 80586
rect 87581 80526 87645 80530
rect 87581 80506 87645 80510
rect 87581 80450 87585 80506
rect 87585 80450 87641 80506
rect 87641 80450 87645 80506
rect 87581 80446 87645 80450
rect 87581 80426 87645 80430
rect 87581 80370 87585 80426
rect 87585 80370 87641 80426
rect 87641 80370 87645 80426
rect 87581 80366 87645 80370
rect 87581 80346 87645 80350
rect 87581 80290 87585 80346
rect 87585 80290 87641 80346
rect 87641 80290 87645 80346
rect 87581 80286 87645 80290
rect 87581 80266 87645 80270
rect 87581 80210 87585 80266
rect 87585 80210 87641 80266
rect 87641 80210 87645 80266
rect 87581 80206 87645 80210
rect 88669 80746 88733 80750
rect 88669 80690 88673 80746
rect 88673 80690 88729 80746
rect 88729 80690 88733 80746
rect 88669 80686 88733 80690
rect 88669 80666 88733 80670
rect 88669 80610 88673 80666
rect 88673 80610 88729 80666
rect 88729 80610 88733 80666
rect 88669 80606 88733 80610
rect 88669 80586 88733 80590
rect 88669 80530 88673 80586
rect 88673 80530 88729 80586
rect 88729 80530 88733 80586
rect 88669 80526 88733 80530
rect 88669 80506 88733 80510
rect 88669 80450 88673 80506
rect 88673 80450 88729 80506
rect 88729 80450 88733 80506
rect 88669 80446 88733 80450
rect 88669 80426 88733 80430
rect 88669 80370 88673 80426
rect 88673 80370 88729 80426
rect 88729 80370 88733 80426
rect 88669 80366 88733 80370
rect 88669 80346 88733 80350
rect 88669 80290 88673 80346
rect 88673 80290 88729 80346
rect 88729 80290 88733 80346
rect 88669 80286 88733 80290
rect 88669 80266 88733 80270
rect 88669 80210 88673 80266
rect 88673 80210 88729 80266
rect 88729 80210 88733 80266
rect 88669 80206 88733 80210
rect 75070 78743 75134 78747
rect 75070 78687 75074 78743
rect 75074 78687 75130 78743
rect 75130 78687 75134 78743
rect 75070 78683 75134 78687
rect 75070 78663 75134 78667
rect 75070 78607 75074 78663
rect 75074 78607 75130 78663
rect 75130 78607 75134 78663
rect 75070 78603 75134 78607
rect 75070 78583 75134 78587
rect 75070 78527 75074 78583
rect 75074 78527 75130 78583
rect 75130 78527 75134 78583
rect 75070 78523 75134 78527
rect 75070 78503 75134 78507
rect 75070 78447 75074 78503
rect 75074 78447 75130 78503
rect 75130 78447 75134 78503
rect 75070 78443 75134 78447
rect 75070 78423 75134 78427
rect 75070 78367 75074 78423
rect 75074 78367 75130 78423
rect 75130 78367 75134 78423
rect 75070 78363 75134 78367
rect 75070 78343 75134 78347
rect 75070 78287 75074 78343
rect 75074 78287 75130 78343
rect 75130 78287 75134 78343
rect 75070 78283 75134 78287
rect 75070 78263 75134 78267
rect 75070 78207 75074 78263
rect 75074 78207 75130 78263
rect 75130 78207 75134 78263
rect 75070 78203 75134 78207
rect 76158 78743 76222 78747
rect 76158 78687 76162 78743
rect 76162 78687 76218 78743
rect 76218 78687 76222 78743
rect 76158 78683 76222 78687
rect 76158 78663 76222 78667
rect 76158 78607 76162 78663
rect 76162 78607 76218 78663
rect 76218 78607 76222 78663
rect 76158 78603 76222 78607
rect 76158 78583 76222 78587
rect 76158 78527 76162 78583
rect 76162 78527 76218 78583
rect 76218 78527 76222 78583
rect 76158 78523 76222 78527
rect 76158 78503 76222 78507
rect 76158 78447 76162 78503
rect 76162 78447 76218 78503
rect 76218 78447 76222 78503
rect 76158 78443 76222 78447
rect 76158 78423 76222 78427
rect 76158 78367 76162 78423
rect 76162 78367 76218 78423
rect 76218 78367 76222 78423
rect 76158 78363 76222 78367
rect 76158 78343 76222 78347
rect 76158 78287 76162 78343
rect 76162 78287 76218 78343
rect 76218 78287 76222 78343
rect 76158 78283 76222 78287
rect 76158 78263 76222 78267
rect 76158 78207 76162 78263
rect 76162 78207 76218 78263
rect 76218 78207 76222 78263
rect 76158 78203 76222 78207
rect 77246 78743 77310 78747
rect 77246 78687 77250 78743
rect 77250 78687 77306 78743
rect 77306 78687 77310 78743
rect 77246 78683 77310 78687
rect 77246 78663 77310 78667
rect 77246 78607 77250 78663
rect 77250 78607 77306 78663
rect 77306 78607 77310 78663
rect 77246 78603 77310 78607
rect 77246 78583 77310 78587
rect 77246 78527 77250 78583
rect 77250 78527 77306 78583
rect 77306 78527 77310 78583
rect 77246 78523 77310 78527
rect 77246 78503 77310 78507
rect 77246 78447 77250 78503
rect 77250 78447 77306 78503
rect 77306 78447 77310 78503
rect 77246 78443 77310 78447
rect 77246 78423 77310 78427
rect 77246 78367 77250 78423
rect 77250 78367 77306 78423
rect 77306 78367 77310 78423
rect 77246 78363 77310 78367
rect 77246 78343 77310 78347
rect 77246 78287 77250 78343
rect 77250 78287 77306 78343
rect 77306 78287 77310 78343
rect 77246 78283 77310 78287
rect 77246 78263 77310 78267
rect 77246 78207 77250 78263
rect 77250 78207 77306 78263
rect 77306 78207 77310 78263
rect 77246 78203 77310 78207
rect 78334 78743 78398 78747
rect 78334 78687 78338 78743
rect 78338 78687 78394 78743
rect 78394 78687 78398 78743
rect 78334 78683 78398 78687
rect 78334 78663 78398 78667
rect 78334 78607 78338 78663
rect 78338 78607 78394 78663
rect 78394 78607 78398 78663
rect 78334 78603 78398 78607
rect 78334 78583 78398 78587
rect 78334 78527 78338 78583
rect 78338 78527 78394 78583
rect 78394 78527 78398 78583
rect 78334 78523 78398 78527
rect 78334 78503 78398 78507
rect 78334 78447 78338 78503
rect 78338 78447 78394 78503
rect 78394 78447 78398 78503
rect 78334 78443 78398 78447
rect 78334 78423 78398 78427
rect 78334 78367 78338 78423
rect 78338 78367 78394 78423
rect 78394 78367 78398 78423
rect 78334 78363 78398 78367
rect 78334 78343 78398 78347
rect 78334 78287 78338 78343
rect 78338 78287 78394 78343
rect 78394 78287 78398 78343
rect 78334 78283 78398 78287
rect 78334 78263 78398 78267
rect 78334 78207 78338 78263
rect 78338 78207 78394 78263
rect 78394 78207 78398 78263
rect 78334 78203 78398 78207
rect 79422 78743 79486 78747
rect 79422 78687 79426 78743
rect 79426 78687 79482 78743
rect 79482 78687 79486 78743
rect 79422 78683 79486 78687
rect 79422 78663 79486 78667
rect 79422 78607 79426 78663
rect 79426 78607 79482 78663
rect 79482 78607 79486 78663
rect 79422 78603 79486 78607
rect 79422 78583 79486 78587
rect 79422 78527 79426 78583
rect 79426 78527 79482 78583
rect 79482 78527 79486 78583
rect 79422 78523 79486 78527
rect 79422 78503 79486 78507
rect 79422 78447 79426 78503
rect 79426 78447 79482 78503
rect 79482 78447 79486 78503
rect 79422 78443 79486 78447
rect 79422 78423 79486 78427
rect 79422 78367 79426 78423
rect 79426 78367 79482 78423
rect 79482 78367 79486 78423
rect 79422 78363 79486 78367
rect 79422 78343 79486 78347
rect 79422 78287 79426 78343
rect 79426 78287 79482 78343
rect 79482 78287 79486 78343
rect 79422 78283 79486 78287
rect 79422 78263 79486 78267
rect 79422 78207 79426 78263
rect 79426 78207 79482 78263
rect 79482 78207 79486 78263
rect 79422 78203 79486 78207
rect 80510 78743 80574 78747
rect 80510 78687 80514 78743
rect 80514 78687 80570 78743
rect 80570 78687 80574 78743
rect 80510 78683 80574 78687
rect 80510 78663 80574 78667
rect 80510 78607 80514 78663
rect 80514 78607 80570 78663
rect 80570 78607 80574 78663
rect 80510 78603 80574 78607
rect 80510 78583 80574 78587
rect 80510 78527 80514 78583
rect 80514 78527 80570 78583
rect 80570 78527 80574 78583
rect 80510 78523 80574 78527
rect 80510 78503 80574 78507
rect 80510 78447 80514 78503
rect 80514 78447 80570 78503
rect 80570 78447 80574 78503
rect 80510 78443 80574 78447
rect 80510 78423 80574 78427
rect 80510 78367 80514 78423
rect 80514 78367 80570 78423
rect 80570 78367 80574 78423
rect 80510 78363 80574 78367
rect 80510 78343 80574 78347
rect 80510 78287 80514 78343
rect 80514 78287 80570 78343
rect 80570 78287 80574 78343
rect 80510 78283 80574 78287
rect 80510 78263 80574 78267
rect 80510 78207 80514 78263
rect 80514 78207 80570 78263
rect 80570 78207 80574 78263
rect 80510 78203 80574 78207
rect 81598 78743 81662 78747
rect 81598 78687 81602 78743
rect 81602 78687 81658 78743
rect 81658 78687 81662 78743
rect 81598 78683 81662 78687
rect 81598 78663 81662 78667
rect 81598 78607 81602 78663
rect 81602 78607 81658 78663
rect 81658 78607 81662 78663
rect 81598 78603 81662 78607
rect 81598 78583 81662 78587
rect 81598 78527 81602 78583
rect 81602 78527 81658 78583
rect 81658 78527 81662 78583
rect 81598 78523 81662 78527
rect 81598 78503 81662 78507
rect 81598 78447 81602 78503
rect 81602 78447 81658 78503
rect 81658 78447 81662 78503
rect 81598 78443 81662 78447
rect 81598 78423 81662 78427
rect 81598 78367 81602 78423
rect 81602 78367 81658 78423
rect 81658 78367 81662 78423
rect 81598 78363 81662 78367
rect 81598 78343 81662 78347
rect 81598 78287 81602 78343
rect 81602 78287 81658 78343
rect 81658 78287 81662 78343
rect 81598 78283 81662 78287
rect 81598 78263 81662 78267
rect 81598 78207 81602 78263
rect 81602 78207 81658 78263
rect 81658 78207 81662 78263
rect 81598 78203 81662 78207
rect 82686 78743 82750 78747
rect 82686 78687 82690 78743
rect 82690 78687 82746 78743
rect 82746 78687 82750 78743
rect 82686 78683 82750 78687
rect 82686 78663 82750 78667
rect 82686 78607 82690 78663
rect 82690 78607 82746 78663
rect 82746 78607 82750 78663
rect 82686 78603 82750 78607
rect 82686 78583 82750 78587
rect 82686 78527 82690 78583
rect 82690 78527 82746 78583
rect 82746 78527 82750 78583
rect 82686 78523 82750 78527
rect 82686 78503 82750 78507
rect 82686 78447 82690 78503
rect 82690 78447 82746 78503
rect 82746 78447 82750 78503
rect 82686 78443 82750 78447
rect 82686 78423 82750 78427
rect 82686 78367 82690 78423
rect 82690 78367 82746 78423
rect 82746 78367 82750 78423
rect 82686 78363 82750 78367
rect 82686 78343 82750 78347
rect 82686 78287 82690 78343
rect 82690 78287 82746 78343
rect 82746 78287 82750 78343
rect 82686 78283 82750 78287
rect 82686 78263 82750 78267
rect 82686 78207 82690 78263
rect 82690 78207 82746 78263
rect 82746 78207 82750 78263
rect 82686 78203 82750 78207
rect 83774 78743 83838 78747
rect 83774 78687 83778 78743
rect 83778 78687 83834 78743
rect 83834 78687 83838 78743
rect 83774 78683 83838 78687
rect 83774 78663 83838 78667
rect 83774 78607 83778 78663
rect 83778 78607 83834 78663
rect 83834 78607 83838 78663
rect 83774 78603 83838 78607
rect 83774 78583 83838 78587
rect 83774 78527 83778 78583
rect 83778 78527 83834 78583
rect 83834 78527 83838 78583
rect 83774 78523 83838 78527
rect 83774 78503 83838 78507
rect 83774 78447 83778 78503
rect 83778 78447 83834 78503
rect 83834 78447 83838 78503
rect 83774 78443 83838 78447
rect 83774 78423 83838 78427
rect 83774 78367 83778 78423
rect 83778 78367 83834 78423
rect 83834 78367 83838 78423
rect 83774 78363 83838 78367
rect 83774 78343 83838 78347
rect 83774 78287 83778 78343
rect 83778 78287 83834 78343
rect 83834 78287 83838 78343
rect 83774 78283 83838 78287
rect 83774 78263 83838 78267
rect 83774 78207 83778 78263
rect 83778 78207 83834 78263
rect 83834 78207 83838 78263
rect 83774 78203 83838 78207
rect 84862 78743 84926 78747
rect 84862 78687 84866 78743
rect 84866 78687 84922 78743
rect 84922 78687 84926 78743
rect 84862 78683 84926 78687
rect 84862 78663 84926 78667
rect 84862 78607 84866 78663
rect 84866 78607 84922 78663
rect 84922 78607 84926 78663
rect 84862 78603 84926 78607
rect 84862 78583 84926 78587
rect 84862 78527 84866 78583
rect 84866 78527 84922 78583
rect 84922 78527 84926 78583
rect 84862 78523 84926 78527
rect 84862 78503 84926 78507
rect 84862 78447 84866 78503
rect 84866 78447 84922 78503
rect 84922 78447 84926 78503
rect 84862 78443 84926 78447
rect 84862 78423 84926 78427
rect 84862 78367 84866 78423
rect 84866 78367 84922 78423
rect 84922 78367 84926 78423
rect 84862 78363 84926 78367
rect 84862 78343 84926 78347
rect 84862 78287 84866 78343
rect 84866 78287 84922 78343
rect 84922 78287 84926 78343
rect 84862 78283 84926 78287
rect 84862 78263 84926 78267
rect 84862 78207 84866 78263
rect 84866 78207 84922 78263
rect 84922 78207 84926 78263
rect 84862 78203 84926 78207
rect 85950 78743 86014 78747
rect 85950 78687 85954 78743
rect 85954 78687 86010 78743
rect 86010 78687 86014 78743
rect 85950 78683 86014 78687
rect 85950 78663 86014 78667
rect 85950 78607 85954 78663
rect 85954 78607 86010 78663
rect 86010 78607 86014 78663
rect 85950 78603 86014 78607
rect 85950 78583 86014 78587
rect 85950 78527 85954 78583
rect 85954 78527 86010 78583
rect 86010 78527 86014 78583
rect 85950 78523 86014 78527
rect 85950 78503 86014 78507
rect 85950 78447 85954 78503
rect 85954 78447 86010 78503
rect 86010 78447 86014 78503
rect 85950 78443 86014 78447
rect 85950 78423 86014 78427
rect 85950 78367 85954 78423
rect 85954 78367 86010 78423
rect 86010 78367 86014 78423
rect 85950 78363 86014 78367
rect 85950 78343 86014 78347
rect 85950 78287 85954 78343
rect 85954 78287 86010 78343
rect 86010 78287 86014 78343
rect 85950 78283 86014 78287
rect 85950 78263 86014 78267
rect 85950 78207 85954 78263
rect 85954 78207 86010 78263
rect 86010 78207 86014 78263
rect 85950 78203 86014 78207
rect 87038 78743 87102 78747
rect 87038 78687 87042 78743
rect 87042 78687 87098 78743
rect 87098 78687 87102 78743
rect 87038 78683 87102 78687
rect 87038 78663 87102 78667
rect 87038 78607 87042 78663
rect 87042 78607 87098 78663
rect 87098 78607 87102 78663
rect 87038 78603 87102 78607
rect 87038 78583 87102 78587
rect 87038 78527 87042 78583
rect 87042 78527 87098 78583
rect 87098 78527 87102 78583
rect 87038 78523 87102 78527
rect 87038 78503 87102 78507
rect 87038 78447 87042 78503
rect 87042 78447 87098 78503
rect 87098 78447 87102 78503
rect 87038 78443 87102 78447
rect 87038 78423 87102 78427
rect 87038 78367 87042 78423
rect 87042 78367 87098 78423
rect 87098 78367 87102 78423
rect 87038 78363 87102 78367
rect 87038 78343 87102 78347
rect 87038 78287 87042 78343
rect 87042 78287 87098 78343
rect 87098 78287 87102 78343
rect 87038 78283 87102 78287
rect 87038 78263 87102 78267
rect 87038 78207 87042 78263
rect 87042 78207 87098 78263
rect 87098 78207 87102 78263
rect 87038 78203 87102 78207
rect 88126 78743 88190 78747
rect 88126 78687 88130 78743
rect 88130 78687 88186 78743
rect 88186 78687 88190 78743
rect 88126 78683 88190 78687
rect 88126 78663 88190 78667
rect 88126 78607 88130 78663
rect 88130 78607 88186 78663
rect 88186 78607 88190 78663
rect 88126 78603 88190 78607
rect 88126 78583 88190 78587
rect 88126 78527 88130 78583
rect 88130 78527 88186 78583
rect 88186 78527 88190 78583
rect 88126 78523 88190 78527
rect 88126 78503 88190 78507
rect 88126 78447 88130 78503
rect 88130 78447 88186 78503
rect 88186 78447 88190 78503
rect 88126 78443 88190 78447
rect 88126 78423 88190 78427
rect 88126 78367 88130 78423
rect 88130 78367 88186 78423
rect 88186 78367 88190 78423
rect 88126 78363 88190 78367
rect 88126 78343 88190 78347
rect 88126 78287 88130 78343
rect 88130 78287 88186 78343
rect 88186 78287 88190 78343
rect 88126 78283 88190 78287
rect 88126 78263 88190 78267
rect 88126 78207 88130 78263
rect 88130 78207 88186 78263
rect 88186 78207 88190 78263
rect 88126 78203 88190 78207
rect 74525 76746 74589 76750
rect 74525 76690 74529 76746
rect 74529 76690 74585 76746
rect 74585 76690 74589 76746
rect 74525 76686 74589 76690
rect 74525 76666 74589 76670
rect 74525 76610 74529 76666
rect 74529 76610 74585 76666
rect 74585 76610 74589 76666
rect 74525 76606 74589 76610
rect 74525 76586 74589 76590
rect 74525 76530 74529 76586
rect 74529 76530 74585 76586
rect 74585 76530 74589 76586
rect 74525 76526 74589 76530
rect 74525 76506 74589 76510
rect 74525 76450 74529 76506
rect 74529 76450 74585 76506
rect 74585 76450 74589 76506
rect 74525 76446 74589 76450
rect 74525 76426 74589 76430
rect 74525 76370 74529 76426
rect 74529 76370 74585 76426
rect 74585 76370 74589 76426
rect 74525 76366 74589 76370
rect 74525 76346 74589 76350
rect 74525 76290 74529 76346
rect 74529 76290 74585 76346
rect 74585 76290 74589 76346
rect 74525 76286 74589 76290
rect 74525 76266 74589 76270
rect 74525 76210 74529 76266
rect 74529 76210 74585 76266
rect 74585 76210 74589 76266
rect 74525 76206 74589 76210
rect 75613 76746 75677 76750
rect 75613 76690 75617 76746
rect 75617 76690 75673 76746
rect 75673 76690 75677 76746
rect 75613 76686 75677 76690
rect 75613 76666 75677 76670
rect 75613 76610 75617 76666
rect 75617 76610 75673 76666
rect 75673 76610 75677 76666
rect 75613 76606 75677 76610
rect 75613 76586 75677 76590
rect 75613 76530 75617 76586
rect 75617 76530 75673 76586
rect 75673 76530 75677 76586
rect 75613 76526 75677 76530
rect 75613 76506 75677 76510
rect 75613 76450 75617 76506
rect 75617 76450 75673 76506
rect 75673 76450 75677 76506
rect 75613 76446 75677 76450
rect 75613 76426 75677 76430
rect 75613 76370 75617 76426
rect 75617 76370 75673 76426
rect 75673 76370 75677 76426
rect 75613 76366 75677 76370
rect 75613 76346 75677 76350
rect 75613 76290 75617 76346
rect 75617 76290 75673 76346
rect 75673 76290 75677 76346
rect 75613 76286 75677 76290
rect 75613 76266 75677 76270
rect 75613 76210 75617 76266
rect 75617 76210 75673 76266
rect 75673 76210 75677 76266
rect 75613 76206 75677 76210
rect 76701 76746 76765 76750
rect 76701 76690 76705 76746
rect 76705 76690 76761 76746
rect 76761 76690 76765 76746
rect 76701 76686 76765 76690
rect 76701 76666 76765 76670
rect 76701 76610 76705 76666
rect 76705 76610 76761 76666
rect 76761 76610 76765 76666
rect 76701 76606 76765 76610
rect 76701 76586 76765 76590
rect 76701 76530 76705 76586
rect 76705 76530 76761 76586
rect 76761 76530 76765 76586
rect 76701 76526 76765 76530
rect 76701 76506 76765 76510
rect 76701 76450 76705 76506
rect 76705 76450 76761 76506
rect 76761 76450 76765 76506
rect 76701 76446 76765 76450
rect 76701 76426 76765 76430
rect 76701 76370 76705 76426
rect 76705 76370 76761 76426
rect 76761 76370 76765 76426
rect 76701 76366 76765 76370
rect 76701 76346 76765 76350
rect 76701 76290 76705 76346
rect 76705 76290 76761 76346
rect 76761 76290 76765 76346
rect 76701 76286 76765 76290
rect 76701 76266 76765 76270
rect 76701 76210 76705 76266
rect 76705 76210 76761 76266
rect 76761 76210 76765 76266
rect 76701 76206 76765 76210
rect 77789 76746 77853 76750
rect 77789 76690 77793 76746
rect 77793 76690 77849 76746
rect 77849 76690 77853 76746
rect 77789 76686 77853 76690
rect 77789 76666 77853 76670
rect 77789 76610 77793 76666
rect 77793 76610 77849 76666
rect 77849 76610 77853 76666
rect 77789 76606 77853 76610
rect 77789 76586 77853 76590
rect 77789 76530 77793 76586
rect 77793 76530 77849 76586
rect 77849 76530 77853 76586
rect 77789 76526 77853 76530
rect 77789 76506 77853 76510
rect 77789 76450 77793 76506
rect 77793 76450 77849 76506
rect 77849 76450 77853 76506
rect 77789 76446 77853 76450
rect 77789 76426 77853 76430
rect 77789 76370 77793 76426
rect 77793 76370 77849 76426
rect 77849 76370 77853 76426
rect 77789 76366 77853 76370
rect 77789 76346 77853 76350
rect 77789 76290 77793 76346
rect 77793 76290 77849 76346
rect 77849 76290 77853 76346
rect 77789 76286 77853 76290
rect 77789 76266 77853 76270
rect 77789 76210 77793 76266
rect 77793 76210 77849 76266
rect 77849 76210 77853 76266
rect 77789 76206 77853 76210
rect 78877 76746 78941 76750
rect 78877 76690 78881 76746
rect 78881 76690 78937 76746
rect 78937 76690 78941 76746
rect 78877 76686 78941 76690
rect 78877 76666 78941 76670
rect 78877 76610 78881 76666
rect 78881 76610 78937 76666
rect 78937 76610 78941 76666
rect 78877 76606 78941 76610
rect 78877 76586 78941 76590
rect 78877 76530 78881 76586
rect 78881 76530 78937 76586
rect 78937 76530 78941 76586
rect 78877 76526 78941 76530
rect 78877 76506 78941 76510
rect 78877 76450 78881 76506
rect 78881 76450 78937 76506
rect 78937 76450 78941 76506
rect 78877 76446 78941 76450
rect 78877 76426 78941 76430
rect 78877 76370 78881 76426
rect 78881 76370 78937 76426
rect 78937 76370 78941 76426
rect 78877 76366 78941 76370
rect 78877 76346 78941 76350
rect 78877 76290 78881 76346
rect 78881 76290 78937 76346
rect 78937 76290 78941 76346
rect 78877 76286 78941 76290
rect 78877 76266 78941 76270
rect 78877 76210 78881 76266
rect 78881 76210 78937 76266
rect 78937 76210 78941 76266
rect 78877 76206 78941 76210
rect 79965 76746 80029 76750
rect 79965 76690 79969 76746
rect 79969 76690 80025 76746
rect 80025 76690 80029 76746
rect 79965 76686 80029 76690
rect 79965 76666 80029 76670
rect 79965 76610 79969 76666
rect 79969 76610 80025 76666
rect 80025 76610 80029 76666
rect 79965 76606 80029 76610
rect 79965 76586 80029 76590
rect 79965 76530 79969 76586
rect 79969 76530 80025 76586
rect 80025 76530 80029 76586
rect 79965 76526 80029 76530
rect 79965 76506 80029 76510
rect 79965 76450 79969 76506
rect 79969 76450 80025 76506
rect 80025 76450 80029 76506
rect 79965 76446 80029 76450
rect 79965 76426 80029 76430
rect 79965 76370 79969 76426
rect 79969 76370 80025 76426
rect 80025 76370 80029 76426
rect 79965 76366 80029 76370
rect 79965 76346 80029 76350
rect 79965 76290 79969 76346
rect 79969 76290 80025 76346
rect 80025 76290 80029 76346
rect 79965 76286 80029 76290
rect 79965 76266 80029 76270
rect 79965 76210 79969 76266
rect 79969 76210 80025 76266
rect 80025 76210 80029 76266
rect 79965 76206 80029 76210
rect 81053 76746 81117 76750
rect 81053 76690 81057 76746
rect 81057 76690 81113 76746
rect 81113 76690 81117 76746
rect 81053 76686 81117 76690
rect 81053 76666 81117 76670
rect 81053 76610 81057 76666
rect 81057 76610 81113 76666
rect 81113 76610 81117 76666
rect 81053 76606 81117 76610
rect 81053 76586 81117 76590
rect 81053 76530 81057 76586
rect 81057 76530 81113 76586
rect 81113 76530 81117 76586
rect 81053 76526 81117 76530
rect 81053 76506 81117 76510
rect 81053 76450 81057 76506
rect 81057 76450 81113 76506
rect 81113 76450 81117 76506
rect 81053 76446 81117 76450
rect 81053 76426 81117 76430
rect 81053 76370 81057 76426
rect 81057 76370 81113 76426
rect 81113 76370 81117 76426
rect 81053 76366 81117 76370
rect 81053 76346 81117 76350
rect 81053 76290 81057 76346
rect 81057 76290 81113 76346
rect 81113 76290 81117 76346
rect 81053 76286 81117 76290
rect 81053 76266 81117 76270
rect 81053 76210 81057 76266
rect 81057 76210 81113 76266
rect 81113 76210 81117 76266
rect 81053 76206 81117 76210
rect 82141 76746 82205 76750
rect 82141 76690 82145 76746
rect 82145 76690 82201 76746
rect 82201 76690 82205 76746
rect 82141 76686 82205 76690
rect 82141 76666 82205 76670
rect 82141 76610 82145 76666
rect 82145 76610 82201 76666
rect 82201 76610 82205 76666
rect 82141 76606 82205 76610
rect 82141 76586 82205 76590
rect 82141 76530 82145 76586
rect 82145 76530 82201 76586
rect 82201 76530 82205 76586
rect 82141 76526 82205 76530
rect 82141 76506 82205 76510
rect 82141 76450 82145 76506
rect 82145 76450 82201 76506
rect 82201 76450 82205 76506
rect 82141 76446 82205 76450
rect 82141 76426 82205 76430
rect 82141 76370 82145 76426
rect 82145 76370 82201 76426
rect 82201 76370 82205 76426
rect 82141 76366 82205 76370
rect 82141 76346 82205 76350
rect 82141 76290 82145 76346
rect 82145 76290 82201 76346
rect 82201 76290 82205 76346
rect 82141 76286 82205 76290
rect 82141 76266 82205 76270
rect 82141 76210 82145 76266
rect 82145 76210 82201 76266
rect 82201 76210 82205 76266
rect 82141 76206 82205 76210
rect 83229 76746 83293 76750
rect 83229 76690 83233 76746
rect 83233 76690 83289 76746
rect 83289 76690 83293 76746
rect 83229 76686 83293 76690
rect 83229 76666 83293 76670
rect 83229 76610 83233 76666
rect 83233 76610 83289 76666
rect 83289 76610 83293 76666
rect 83229 76606 83293 76610
rect 83229 76586 83293 76590
rect 83229 76530 83233 76586
rect 83233 76530 83289 76586
rect 83289 76530 83293 76586
rect 83229 76526 83293 76530
rect 83229 76506 83293 76510
rect 83229 76450 83233 76506
rect 83233 76450 83289 76506
rect 83289 76450 83293 76506
rect 83229 76446 83293 76450
rect 83229 76426 83293 76430
rect 83229 76370 83233 76426
rect 83233 76370 83289 76426
rect 83289 76370 83293 76426
rect 83229 76366 83293 76370
rect 83229 76346 83293 76350
rect 83229 76290 83233 76346
rect 83233 76290 83289 76346
rect 83289 76290 83293 76346
rect 83229 76286 83293 76290
rect 83229 76266 83293 76270
rect 83229 76210 83233 76266
rect 83233 76210 83289 76266
rect 83289 76210 83293 76266
rect 83229 76206 83293 76210
rect 84317 76746 84381 76750
rect 84317 76690 84321 76746
rect 84321 76690 84377 76746
rect 84377 76690 84381 76746
rect 84317 76686 84381 76690
rect 84317 76666 84381 76670
rect 84317 76610 84321 76666
rect 84321 76610 84377 76666
rect 84377 76610 84381 76666
rect 84317 76606 84381 76610
rect 84317 76586 84381 76590
rect 84317 76530 84321 76586
rect 84321 76530 84377 76586
rect 84377 76530 84381 76586
rect 84317 76526 84381 76530
rect 84317 76506 84381 76510
rect 84317 76450 84321 76506
rect 84321 76450 84377 76506
rect 84377 76450 84381 76506
rect 84317 76446 84381 76450
rect 84317 76426 84381 76430
rect 84317 76370 84321 76426
rect 84321 76370 84377 76426
rect 84377 76370 84381 76426
rect 84317 76366 84381 76370
rect 84317 76346 84381 76350
rect 84317 76290 84321 76346
rect 84321 76290 84377 76346
rect 84377 76290 84381 76346
rect 84317 76286 84381 76290
rect 84317 76266 84381 76270
rect 84317 76210 84321 76266
rect 84321 76210 84377 76266
rect 84377 76210 84381 76266
rect 84317 76206 84381 76210
rect 85405 76746 85469 76750
rect 85405 76690 85409 76746
rect 85409 76690 85465 76746
rect 85465 76690 85469 76746
rect 85405 76686 85469 76690
rect 85405 76666 85469 76670
rect 85405 76610 85409 76666
rect 85409 76610 85465 76666
rect 85465 76610 85469 76666
rect 85405 76606 85469 76610
rect 85405 76586 85469 76590
rect 85405 76530 85409 76586
rect 85409 76530 85465 76586
rect 85465 76530 85469 76586
rect 85405 76526 85469 76530
rect 85405 76506 85469 76510
rect 85405 76450 85409 76506
rect 85409 76450 85465 76506
rect 85465 76450 85469 76506
rect 85405 76446 85469 76450
rect 85405 76426 85469 76430
rect 85405 76370 85409 76426
rect 85409 76370 85465 76426
rect 85465 76370 85469 76426
rect 85405 76366 85469 76370
rect 85405 76346 85469 76350
rect 85405 76290 85409 76346
rect 85409 76290 85465 76346
rect 85465 76290 85469 76346
rect 85405 76286 85469 76290
rect 85405 76266 85469 76270
rect 85405 76210 85409 76266
rect 85409 76210 85465 76266
rect 85465 76210 85469 76266
rect 85405 76206 85469 76210
rect 86493 76746 86557 76750
rect 86493 76690 86497 76746
rect 86497 76690 86553 76746
rect 86553 76690 86557 76746
rect 86493 76686 86557 76690
rect 86493 76666 86557 76670
rect 86493 76610 86497 76666
rect 86497 76610 86553 76666
rect 86553 76610 86557 76666
rect 86493 76606 86557 76610
rect 86493 76586 86557 76590
rect 86493 76530 86497 76586
rect 86497 76530 86553 76586
rect 86553 76530 86557 76586
rect 86493 76526 86557 76530
rect 86493 76506 86557 76510
rect 86493 76450 86497 76506
rect 86497 76450 86553 76506
rect 86553 76450 86557 76506
rect 86493 76446 86557 76450
rect 86493 76426 86557 76430
rect 86493 76370 86497 76426
rect 86497 76370 86553 76426
rect 86553 76370 86557 76426
rect 86493 76366 86557 76370
rect 86493 76346 86557 76350
rect 86493 76290 86497 76346
rect 86497 76290 86553 76346
rect 86553 76290 86557 76346
rect 86493 76286 86557 76290
rect 86493 76266 86557 76270
rect 86493 76210 86497 76266
rect 86497 76210 86553 76266
rect 86553 76210 86557 76266
rect 86493 76206 86557 76210
rect 87581 76746 87645 76750
rect 87581 76690 87585 76746
rect 87585 76690 87641 76746
rect 87641 76690 87645 76746
rect 87581 76686 87645 76690
rect 87581 76666 87645 76670
rect 87581 76610 87585 76666
rect 87585 76610 87641 76666
rect 87641 76610 87645 76666
rect 87581 76606 87645 76610
rect 87581 76586 87645 76590
rect 87581 76530 87585 76586
rect 87585 76530 87641 76586
rect 87641 76530 87645 76586
rect 87581 76526 87645 76530
rect 87581 76506 87645 76510
rect 87581 76450 87585 76506
rect 87585 76450 87641 76506
rect 87641 76450 87645 76506
rect 87581 76446 87645 76450
rect 87581 76426 87645 76430
rect 87581 76370 87585 76426
rect 87585 76370 87641 76426
rect 87641 76370 87645 76426
rect 87581 76366 87645 76370
rect 87581 76346 87645 76350
rect 87581 76290 87585 76346
rect 87585 76290 87641 76346
rect 87641 76290 87645 76346
rect 87581 76286 87645 76290
rect 87581 76266 87645 76270
rect 87581 76210 87585 76266
rect 87585 76210 87641 76266
rect 87641 76210 87645 76266
rect 87581 76206 87645 76210
rect 88669 76746 88733 76750
rect 88669 76690 88673 76746
rect 88673 76690 88729 76746
rect 88729 76690 88733 76746
rect 88669 76686 88733 76690
rect 88669 76666 88733 76670
rect 88669 76610 88673 76666
rect 88673 76610 88729 76666
rect 88729 76610 88733 76666
rect 88669 76606 88733 76610
rect 88669 76586 88733 76590
rect 88669 76530 88673 76586
rect 88673 76530 88729 76586
rect 88729 76530 88733 76586
rect 88669 76526 88733 76530
rect 88669 76506 88733 76510
rect 88669 76450 88673 76506
rect 88673 76450 88729 76506
rect 88729 76450 88733 76506
rect 88669 76446 88733 76450
rect 88669 76426 88733 76430
rect 88669 76370 88673 76426
rect 88673 76370 88729 76426
rect 88729 76370 88733 76426
rect 88669 76366 88733 76370
rect 88669 76346 88733 76350
rect 88669 76290 88673 76346
rect 88673 76290 88729 76346
rect 88729 76290 88733 76346
rect 88669 76286 88733 76290
rect 88669 76266 88733 76270
rect 88669 76210 88673 76266
rect 88673 76210 88729 76266
rect 88729 76210 88733 76266
rect 88669 76206 88733 76210
rect 75070 74743 75134 74747
rect 75070 74687 75074 74743
rect 75074 74687 75130 74743
rect 75130 74687 75134 74743
rect 75070 74683 75134 74687
rect 75070 74663 75134 74667
rect 75070 74607 75074 74663
rect 75074 74607 75130 74663
rect 75130 74607 75134 74663
rect 75070 74603 75134 74607
rect 75070 74583 75134 74587
rect 75070 74527 75074 74583
rect 75074 74527 75130 74583
rect 75130 74527 75134 74583
rect 75070 74523 75134 74527
rect 75070 74503 75134 74507
rect 75070 74447 75074 74503
rect 75074 74447 75130 74503
rect 75130 74447 75134 74503
rect 75070 74443 75134 74447
rect 75070 74423 75134 74427
rect 75070 74367 75074 74423
rect 75074 74367 75130 74423
rect 75130 74367 75134 74423
rect 75070 74363 75134 74367
rect 75070 74343 75134 74347
rect 75070 74287 75074 74343
rect 75074 74287 75130 74343
rect 75130 74287 75134 74343
rect 75070 74283 75134 74287
rect 75070 74263 75134 74267
rect 75070 74207 75074 74263
rect 75074 74207 75130 74263
rect 75130 74207 75134 74263
rect 75070 74203 75134 74207
rect 77246 74743 77310 74747
rect 77246 74687 77250 74743
rect 77250 74687 77306 74743
rect 77306 74687 77310 74743
rect 77246 74683 77310 74687
rect 77246 74663 77310 74667
rect 77246 74607 77250 74663
rect 77250 74607 77306 74663
rect 77306 74607 77310 74663
rect 77246 74603 77310 74607
rect 77246 74583 77310 74587
rect 77246 74527 77250 74583
rect 77250 74527 77306 74583
rect 77306 74527 77310 74583
rect 77246 74523 77310 74527
rect 77246 74503 77310 74507
rect 77246 74447 77250 74503
rect 77250 74447 77306 74503
rect 77306 74447 77310 74503
rect 77246 74443 77310 74447
rect 77246 74423 77310 74427
rect 77246 74367 77250 74423
rect 77250 74367 77306 74423
rect 77306 74367 77310 74423
rect 77246 74363 77310 74367
rect 77246 74343 77310 74347
rect 77246 74287 77250 74343
rect 77250 74287 77306 74343
rect 77306 74287 77310 74343
rect 77246 74283 77310 74287
rect 77246 74263 77310 74267
rect 77246 74207 77250 74263
rect 77250 74207 77306 74263
rect 77306 74207 77310 74263
rect 77246 74203 77310 74207
rect 78334 74743 78398 74747
rect 78334 74687 78338 74743
rect 78338 74687 78394 74743
rect 78394 74687 78398 74743
rect 78334 74683 78398 74687
rect 78334 74663 78398 74667
rect 78334 74607 78338 74663
rect 78338 74607 78394 74663
rect 78394 74607 78398 74663
rect 78334 74603 78398 74607
rect 78334 74583 78398 74587
rect 78334 74527 78338 74583
rect 78338 74527 78394 74583
rect 78394 74527 78398 74583
rect 78334 74523 78398 74527
rect 78334 74503 78398 74507
rect 78334 74447 78338 74503
rect 78338 74447 78394 74503
rect 78394 74447 78398 74503
rect 78334 74443 78398 74447
rect 78334 74423 78398 74427
rect 78334 74367 78338 74423
rect 78338 74367 78394 74423
rect 78394 74367 78398 74423
rect 78334 74363 78398 74367
rect 78334 74343 78398 74347
rect 78334 74287 78338 74343
rect 78338 74287 78394 74343
rect 78394 74287 78398 74343
rect 78334 74283 78398 74287
rect 78334 74263 78398 74267
rect 78334 74207 78338 74263
rect 78338 74207 78394 74263
rect 78394 74207 78398 74263
rect 78334 74203 78398 74207
rect 80510 74743 80574 74747
rect 80510 74687 80514 74743
rect 80514 74687 80570 74743
rect 80570 74687 80574 74743
rect 80510 74683 80574 74687
rect 80510 74663 80574 74667
rect 80510 74607 80514 74663
rect 80514 74607 80570 74663
rect 80570 74607 80574 74663
rect 80510 74603 80574 74607
rect 80510 74583 80574 74587
rect 80510 74527 80514 74583
rect 80514 74527 80570 74583
rect 80570 74527 80574 74583
rect 80510 74523 80574 74527
rect 80510 74503 80574 74507
rect 80510 74447 80514 74503
rect 80514 74447 80570 74503
rect 80570 74447 80574 74503
rect 80510 74443 80574 74447
rect 80510 74423 80574 74427
rect 80510 74367 80514 74423
rect 80514 74367 80570 74423
rect 80570 74367 80574 74423
rect 80510 74363 80574 74367
rect 80510 74343 80574 74347
rect 80510 74287 80514 74343
rect 80514 74287 80570 74343
rect 80570 74287 80574 74343
rect 80510 74283 80574 74287
rect 80510 74263 80574 74267
rect 80510 74207 80514 74263
rect 80514 74207 80570 74263
rect 80570 74207 80574 74263
rect 80510 74203 80574 74207
rect 81598 74743 81662 74747
rect 81598 74687 81602 74743
rect 81602 74687 81658 74743
rect 81658 74687 81662 74743
rect 81598 74683 81662 74687
rect 81598 74663 81662 74667
rect 81598 74607 81602 74663
rect 81602 74607 81658 74663
rect 81658 74607 81662 74663
rect 81598 74603 81662 74607
rect 81598 74583 81662 74587
rect 81598 74527 81602 74583
rect 81602 74527 81658 74583
rect 81658 74527 81662 74583
rect 81598 74523 81662 74527
rect 81598 74503 81662 74507
rect 81598 74447 81602 74503
rect 81602 74447 81658 74503
rect 81658 74447 81662 74503
rect 81598 74443 81662 74447
rect 81598 74423 81662 74427
rect 81598 74367 81602 74423
rect 81602 74367 81658 74423
rect 81658 74367 81662 74423
rect 81598 74363 81662 74367
rect 81598 74343 81662 74347
rect 81598 74287 81602 74343
rect 81602 74287 81658 74343
rect 81658 74287 81662 74343
rect 81598 74283 81662 74287
rect 81598 74263 81662 74267
rect 81598 74207 81602 74263
rect 81602 74207 81658 74263
rect 81658 74207 81662 74263
rect 81598 74203 81662 74207
rect 82686 74743 82750 74747
rect 82686 74687 82690 74743
rect 82690 74687 82746 74743
rect 82746 74687 82750 74743
rect 82686 74683 82750 74687
rect 82686 74663 82750 74667
rect 82686 74607 82690 74663
rect 82690 74607 82746 74663
rect 82746 74607 82750 74663
rect 82686 74603 82750 74607
rect 82686 74583 82750 74587
rect 82686 74527 82690 74583
rect 82690 74527 82746 74583
rect 82746 74527 82750 74583
rect 82686 74523 82750 74527
rect 82686 74503 82750 74507
rect 82686 74447 82690 74503
rect 82690 74447 82746 74503
rect 82746 74447 82750 74503
rect 82686 74443 82750 74447
rect 82686 74423 82750 74427
rect 82686 74367 82690 74423
rect 82690 74367 82746 74423
rect 82746 74367 82750 74423
rect 82686 74363 82750 74367
rect 82686 74343 82750 74347
rect 82686 74287 82690 74343
rect 82690 74287 82746 74343
rect 82746 74287 82750 74343
rect 82686 74283 82750 74287
rect 82686 74263 82750 74267
rect 82686 74207 82690 74263
rect 82690 74207 82746 74263
rect 82746 74207 82750 74263
rect 82686 74203 82750 74207
rect 84862 74743 84926 74747
rect 84862 74687 84866 74743
rect 84866 74687 84922 74743
rect 84922 74687 84926 74743
rect 84862 74683 84926 74687
rect 84862 74663 84926 74667
rect 84862 74607 84866 74663
rect 84866 74607 84922 74663
rect 84922 74607 84926 74663
rect 84862 74603 84926 74607
rect 84862 74583 84926 74587
rect 84862 74527 84866 74583
rect 84866 74527 84922 74583
rect 84922 74527 84926 74583
rect 84862 74523 84926 74527
rect 84862 74503 84926 74507
rect 84862 74447 84866 74503
rect 84866 74447 84922 74503
rect 84922 74447 84926 74503
rect 84862 74443 84926 74447
rect 84862 74423 84926 74427
rect 84862 74367 84866 74423
rect 84866 74367 84922 74423
rect 84922 74367 84926 74423
rect 84862 74363 84926 74367
rect 84862 74343 84926 74347
rect 84862 74287 84866 74343
rect 84866 74287 84922 74343
rect 84922 74287 84926 74343
rect 84862 74283 84926 74287
rect 84862 74263 84926 74267
rect 84862 74207 84866 74263
rect 84866 74207 84922 74263
rect 84922 74207 84926 74263
rect 84862 74203 84926 74207
rect 85950 74743 86014 74747
rect 85950 74687 85954 74743
rect 85954 74687 86010 74743
rect 86010 74687 86014 74743
rect 85950 74683 86014 74687
rect 85950 74663 86014 74667
rect 85950 74607 85954 74663
rect 85954 74607 86010 74663
rect 86010 74607 86014 74663
rect 85950 74603 86014 74607
rect 85950 74583 86014 74587
rect 85950 74527 85954 74583
rect 85954 74527 86010 74583
rect 86010 74527 86014 74583
rect 85950 74523 86014 74527
rect 85950 74503 86014 74507
rect 85950 74447 85954 74503
rect 85954 74447 86010 74503
rect 86010 74447 86014 74503
rect 85950 74443 86014 74447
rect 85950 74423 86014 74427
rect 85950 74367 85954 74423
rect 85954 74367 86010 74423
rect 86010 74367 86014 74423
rect 85950 74363 86014 74367
rect 85950 74343 86014 74347
rect 85950 74287 85954 74343
rect 85954 74287 86010 74343
rect 86010 74287 86014 74343
rect 85950 74283 86014 74287
rect 85950 74263 86014 74267
rect 85950 74207 85954 74263
rect 85954 74207 86010 74263
rect 86010 74207 86014 74263
rect 85950 74203 86014 74207
rect 88126 74743 88190 74747
rect 88126 74687 88130 74743
rect 88130 74687 88186 74743
rect 88186 74687 88190 74743
rect 88126 74683 88190 74687
rect 88126 74663 88190 74667
rect 88126 74607 88130 74663
rect 88130 74607 88186 74663
rect 88186 74607 88190 74663
rect 88126 74603 88190 74607
rect 88126 74583 88190 74587
rect 88126 74527 88130 74583
rect 88130 74527 88186 74583
rect 88186 74527 88190 74583
rect 88126 74523 88190 74527
rect 88126 74503 88190 74507
rect 88126 74447 88130 74503
rect 88130 74447 88186 74503
rect 88186 74447 88190 74503
rect 88126 74443 88190 74447
rect 88126 74423 88190 74427
rect 88126 74367 88130 74423
rect 88130 74367 88186 74423
rect 88186 74367 88190 74423
rect 88126 74363 88190 74367
rect 88126 74343 88190 74347
rect 88126 74287 88130 74343
rect 88130 74287 88186 74343
rect 88186 74287 88190 74343
rect 88126 74283 88190 74287
rect 88126 74263 88190 74267
rect 88126 74207 88130 74263
rect 88130 74207 88186 74263
rect 88186 74207 88190 74263
rect 88126 74203 88190 74207
rect 74525 72746 74589 72750
rect 74525 72690 74529 72746
rect 74529 72690 74585 72746
rect 74585 72690 74589 72746
rect 74525 72686 74589 72690
rect 74525 72666 74589 72670
rect 74525 72610 74529 72666
rect 74529 72610 74585 72666
rect 74585 72610 74589 72666
rect 74525 72606 74589 72610
rect 74525 72586 74589 72590
rect 74525 72530 74529 72586
rect 74529 72530 74585 72586
rect 74585 72530 74589 72586
rect 74525 72526 74589 72530
rect 74525 72506 74589 72510
rect 74525 72450 74529 72506
rect 74529 72450 74585 72506
rect 74585 72450 74589 72506
rect 74525 72446 74589 72450
rect 74525 72426 74589 72430
rect 74525 72370 74529 72426
rect 74529 72370 74585 72426
rect 74585 72370 74589 72426
rect 74525 72366 74589 72370
rect 74525 72346 74589 72350
rect 74525 72290 74529 72346
rect 74529 72290 74585 72346
rect 74585 72290 74589 72346
rect 74525 72286 74589 72290
rect 74525 72266 74589 72270
rect 74525 72210 74529 72266
rect 74529 72210 74585 72266
rect 74585 72210 74589 72266
rect 74525 72206 74589 72210
rect 75613 72746 75677 72750
rect 75613 72690 75617 72746
rect 75617 72690 75673 72746
rect 75673 72690 75677 72746
rect 75613 72686 75677 72690
rect 75613 72666 75677 72670
rect 75613 72610 75617 72666
rect 75617 72610 75673 72666
rect 75673 72610 75677 72666
rect 75613 72606 75677 72610
rect 75613 72586 75677 72590
rect 75613 72530 75617 72586
rect 75617 72530 75673 72586
rect 75673 72530 75677 72586
rect 75613 72526 75677 72530
rect 75613 72506 75677 72510
rect 75613 72450 75617 72506
rect 75617 72450 75673 72506
rect 75673 72450 75677 72506
rect 75613 72446 75677 72450
rect 75613 72426 75677 72430
rect 75613 72370 75617 72426
rect 75617 72370 75673 72426
rect 75673 72370 75677 72426
rect 75613 72366 75677 72370
rect 75613 72346 75677 72350
rect 75613 72290 75617 72346
rect 75617 72290 75673 72346
rect 75673 72290 75677 72346
rect 75613 72286 75677 72290
rect 75613 72266 75677 72270
rect 75613 72210 75617 72266
rect 75617 72210 75673 72266
rect 75673 72210 75677 72266
rect 75613 72206 75677 72210
rect 76701 72746 76765 72750
rect 76701 72690 76705 72746
rect 76705 72690 76761 72746
rect 76761 72690 76765 72746
rect 76701 72686 76765 72690
rect 76701 72666 76765 72670
rect 76701 72610 76705 72666
rect 76705 72610 76761 72666
rect 76761 72610 76765 72666
rect 76701 72606 76765 72610
rect 76701 72586 76765 72590
rect 76701 72530 76705 72586
rect 76705 72530 76761 72586
rect 76761 72530 76765 72586
rect 76701 72526 76765 72530
rect 76701 72506 76765 72510
rect 76701 72450 76705 72506
rect 76705 72450 76761 72506
rect 76761 72450 76765 72506
rect 76701 72446 76765 72450
rect 76701 72426 76765 72430
rect 76701 72370 76705 72426
rect 76705 72370 76761 72426
rect 76761 72370 76765 72426
rect 76701 72366 76765 72370
rect 76701 72346 76765 72350
rect 76701 72290 76705 72346
rect 76705 72290 76761 72346
rect 76761 72290 76765 72346
rect 76701 72286 76765 72290
rect 76701 72266 76765 72270
rect 76701 72210 76705 72266
rect 76705 72210 76761 72266
rect 76761 72210 76765 72266
rect 76701 72206 76765 72210
rect 77789 72746 77853 72750
rect 77789 72690 77793 72746
rect 77793 72690 77849 72746
rect 77849 72690 77853 72746
rect 77789 72686 77853 72690
rect 77789 72666 77853 72670
rect 77789 72610 77793 72666
rect 77793 72610 77849 72666
rect 77849 72610 77853 72666
rect 77789 72606 77853 72610
rect 77789 72586 77853 72590
rect 77789 72530 77793 72586
rect 77793 72530 77849 72586
rect 77849 72530 77853 72586
rect 77789 72526 77853 72530
rect 77789 72506 77853 72510
rect 77789 72450 77793 72506
rect 77793 72450 77849 72506
rect 77849 72450 77853 72506
rect 77789 72446 77853 72450
rect 77789 72426 77853 72430
rect 77789 72370 77793 72426
rect 77793 72370 77849 72426
rect 77849 72370 77853 72426
rect 77789 72366 77853 72370
rect 77789 72346 77853 72350
rect 77789 72290 77793 72346
rect 77793 72290 77849 72346
rect 77849 72290 77853 72346
rect 77789 72286 77853 72290
rect 77789 72266 77853 72270
rect 77789 72210 77793 72266
rect 77793 72210 77849 72266
rect 77849 72210 77853 72266
rect 77789 72206 77853 72210
rect 78877 72746 78941 72750
rect 78877 72690 78881 72746
rect 78881 72690 78937 72746
rect 78937 72690 78941 72746
rect 78877 72686 78941 72690
rect 78877 72666 78941 72670
rect 78877 72610 78881 72666
rect 78881 72610 78937 72666
rect 78937 72610 78941 72666
rect 78877 72606 78941 72610
rect 78877 72586 78941 72590
rect 78877 72530 78881 72586
rect 78881 72530 78937 72586
rect 78937 72530 78941 72586
rect 78877 72526 78941 72530
rect 78877 72506 78941 72510
rect 78877 72450 78881 72506
rect 78881 72450 78937 72506
rect 78937 72450 78941 72506
rect 78877 72446 78941 72450
rect 78877 72426 78941 72430
rect 78877 72370 78881 72426
rect 78881 72370 78937 72426
rect 78937 72370 78941 72426
rect 78877 72366 78941 72370
rect 78877 72346 78941 72350
rect 78877 72290 78881 72346
rect 78881 72290 78937 72346
rect 78937 72290 78941 72346
rect 78877 72286 78941 72290
rect 78877 72266 78941 72270
rect 78877 72210 78881 72266
rect 78881 72210 78937 72266
rect 78937 72210 78941 72266
rect 78877 72206 78941 72210
rect 79965 72746 80029 72750
rect 79965 72690 79969 72746
rect 79969 72690 80025 72746
rect 80025 72690 80029 72746
rect 79965 72686 80029 72690
rect 79965 72666 80029 72670
rect 79965 72610 79969 72666
rect 79969 72610 80025 72666
rect 80025 72610 80029 72666
rect 79965 72606 80029 72610
rect 79965 72586 80029 72590
rect 79965 72530 79969 72586
rect 79969 72530 80025 72586
rect 80025 72530 80029 72586
rect 79965 72526 80029 72530
rect 79965 72506 80029 72510
rect 79965 72450 79969 72506
rect 79969 72450 80025 72506
rect 80025 72450 80029 72506
rect 79965 72446 80029 72450
rect 79965 72426 80029 72430
rect 79965 72370 79969 72426
rect 79969 72370 80025 72426
rect 80025 72370 80029 72426
rect 79965 72366 80029 72370
rect 79965 72346 80029 72350
rect 79965 72290 79969 72346
rect 79969 72290 80025 72346
rect 80025 72290 80029 72346
rect 79965 72286 80029 72290
rect 79965 72266 80029 72270
rect 79965 72210 79969 72266
rect 79969 72210 80025 72266
rect 80025 72210 80029 72266
rect 79965 72206 80029 72210
rect 81053 72746 81117 72750
rect 81053 72690 81057 72746
rect 81057 72690 81113 72746
rect 81113 72690 81117 72746
rect 81053 72686 81117 72690
rect 81053 72666 81117 72670
rect 81053 72610 81057 72666
rect 81057 72610 81113 72666
rect 81113 72610 81117 72666
rect 81053 72606 81117 72610
rect 81053 72586 81117 72590
rect 81053 72530 81057 72586
rect 81057 72530 81113 72586
rect 81113 72530 81117 72586
rect 81053 72526 81117 72530
rect 81053 72506 81117 72510
rect 81053 72450 81057 72506
rect 81057 72450 81113 72506
rect 81113 72450 81117 72506
rect 81053 72446 81117 72450
rect 81053 72426 81117 72430
rect 81053 72370 81057 72426
rect 81057 72370 81113 72426
rect 81113 72370 81117 72426
rect 81053 72366 81117 72370
rect 81053 72346 81117 72350
rect 81053 72290 81057 72346
rect 81057 72290 81113 72346
rect 81113 72290 81117 72346
rect 81053 72286 81117 72290
rect 81053 72266 81117 72270
rect 81053 72210 81057 72266
rect 81057 72210 81113 72266
rect 81113 72210 81117 72266
rect 81053 72206 81117 72210
rect 86493 72746 86557 72750
rect 86493 72690 86497 72746
rect 86497 72690 86553 72746
rect 86553 72690 86557 72746
rect 86493 72686 86557 72690
rect 86493 72666 86557 72670
rect 86493 72610 86497 72666
rect 86497 72610 86553 72666
rect 86553 72610 86557 72666
rect 86493 72606 86557 72610
rect 86493 72586 86557 72590
rect 86493 72530 86497 72586
rect 86497 72530 86553 72586
rect 86553 72530 86557 72586
rect 86493 72526 86557 72530
rect 86493 72506 86557 72510
rect 86493 72450 86497 72506
rect 86497 72450 86553 72506
rect 86553 72450 86557 72506
rect 86493 72446 86557 72450
rect 86493 72426 86557 72430
rect 86493 72370 86497 72426
rect 86497 72370 86553 72426
rect 86553 72370 86557 72426
rect 86493 72366 86557 72370
rect 86493 72346 86557 72350
rect 86493 72290 86497 72346
rect 86497 72290 86553 72346
rect 86553 72290 86557 72346
rect 86493 72286 86557 72290
rect 86493 72266 86557 72270
rect 86493 72210 86497 72266
rect 86497 72210 86553 72266
rect 86553 72210 86557 72266
rect 86493 72206 86557 72210
rect 87581 72746 87645 72750
rect 87581 72690 87585 72746
rect 87585 72690 87641 72746
rect 87641 72690 87645 72746
rect 87581 72686 87645 72690
rect 87581 72666 87645 72670
rect 87581 72610 87585 72666
rect 87585 72610 87641 72666
rect 87641 72610 87645 72666
rect 87581 72606 87645 72610
rect 87581 72586 87645 72590
rect 87581 72530 87585 72586
rect 87585 72530 87641 72586
rect 87641 72530 87645 72586
rect 87581 72526 87645 72530
rect 87581 72506 87645 72510
rect 87581 72450 87585 72506
rect 87585 72450 87641 72506
rect 87641 72450 87645 72506
rect 87581 72446 87645 72450
rect 87581 72426 87645 72430
rect 87581 72370 87585 72426
rect 87585 72370 87641 72426
rect 87641 72370 87645 72426
rect 87581 72366 87645 72370
rect 87581 72346 87645 72350
rect 87581 72290 87585 72346
rect 87585 72290 87641 72346
rect 87641 72290 87645 72346
rect 87581 72286 87645 72290
rect 87581 72266 87645 72270
rect 87581 72210 87585 72266
rect 87585 72210 87641 72266
rect 87641 72210 87645 72266
rect 87581 72206 87645 72210
rect 88669 72746 88733 72750
rect 88669 72690 88673 72746
rect 88673 72690 88729 72746
rect 88729 72690 88733 72746
rect 88669 72686 88733 72690
rect 88669 72666 88733 72670
rect 88669 72610 88673 72666
rect 88673 72610 88729 72666
rect 88729 72610 88733 72666
rect 88669 72606 88733 72610
rect 88669 72586 88733 72590
rect 88669 72530 88673 72586
rect 88673 72530 88729 72586
rect 88729 72530 88733 72586
rect 88669 72526 88733 72530
rect 88669 72506 88733 72510
rect 88669 72450 88673 72506
rect 88673 72450 88729 72506
rect 88729 72450 88733 72506
rect 88669 72446 88733 72450
rect 88669 72426 88733 72430
rect 88669 72370 88673 72426
rect 88673 72370 88729 72426
rect 88729 72370 88733 72426
rect 88669 72366 88733 72370
rect 88669 72346 88733 72350
rect 88669 72290 88673 72346
rect 88673 72290 88729 72346
rect 88729 72290 88733 72346
rect 88669 72286 88733 72290
rect 88669 72266 88733 72270
rect 88669 72210 88673 72266
rect 88673 72210 88729 72266
rect 88729 72210 88733 72266
rect 88669 72206 88733 72210
rect 45733 71214 45797 71278
rect 50683 71214 50747 71278
rect 30023 67296 30087 67300
rect 30023 67240 30027 67296
rect 30027 67240 30083 67296
rect 30083 67240 30087 67296
rect 30023 67236 30087 67240
rect 30023 67216 30087 67220
rect 30023 67160 30027 67216
rect 30027 67160 30083 67216
rect 30083 67160 30087 67216
rect 30023 67156 30087 67160
rect 30023 67136 30087 67140
rect 30023 67080 30027 67136
rect 30027 67080 30083 67136
rect 30083 67080 30087 67136
rect 30023 67076 30087 67080
rect 30023 67056 30087 67060
rect 30023 67000 30027 67056
rect 30027 67000 30083 67056
rect 30083 67000 30087 67056
rect 30023 66996 30087 67000
rect 30023 66976 30087 66980
rect 30023 66920 30027 66976
rect 30027 66920 30083 66976
rect 30083 66920 30087 66976
rect 30023 66916 30087 66920
rect 30023 66896 30087 66900
rect 30023 66840 30027 66896
rect 30027 66840 30083 66896
rect 30083 66840 30087 66896
rect 30023 66836 30087 66840
rect 30023 66155 30087 66159
rect 30023 66099 30027 66155
rect 30027 66099 30083 66155
rect 30083 66099 30087 66155
rect 30023 66095 30087 66099
rect 30023 66075 30087 66079
rect 30023 66019 30027 66075
rect 30027 66019 30083 66075
rect 30083 66019 30087 66075
rect 30023 66015 30087 66019
rect 30023 65995 30087 65999
rect 30023 65939 30027 65995
rect 30027 65939 30083 65995
rect 30083 65939 30087 65995
rect 30023 65935 30087 65939
rect 30023 65915 30087 65919
rect 30023 65859 30027 65915
rect 30027 65859 30083 65915
rect 30083 65859 30087 65915
rect 30023 65855 30087 65859
rect 30023 65835 30087 65839
rect 30023 65779 30027 65835
rect 30027 65779 30083 65835
rect 30083 65779 30087 65835
rect 30023 65775 30087 65779
rect 30023 65755 30087 65759
rect 30023 65699 30027 65755
rect 30027 65699 30083 65755
rect 30083 65699 30087 65755
rect 30023 65695 30087 65699
rect 30023 65675 30087 65679
rect 30023 65619 30027 65675
rect 30027 65619 30083 65675
rect 30083 65619 30087 65675
rect 30023 65615 30087 65619
rect 30023 65595 30087 65599
rect 30023 65539 30027 65595
rect 30027 65539 30083 65595
rect 30083 65539 30087 65595
rect 30023 65535 30087 65539
rect 30023 65515 30087 65519
rect 30023 65459 30027 65515
rect 30027 65459 30083 65515
rect 30083 65459 30087 65515
rect 30023 65455 30087 65459
rect 30023 65435 30087 65439
rect 30023 65379 30027 65435
rect 30027 65379 30083 65435
rect 30083 65379 30087 65435
rect 30023 65375 30087 65379
rect 30023 65355 30087 65359
rect 30023 65299 30027 65355
rect 30027 65299 30083 65355
rect 30083 65299 30087 65355
rect 30023 65295 30087 65299
rect 30023 65275 30087 65279
rect 30023 65219 30027 65275
rect 30027 65219 30083 65275
rect 30083 65219 30087 65275
rect 30023 65215 30087 65219
rect 30023 65195 30087 65199
rect 30023 65139 30027 65195
rect 30027 65139 30083 65195
rect 30083 65139 30087 65195
rect 30023 65135 30087 65139
rect 30023 65115 30087 65119
rect 30023 65059 30027 65115
rect 30027 65059 30083 65115
rect 30083 65059 30087 65115
rect 30023 65055 30087 65059
rect 30028 64629 30092 64633
rect 30028 64573 30032 64629
rect 30032 64573 30088 64629
rect 30088 64573 30092 64629
rect 30028 64569 30092 64573
rect 30028 64549 30092 64553
rect 30028 64493 30032 64549
rect 30032 64493 30088 64549
rect 30088 64493 30092 64549
rect 30028 64489 30092 64493
rect 30028 64469 30092 64473
rect 30028 64413 30032 64469
rect 30032 64413 30088 64469
rect 30088 64413 30092 64469
rect 30028 64409 30092 64413
rect 30028 64389 30092 64393
rect 30028 64333 30032 64389
rect 30032 64333 30088 64389
rect 30088 64333 30092 64389
rect 30028 64329 30092 64333
rect 30028 64309 30092 64313
rect 30028 64253 30032 64309
rect 30032 64253 30088 64309
rect 30088 64253 30092 64309
rect 30028 64249 30092 64253
rect 30028 64229 30092 64233
rect 30028 64173 30032 64229
rect 30032 64173 30088 64229
rect 30088 64173 30092 64229
rect 30028 64169 30092 64173
rect 30028 64149 30092 64153
rect 30028 64093 30032 64149
rect 30032 64093 30088 64149
rect 30088 64093 30092 64149
rect 30028 64089 30092 64093
rect 30028 64069 30092 64073
rect 30028 64013 30032 64069
rect 30032 64013 30088 64069
rect 30088 64013 30092 64069
rect 30028 64009 30092 64013
rect 30028 63989 30092 63993
rect 30028 63933 30032 63989
rect 30032 63933 30088 63989
rect 30088 63933 30092 63989
rect 30028 63929 30092 63933
rect 30028 63909 30092 63913
rect 30028 63853 30032 63909
rect 30032 63853 30088 63909
rect 30088 63853 30092 63909
rect 30028 63849 30092 63853
rect 30028 63829 30092 63833
rect 30028 63773 30032 63829
rect 30032 63773 30088 63829
rect 30088 63773 30092 63829
rect 30028 63769 30092 63773
rect 30028 63749 30092 63753
rect 30028 63693 30032 63749
rect 30032 63693 30088 63749
rect 30088 63693 30092 63749
rect 30028 63689 30092 63693
rect 30028 63669 30092 63673
rect 30028 63613 30032 63669
rect 30032 63613 30088 63669
rect 30088 63613 30092 63669
rect 30028 63609 30092 63613
rect 30028 63589 30092 63593
rect 30028 63533 30032 63589
rect 30032 63533 30088 63589
rect 30088 63533 30092 63589
rect 30028 63529 30092 63533
rect 25282 63166 25346 63170
rect 25282 63110 25286 63166
rect 25286 63110 25342 63166
rect 25342 63110 25346 63166
rect 25282 63106 25346 63110
rect 25282 63086 25346 63090
rect 25282 63030 25286 63086
rect 25286 63030 25342 63086
rect 25342 63030 25346 63086
rect 25282 63026 25346 63030
rect 25282 63006 25346 63010
rect 25282 62950 25286 63006
rect 25286 62950 25342 63006
rect 25342 62950 25346 63006
rect 25282 62946 25346 62950
rect 25282 62926 25346 62930
rect 25282 62870 25286 62926
rect 25286 62870 25342 62926
rect 25342 62870 25346 62926
rect 25282 62866 25346 62870
rect 30022 63126 30086 63130
rect 30022 63070 30026 63126
rect 30026 63070 30082 63126
rect 30082 63070 30086 63126
rect 30022 63066 30086 63070
rect 30022 63046 30086 63050
rect 30022 62990 30026 63046
rect 30026 62990 30082 63046
rect 30082 62990 30086 63046
rect 30022 62986 30086 62990
rect 30022 62966 30086 62970
rect 30022 62910 30026 62966
rect 30026 62910 30082 62966
rect 30082 62910 30086 62966
rect 30022 62906 30086 62910
rect 30022 62886 30086 62890
rect 30022 62830 30026 62886
rect 30026 62830 30082 62886
rect 30082 62830 30086 62886
rect 30022 62826 30086 62830
rect 30022 62806 30086 62810
rect 30022 62750 30026 62806
rect 30026 62750 30082 62806
rect 30082 62750 30086 62806
rect 30022 62746 30086 62750
rect 30022 62726 30086 62730
rect 30022 62670 30026 62726
rect 30026 62670 30082 62726
rect 30082 62670 30086 62726
rect 30022 62666 30086 62670
rect 25283 62627 25347 62631
rect 25283 62571 25287 62627
rect 25287 62571 25343 62627
rect 25343 62571 25347 62627
rect 25283 62567 25347 62571
rect 25283 62547 25347 62551
rect 25283 62491 25287 62547
rect 25287 62491 25343 62547
rect 25343 62491 25347 62547
rect 25283 62487 25347 62491
rect 25283 62467 25347 62471
rect 25283 62411 25287 62467
rect 25287 62411 25343 62467
rect 25343 62411 25347 62467
rect 25283 62407 25347 62411
rect 30022 62646 30086 62650
rect 30022 62590 30026 62646
rect 30026 62590 30082 62646
rect 30082 62590 30086 62646
rect 30022 62586 30086 62590
rect 30022 62566 30086 62570
rect 30022 62510 30026 62566
rect 30026 62510 30082 62566
rect 30082 62510 30086 62566
rect 30022 62506 30086 62510
rect 25283 62387 25347 62391
rect 25283 62331 25287 62387
rect 25287 62331 25343 62387
rect 25343 62331 25347 62387
rect 25283 62327 25347 62331
rect 27480 62431 27544 62435
rect 27480 62375 27484 62431
rect 27484 62375 27540 62431
rect 27540 62375 27544 62431
rect 27480 62371 27544 62375
rect 27560 62431 27624 62435
rect 27560 62375 27564 62431
rect 27564 62375 27620 62431
rect 27620 62375 27624 62431
rect 27560 62371 27624 62375
rect 27640 62431 27704 62435
rect 27640 62375 27644 62431
rect 27644 62375 27700 62431
rect 27700 62375 27704 62431
rect 27640 62371 27704 62375
rect 27720 62431 27784 62435
rect 27720 62375 27724 62431
rect 27724 62375 27780 62431
rect 27780 62375 27784 62431
rect 27720 62371 27784 62375
rect 27800 62431 27864 62435
rect 27800 62375 27804 62431
rect 27804 62375 27860 62431
rect 27860 62375 27864 62431
rect 27800 62371 27864 62375
rect 27880 62431 27944 62435
rect 27880 62375 27884 62431
rect 27884 62375 27940 62431
rect 27940 62375 27944 62431
rect 27880 62371 27944 62375
rect 30022 62486 30086 62490
rect 30022 62430 30026 62486
rect 30026 62430 30082 62486
rect 30082 62430 30086 62486
rect 30022 62426 30086 62430
rect 25283 62307 25347 62311
rect 25283 62251 25287 62307
rect 25287 62251 25343 62307
rect 25343 62251 25347 62307
rect 25283 62247 25347 62251
rect 30022 62406 30086 62410
rect 30022 62350 30026 62406
rect 30026 62350 30082 62406
rect 30082 62350 30086 62406
rect 30022 62346 30086 62350
rect 30022 62326 30086 62330
rect 30022 62270 30026 62326
rect 30026 62270 30082 62326
rect 30082 62270 30086 62326
rect 30022 62266 30086 62270
rect 25283 62227 25347 62231
rect 25283 62171 25287 62227
rect 25287 62171 25343 62227
rect 25343 62171 25347 62227
rect 25283 62167 25347 62171
rect 75070 70743 75134 70747
rect 75070 70687 75074 70743
rect 75074 70687 75130 70743
rect 75130 70687 75134 70743
rect 75070 70683 75134 70687
rect 46607 70591 46671 70655
rect 50683 70591 50747 70655
rect 75070 70663 75134 70667
rect 75070 70607 75074 70663
rect 75074 70607 75130 70663
rect 75130 70607 75134 70663
rect 75070 70603 75134 70607
rect 75070 70583 75134 70587
rect 75070 70527 75074 70583
rect 75074 70527 75130 70583
rect 75130 70527 75134 70583
rect 75070 70523 75134 70527
rect 75070 70503 75134 70507
rect 75070 70447 75074 70503
rect 75074 70447 75130 70503
rect 75130 70447 75134 70503
rect 75070 70443 75134 70447
rect 75070 70423 75134 70427
rect 75070 70367 75074 70423
rect 75074 70367 75130 70423
rect 75130 70367 75134 70423
rect 75070 70363 75134 70367
rect 43625 67079 43689 67083
rect 43625 67023 43629 67079
rect 43629 67023 43685 67079
rect 43685 67023 43689 67079
rect 43625 67019 43689 67023
rect 47886 67019 47950 67083
rect 44401 66416 44465 66420
rect 44401 66360 44405 66416
rect 44405 66360 44461 66416
rect 44461 66360 44465 66416
rect 44401 66356 44465 66360
rect 47025 66356 47089 66420
rect 35619 66181 35683 66185
rect 35619 66125 35623 66181
rect 35623 66125 35679 66181
rect 35679 66125 35683 66181
rect 35619 66121 35683 66125
rect 51199 70256 51343 70260
rect 51199 63880 51203 70256
rect 51203 63880 51339 70256
rect 51339 63880 51343 70256
rect 75070 70343 75134 70347
rect 75070 70287 75074 70343
rect 75074 70287 75130 70343
rect 75130 70287 75134 70343
rect 75070 70283 75134 70287
rect 75070 70263 75134 70267
rect 75070 70207 75074 70263
rect 75074 70207 75130 70263
rect 75130 70207 75134 70263
rect 75070 70203 75134 70207
rect 76158 70743 76222 70747
rect 76158 70687 76162 70743
rect 76162 70687 76218 70743
rect 76218 70687 76222 70743
rect 76158 70683 76222 70687
rect 76158 70663 76222 70667
rect 76158 70607 76162 70663
rect 76162 70607 76218 70663
rect 76218 70607 76222 70663
rect 76158 70603 76222 70607
rect 76158 70583 76222 70587
rect 76158 70527 76162 70583
rect 76162 70527 76218 70583
rect 76218 70527 76222 70583
rect 76158 70523 76222 70527
rect 76158 70503 76222 70507
rect 76158 70447 76162 70503
rect 76162 70447 76218 70503
rect 76218 70447 76222 70503
rect 76158 70443 76222 70447
rect 76158 70423 76222 70427
rect 76158 70367 76162 70423
rect 76162 70367 76218 70423
rect 76218 70367 76222 70423
rect 76158 70363 76222 70367
rect 76158 70343 76222 70347
rect 76158 70287 76162 70343
rect 76162 70287 76218 70343
rect 76218 70287 76222 70343
rect 76158 70283 76222 70287
rect 76158 70263 76222 70267
rect 76158 70207 76162 70263
rect 76162 70207 76218 70263
rect 76218 70207 76222 70263
rect 76158 70203 76222 70207
rect 77246 70743 77310 70747
rect 77246 70687 77250 70743
rect 77250 70687 77306 70743
rect 77306 70687 77310 70743
rect 77246 70683 77310 70687
rect 77246 70663 77310 70667
rect 77246 70607 77250 70663
rect 77250 70607 77306 70663
rect 77306 70607 77310 70663
rect 77246 70603 77310 70607
rect 77246 70583 77310 70587
rect 77246 70527 77250 70583
rect 77250 70527 77306 70583
rect 77306 70527 77310 70583
rect 77246 70523 77310 70527
rect 77246 70503 77310 70507
rect 77246 70447 77250 70503
rect 77250 70447 77306 70503
rect 77306 70447 77310 70503
rect 77246 70443 77310 70447
rect 77246 70423 77310 70427
rect 77246 70367 77250 70423
rect 77250 70367 77306 70423
rect 77306 70367 77310 70423
rect 77246 70363 77310 70367
rect 77246 70343 77310 70347
rect 77246 70287 77250 70343
rect 77250 70287 77306 70343
rect 77306 70287 77310 70343
rect 77246 70283 77310 70287
rect 77246 70263 77310 70267
rect 77246 70207 77250 70263
rect 77250 70207 77306 70263
rect 77306 70207 77310 70263
rect 77246 70203 77310 70207
rect 78334 70743 78398 70747
rect 78334 70687 78338 70743
rect 78338 70687 78394 70743
rect 78394 70687 78398 70743
rect 78334 70683 78398 70687
rect 78334 70663 78398 70667
rect 78334 70607 78338 70663
rect 78338 70607 78394 70663
rect 78394 70607 78398 70663
rect 78334 70603 78398 70607
rect 78334 70583 78398 70587
rect 78334 70527 78338 70583
rect 78338 70527 78394 70583
rect 78394 70527 78398 70583
rect 78334 70523 78398 70527
rect 78334 70503 78398 70507
rect 78334 70447 78338 70503
rect 78338 70447 78394 70503
rect 78394 70447 78398 70503
rect 78334 70443 78398 70447
rect 78334 70423 78398 70427
rect 78334 70367 78338 70423
rect 78338 70367 78394 70423
rect 78394 70367 78398 70423
rect 78334 70363 78398 70367
rect 78334 70343 78398 70347
rect 78334 70287 78338 70343
rect 78338 70287 78394 70343
rect 78394 70287 78398 70343
rect 78334 70283 78398 70287
rect 78334 70263 78398 70267
rect 78334 70207 78338 70263
rect 78338 70207 78394 70263
rect 78394 70207 78398 70263
rect 78334 70203 78398 70207
rect 79422 70743 79486 70747
rect 79422 70687 79426 70743
rect 79426 70687 79482 70743
rect 79482 70687 79486 70743
rect 79422 70683 79486 70687
rect 79422 70663 79486 70667
rect 79422 70607 79426 70663
rect 79426 70607 79482 70663
rect 79482 70607 79486 70663
rect 79422 70603 79486 70607
rect 79422 70583 79486 70587
rect 79422 70527 79426 70583
rect 79426 70527 79482 70583
rect 79482 70527 79486 70583
rect 79422 70523 79486 70527
rect 79422 70503 79486 70507
rect 79422 70447 79426 70503
rect 79426 70447 79482 70503
rect 79482 70447 79486 70503
rect 79422 70443 79486 70447
rect 79422 70423 79486 70427
rect 79422 70367 79426 70423
rect 79426 70367 79482 70423
rect 79482 70367 79486 70423
rect 79422 70363 79486 70367
rect 79422 70343 79486 70347
rect 79422 70287 79426 70343
rect 79426 70287 79482 70343
rect 79482 70287 79486 70343
rect 79422 70283 79486 70287
rect 79422 70263 79486 70267
rect 79422 70207 79426 70263
rect 79426 70207 79482 70263
rect 79482 70207 79486 70263
rect 79422 70203 79486 70207
rect 81598 70743 81662 70747
rect 81598 70687 81602 70743
rect 81602 70687 81658 70743
rect 81658 70687 81662 70743
rect 81598 70683 81662 70687
rect 81598 70663 81662 70667
rect 81598 70607 81602 70663
rect 81602 70607 81658 70663
rect 81658 70607 81662 70663
rect 81598 70603 81662 70607
rect 81598 70583 81662 70587
rect 81598 70527 81602 70583
rect 81602 70527 81658 70583
rect 81658 70527 81662 70583
rect 81598 70523 81662 70527
rect 81598 70503 81662 70507
rect 81598 70447 81602 70503
rect 81602 70447 81658 70503
rect 81658 70447 81662 70503
rect 81598 70443 81662 70447
rect 81598 70423 81662 70427
rect 81598 70367 81602 70423
rect 81602 70367 81658 70423
rect 81658 70367 81662 70423
rect 81598 70363 81662 70367
rect 81598 70343 81662 70347
rect 81598 70287 81602 70343
rect 81602 70287 81658 70343
rect 81658 70287 81662 70343
rect 81598 70283 81662 70287
rect 81598 70263 81662 70267
rect 81598 70207 81602 70263
rect 81602 70207 81658 70263
rect 81658 70207 81662 70263
rect 81598 70203 81662 70207
rect 82686 70743 82750 70747
rect 82686 70687 82690 70743
rect 82690 70687 82746 70743
rect 82746 70687 82750 70743
rect 82686 70683 82750 70687
rect 82686 70663 82750 70667
rect 82686 70607 82690 70663
rect 82690 70607 82746 70663
rect 82746 70607 82750 70663
rect 82686 70603 82750 70607
rect 82686 70583 82750 70587
rect 82686 70527 82690 70583
rect 82690 70527 82746 70583
rect 82746 70527 82750 70583
rect 82686 70523 82750 70527
rect 82686 70503 82750 70507
rect 82686 70447 82690 70503
rect 82690 70447 82746 70503
rect 82746 70447 82750 70503
rect 82686 70443 82750 70447
rect 82686 70423 82750 70427
rect 82686 70367 82690 70423
rect 82690 70367 82746 70423
rect 82746 70367 82750 70423
rect 82686 70363 82750 70367
rect 82686 70343 82750 70347
rect 82686 70287 82690 70343
rect 82690 70287 82746 70343
rect 82746 70287 82750 70343
rect 82686 70283 82750 70287
rect 82686 70263 82750 70267
rect 82686 70207 82690 70263
rect 82690 70207 82746 70263
rect 82746 70207 82750 70263
rect 82686 70203 82750 70207
rect 83774 70743 83838 70747
rect 83774 70687 83778 70743
rect 83778 70687 83834 70743
rect 83834 70687 83838 70743
rect 83774 70683 83838 70687
rect 83774 70663 83838 70667
rect 83774 70607 83778 70663
rect 83778 70607 83834 70663
rect 83834 70607 83838 70663
rect 83774 70603 83838 70607
rect 83774 70583 83838 70587
rect 83774 70527 83778 70583
rect 83778 70527 83834 70583
rect 83834 70527 83838 70583
rect 83774 70523 83838 70527
rect 83774 70503 83838 70507
rect 83774 70447 83778 70503
rect 83778 70447 83834 70503
rect 83834 70447 83838 70503
rect 83774 70443 83838 70447
rect 83774 70423 83838 70427
rect 83774 70367 83778 70423
rect 83778 70367 83834 70423
rect 83834 70367 83838 70423
rect 83774 70363 83838 70367
rect 83774 70343 83838 70347
rect 83774 70287 83778 70343
rect 83778 70287 83834 70343
rect 83834 70287 83838 70343
rect 83774 70283 83838 70287
rect 83774 70263 83838 70267
rect 83774 70207 83778 70263
rect 83778 70207 83834 70263
rect 83834 70207 83838 70263
rect 83774 70203 83838 70207
rect 84862 70743 84926 70747
rect 84862 70687 84866 70743
rect 84866 70687 84922 70743
rect 84922 70687 84926 70743
rect 84862 70683 84926 70687
rect 84862 70663 84926 70667
rect 84862 70607 84866 70663
rect 84866 70607 84922 70663
rect 84922 70607 84926 70663
rect 84862 70603 84926 70607
rect 84862 70583 84926 70587
rect 84862 70527 84866 70583
rect 84866 70527 84922 70583
rect 84922 70527 84926 70583
rect 84862 70523 84926 70527
rect 84862 70503 84926 70507
rect 84862 70447 84866 70503
rect 84866 70447 84922 70503
rect 84922 70447 84926 70503
rect 84862 70443 84926 70447
rect 84862 70423 84926 70427
rect 84862 70367 84866 70423
rect 84866 70367 84922 70423
rect 84922 70367 84926 70423
rect 84862 70363 84926 70367
rect 84862 70343 84926 70347
rect 84862 70287 84866 70343
rect 84866 70287 84922 70343
rect 84922 70287 84926 70343
rect 84862 70283 84926 70287
rect 84862 70263 84926 70267
rect 84862 70207 84866 70263
rect 84866 70207 84922 70263
rect 84922 70207 84926 70263
rect 84862 70203 84926 70207
rect 85950 70743 86014 70747
rect 85950 70687 85954 70743
rect 85954 70687 86010 70743
rect 86010 70687 86014 70743
rect 85950 70683 86014 70687
rect 85950 70663 86014 70667
rect 85950 70607 85954 70663
rect 85954 70607 86010 70663
rect 86010 70607 86014 70663
rect 85950 70603 86014 70607
rect 85950 70583 86014 70587
rect 85950 70527 85954 70583
rect 85954 70527 86010 70583
rect 86010 70527 86014 70583
rect 85950 70523 86014 70527
rect 85950 70503 86014 70507
rect 85950 70447 85954 70503
rect 85954 70447 86010 70503
rect 86010 70447 86014 70503
rect 85950 70443 86014 70447
rect 85950 70423 86014 70427
rect 85950 70367 85954 70423
rect 85954 70367 86010 70423
rect 86010 70367 86014 70423
rect 85950 70363 86014 70367
rect 85950 70343 86014 70347
rect 85950 70287 85954 70343
rect 85954 70287 86010 70343
rect 86010 70287 86014 70343
rect 85950 70283 86014 70287
rect 85950 70263 86014 70267
rect 85950 70207 85954 70263
rect 85954 70207 86010 70263
rect 86010 70207 86014 70263
rect 85950 70203 86014 70207
rect 87038 70743 87102 70747
rect 87038 70687 87042 70743
rect 87042 70687 87098 70743
rect 87098 70687 87102 70743
rect 87038 70683 87102 70687
rect 87038 70663 87102 70667
rect 87038 70607 87042 70663
rect 87042 70607 87098 70663
rect 87098 70607 87102 70663
rect 87038 70603 87102 70607
rect 87038 70583 87102 70587
rect 87038 70527 87042 70583
rect 87042 70527 87098 70583
rect 87098 70527 87102 70583
rect 87038 70523 87102 70527
rect 87038 70503 87102 70507
rect 87038 70447 87042 70503
rect 87042 70447 87098 70503
rect 87098 70447 87102 70503
rect 87038 70443 87102 70447
rect 87038 70423 87102 70427
rect 87038 70367 87042 70423
rect 87042 70367 87098 70423
rect 87098 70367 87102 70423
rect 87038 70363 87102 70367
rect 87038 70343 87102 70347
rect 87038 70287 87042 70343
rect 87042 70287 87098 70343
rect 87098 70287 87102 70343
rect 87038 70283 87102 70287
rect 87038 70263 87102 70267
rect 87038 70207 87042 70263
rect 87042 70207 87098 70263
rect 87098 70207 87102 70263
rect 87038 70203 87102 70207
rect 88126 70743 88190 70747
rect 88126 70687 88130 70743
rect 88130 70687 88186 70743
rect 88186 70687 88190 70743
rect 88126 70683 88190 70687
rect 88126 70663 88190 70667
rect 88126 70607 88130 70663
rect 88130 70607 88186 70663
rect 88186 70607 88190 70663
rect 88126 70603 88190 70607
rect 88126 70583 88190 70587
rect 88126 70527 88130 70583
rect 88130 70527 88186 70583
rect 88186 70527 88190 70583
rect 88126 70523 88190 70527
rect 88126 70503 88190 70507
rect 88126 70447 88130 70503
rect 88130 70447 88186 70503
rect 88186 70447 88190 70503
rect 88126 70443 88190 70447
rect 88126 70423 88190 70427
rect 88126 70367 88130 70423
rect 88130 70367 88186 70423
rect 88186 70367 88190 70423
rect 88126 70363 88190 70367
rect 88126 70343 88190 70347
rect 88126 70287 88130 70343
rect 88130 70287 88186 70343
rect 88186 70287 88190 70343
rect 88126 70283 88190 70287
rect 88126 70263 88190 70267
rect 88126 70207 88130 70263
rect 88130 70207 88186 70263
rect 88186 70207 88190 70263
rect 88126 70203 88190 70207
rect 57473 69851 57617 69855
rect 57473 68355 57477 69851
rect 57477 68355 57613 69851
rect 57613 68355 57617 69851
rect 57473 68351 57617 68355
rect 51199 63876 51343 63880
rect 57454 65389 57598 65393
rect 57454 63893 57458 65389
rect 57458 63893 57594 65389
rect 57594 63893 57598 65389
rect 57454 63889 57598 63893
rect 67307 70127 67611 70131
rect 67307 63911 67311 70127
rect 67311 63911 67607 70127
rect 67607 63911 67611 70127
rect 67307 63907 67611 63911
rect 75339 69766 75403 69770
rect 75339 69710 75343 69766
rect 75343 69710 75399 69766
rect 75399 69710 75403 69766
rect 75339 69706 75403 69710
rect 75885 69766 75949 69770
rect 75885 69710 75889 69766
rect 75889 69710 75945 69766
rect 75945 69710 75949 69766
rect 75885 69706 75949 69710
rect 76431 69757 76495 69761
rect 76431 69701 76435 69757
rect 76435 69701 76491 69757
rect 76491 69701 76495 69757
rect 76431 69697 76495 69701
rect 76976 69756 77040 69760
rect 76976 69700 76980 69756
rect 76980 69700 77036 69756
rect 77036 69700 77040 69756
rect 76976 69696 77040 69700
rect 78607 69744 78671 69748
rect 78607 69688 78611 69744
rect 78611 69688 78667 69744
rect 78667 69688 78671 69744
rect 78607 69684 78671 69688
rect 79150 69741 79214 69745
rect 79150 69685 79154 69741
rect 79154 69685 79210 69741
rect 79210 69685 79214 69741
rect 79150 69681 79214 69685
rect 79692 69740 79756 69744
rect 79692 69684 79696 69740
rect 79696 69684 79752 69740
rect 79752 69684 79756 69740
rect 79692 69680 79756 69684
rect 80239 69745 80303 69749
rect 80239 69689 80243 69745
rect 80243 69689 80299 69745
rect 80299 69689 80303 69745
rect 80239 69685 80303 69689
rect 82957 69756 83021 69760
rect 82957 69700 82961 69756
rect 82961 69700 83017 69756
rect 83017 69700 83021 69756
rect 82957 69696 83021 69700
rect 83500 69760 83564 69764
rect 83500 69704 83504 69760
rect 83504 69704 83560 69760
rect 83560 69704 83564 69760
rect 83500 69700 83564 69704
rect 84042 69754 84106 69758
rect 84042 69698 84046 69754
rect 84046 69698 84102 69754
rect 84102 69698 84106 69754
rect 84042 69694 84106 69698
rect 84599 69745 84663 69749
rect 84599 69689 84603 69745
rect 84603 69689 84659 69745
rect 84659 69689 84663 69745
rect 84599 69685 84663 69689
rect 86223 69756 86287 69760
rect 86223 69700 86227 69756
rect 86227 69700 86283 69756
rect 86283 69700 86287 69756
rect 86223 69696 86287 69700
rect 86767 69749 86831 69753
rect 86767 69693 86771 69749
rect 86771 69693 86827 69749
rect 86827 69693 86831 69749
rect 86767 69689 86831 69693
rect 87317 69753 87381 69757
rect 87317 69697 87321 69753
rect 87321 69697 87377 69753
rect 87377 69697 87381 69753
rect 87317 69693 87381 69697
rect 87850 69753 87914 69757
rect 87850 69697 87854 69753
rect 87854 69697 87910 69753
rect 87910 69697 87914 69753
rect 87850 69693 87914 69697
rect 75885 69030 75949 69094
rect 101852 69090 101916 69094
rect 101852 69034 101856 69090
rect 101856 69034 101912 69090
rect 101912 69034 101916 69090
rect 101852 69030 101916 69034
rect 101932 69090 101996 69094
rect 101932 69034 101936 69090
rect 101936 69034 101992 69090
rect 101992 69034 101996 69090
rect 101932 69030 101996 69034
rect 102012 69090 102076 69094
rect 102012 69034 102016 69090
rect 102016 69034 102072 69090
rect 102072 69034 102076 69090
rect 102012 69030 102076 69034
rect 102092 69090 102156 69094
rect 102092 69034 102096 69090
rect 102096 69034 102152 69090
rect 102152 69034 102156 69090
rect 102092 69030 102156 69034
rect 102172 69090 102236 69094
rect 102172 69034 102176 69090
rect 102176 69034 102232 69090
rect 102232 69034 102236 69090
rect 102172 69030 102236 69034
rect 102252 69090 102316 69094
rect 102252 69034 102256 69090
rect 102256 69034 102312 69090
rect 102312 69034 102316 69090
rect 102252 69030 102316 69034
rect 102332 69090 102396 69094
rect 102332 69034 102336 69090
rect 102336 69034 102392 69090
rect 102392 69034 102396 69090
rect 102332 69030 102396 69034
rect 82957 68849 83021 68913
rect 75339 68659 75403 68723
rect 83500 68484 83564 68548
rect 98637 68544 98701 68548
rect 98637 68488 98641 68544
rect 98641 68488 98697 68544
rect 98697 68488 98701 68544
rect 98637 68484 98701 68488
rect 98717 68544 98781 68548
rect 98717 68488 98721 68544
rect 98721 68488 98777 68544
rect 98777 68488 98781 68544
rect 98717 68484 98781 68488
rect 98797 68544 98861 68548
rect 98797 68488 98801 68544
rect 98801 68488 98857 68544
rect 98857 68488 98861 68544
rect 98797 68484 98861 68488
rect 98877 68544 98941 68548
rect 98877 68488 98881 68544
rect 98881 68488 98937 68544
rect 98937 68488 98941 68544
rect 98877 68484 98941 68488
rect 79691 67880 79755 67944
rect 101891 67939 101955 67943
rect 101891 67883 101895 67939
rect 101895 67883 101951 67939
rect 101951 67883 101955 67939
rect 101891 67879 101955 67883
rect 101971 67939 102035 67943
rect 101971 67883 101975 67939
rect 101975 67883 102031 67939
rect 102031 67883 102035 67939
rect 101971 67879 102035 67883
rect 102051 67939 102115 67943
rect 102051 67883 102055 67939
rect 102055 67883 102111 67939
rect 102111 67883 102115 67939
rect 102051 67879 102115 67883
rect 102131 67939 102195 67943
rect 102131 67883 102135 67939
rect 102135 67883 102191 67939
rect 102191 67883 102195 67939
rect 102131 67879 102195 67883
rect 102211 67939 102275 67943
rect 102211 67883 102215 67939
rect 102215 67883 102271 67939
rect 102271 67883 102275 67939
rect 102211 67879 102275 67883
rect 102291 67939 102355 67943
rect 102291 67883 102295 67939
rect 102295 67883 102351 67939
rect 102351 67883 102355 67939
rect 102291 67879 102355 67883
rect 87850 67699 87914 67763
rect 80239 67509 80303 67573
rect 87316 67333 87380 67397
rect 98635 67394 98699 67398
rect 98635 67338 98639 67394
rect 98639 67338 98695 67394
rect 98695 67338 98699 67394
rect 98635 67334 98699 67338
rect 98715 67394 98779 67398
rect 98715 67338 98719 67394
rect 98719 67338 98775 67394
rect 98775 67338 98779 67394
rect 98715 67334 98779 67338
rect 98795 67394 98859 67398
rect 98795 67338 98799 67394
rect 98799 67338 98855 67394
rect 98855 67338 98859 67394
rect 98795 67334 98859 67338
rect 98875 67394 98939 67398
rect 98875 67338 98879 67394
rect 98879 67338 98935 67394
rect 98935 67338 98939 67394
rect 98875 67334 98939 67338
rect 76976 65340 77040 65404
rect 101881 65397 101945 65401
rect 101881 65341 101885 65397
rect 101885 65341 101941 65397
rect 101941 65341 101945 65397
rect 101881 65337 101945 65341
rect 101961 65397 102025 65401
rect 101961 65341 101965 65397
rect 101965 65341 102021 65397
rect 102021 65341 102025 65397
rect 101961 65337 102025 65341
rect 102041 65397 102105 65401
rect 102041 65341 102045 65397
rect 102045 65341 102101 65397
rect 102101 65341 102105 65397
rect 102041 65337 102105 65341
rect 102121 65397 102185 65401
rect 102121 65341 102125 65397
rect 102125 65341 102181 65397
rect 102181 65341 102185 65397
rect 102121 65337 102185 65341
rect 102201 65397 102265 65401
rect 102201 65341 102205 65397
rect 102205 65341 102261 65397
rect 102261 65341 102265 65397
rect 102201 65337 102265 65341
rect 102281 65397 102345 65401
rect 102281 65341 102285 65397
rect 102285 65341 102341 65397
rect 102341 65341 102345 65397
rect 102281 65337 102345 65341
rect 84042 65159 84106 65223
rect 76431 64969 76495 65033
rect 84599 64794 84663 64858
rect 98553 64853 98617 64857
rect 98553 64797 98557 64853
rect 98557 64797 98613 64853
rect 98613 64797 98617 64853
rect 98553 64793 98617 64797
rect 98633 64853 98697 64857
rect 98633 64797 98637 64853
rect 98637 64797 98693 64853
rect 98693 64797 98697 64853
rect 98633 64793 98697 64797
rect 98713 64853 98777 64857
rect 98713 64797 98717 64853
rect 98717 64797 98773 64853
rect 98773 64797 98777 64853
rect 98713 64793 98777 64797
rect 98793 64853 98857 64857
rect 98793 64797 98797 64853
rect 98797 64797 98853 64853
rect 98853 64797 98857 64853
rect 98793 64793 98857 64797
rect 78607 64070 78671 64134
rect 101881 64127 101945 64131
rect 101881 64071 101885 64127
rect 101885 64071 101941 64127
rect 101941 64071 101945 64127
rect 101881 64067 101945 64071
rect 101961 64127 102025 64131
rect 101961 64071 101965 64127
rect 101965 64071 102021 64127
rect 102021 64071 102025 64127
rect 101961 64067 102025 64071
rect 102041 64127 102105 64131
rect 102041 64071 102045 64127
rect 102045 64071 102101 64127
rect 102101 64071 102105 64127
rect 102041 64067 102105 64071
rect 102121 64127 102185 64131
rect 102121 64071 102125 64127
rect 102125 64071 102181 64127
rect 102181 64071 102185 64127
rect 102121 64067 102185 64071
rect 102201 64127 102265 64131
rect 102201 64071 102205 64127
rect 102205 64071 102261 64127
rect 102261 64071 102265 64127
rect 102201 64067 102265 64071
rect 102281 64127 102345 64131
rect 102281 64071 102285 64127
rect 102285 64071 102341 64127
rect 102341 64071 102345 64127
rect 102281 64067 102345 64071
rect 86767 63889 86831 63953
rect 51426 63846 56930 63850
rect 51426 63710 51430 63846
rect 51430 63710 56926 63846
rect 56926 63710 56930 63846
rect 51426 63706 56930 63710
rect 79151 63699 79215 63763
rect 86223 63524 86287 63588
rect 98551 63584 98615 63588
rect 98551 63528 98555 63584
rect 98555 63528 98611 63584
rect 98611 63528 98615 63584
rect 98551 63524 98615 63528
rect 98631 63584 98695 63588
rect 98631 63528 98635 63584
rect 98635 63528 98691 63584
rect 98691 63528 98695 63584
rect 98631 63524 98695 63528
rect 98711 63584 98775 63588
rect 98711 63528 98715 63584
rect 98715 63528 98771 63584
rect 98771 63528 98775 63584
rect 98711 63524 98775 63528
rect 98791 63584 98855 63588
rect 98791 63528 98795 63584
rect 98795 63528 98851 63584
rect 98851 63528 98855 63584
rect 98791 63524 98855 63528
rect 38217 63520 38281 63524
rect 38217 63464 38221 63520
rect 38221 63464 38277 63520
rect 38277 63464 38281 63520
rect 38217 63460 38281 63464
rect 38217 63440 38281 63444
rect 38217 63384 38221 63440
rect 38221 63384 38277 63440
rect 38277 63384 38281 63440
rect 38217 63380 38281 63384
rect 38217 63360 38281 63364
rect 38217 63304 38221 63360
rect 38221 63304 38277 63360
rect 38277 63304 38281 63360
rect 38217 63300 38281 63304
rect 38217 63280 38281 63284
rect 38217 63224 38221 63280
rect 38221 63224 38277 63280
rect 38277 63224 38281 63280
rect 38217 63220 38281 63224
rect 38217 63200 38281 63204
rect 38217 63144 38221 63200
rect 38221 63144 38277 63200
rect 38277 63144 38281 63200
rect 38217 63140 38281 63144
rect 38217 63120 38281 63124
rect 38217 63064 38221 63120
rect 38221 63064 38277 63120
rect 38277 63064 38281 63120
rect 38217 63060 38281 63064
rect 38217 63040 38281 63044
rect 38217 62984 38221 63040
rect 38221 62984 38277 63040
rect 38277 62984 38281 63040
rect 38217 62980 38281 62984
rect 38217 62960 38281 62964
rect 38217 62904 38221 62960
rect 38221 62904 38277 62960
rect 38277 62904 38281 62960
rect 38217 62900 38281 62904
rect 38217 62880 38281 62884
rect 38217 62824 38221 62880
rect 38221 62824 38277 62880
rect 38277 62824 38281 62880
rect 38217 62820 38281 62824
rect 59616 62891 59680 62895
rect 59616 62835 59620 62891
rect 59620 62835 59676 62891
rect 59676 62835 59680 62891
rect 59616 62831 59680 62835
rect 38217 62800 38281 62804
rect 38217 62744 38221 62800
rect 38221 62744 38277 62800
rect 38277 62744 38281 62800
rect 38217 62740 38281 62744
rect 45381 62748 45445 62812
rect 52381 62748 52445 62812
rect 38217 62720 38281 62724
rect 38217 62664 38221 62720
rect 38221 62664 38277 62720
rect 38277 62664 38281 62720
rect 38217 62660 38281 62664
rect 38217 62640 38281 62644
rect 38217 62584 38221 62640
rect 38221 62584 38277 62640
rect 38277 62584 38281 62640
rect 38217 62580 38281 62584
rect 38217 62560 38281 62564
rect 38217 62504 38221 62560
rect 38221 62504 38277 62560
rect 38277 62504 38281 62560
rect 38217 62500 38281 62504
rect 38217 62480 38281 62484
rect 38217 62424 38221 62480
rect 38221 62424 38277 62480
rect 38277 62424 38281 62480
rect 38217 62420 38281 62424
rect 38217 62400 38281 62404
rect 38217 62344 38221 62400
rect 38221 62344 38277 62400
rect 38277 62344 38281 62400
rect 38217 62340 38281 62344
rect 38217 62320 38281 62324
rect 38217 62264 38221 62320
rect 38221 62264 38277 62320
rect 38277 62264 38281 62320
rect 38217 62260 38281 62264
rect 38217 62240 38281 62244
rect 38217 62184 38221 62240
rect 38221 62184 38277 62240
rect 38277 62184 38281 62240
rect 38217 62180 38281 62184
rect 38217 62160 38281 62164
rect 38217 62104 38221 62160
rect 38221 62104 38277 62160
rect 38277 62104 38281 62160
rect 38217 62100 38281 62104
rect 38217 62080 38281 62084
rect 38217 62024 38221 62080
rect 38221 62024 38277 62080
rect 38277 62024 38281 62080
rect 38217 62020 38281 62024
rect 38217 62000 38281 62004
rect 38217 61944 38221 62000
rect 38221 61944 38277 62000
rect 38277 61944 38281 62000
rect 38217 61940 38281 61944
rect 38217 61920 38281 61924
rect 38217 61864 38221 61920
rect 38221 61864 38277 61920
rect 38277 61864 38281 61920
rect 38217 61860 38281 61864
rect 38217 61840 38281 61844
rect 38217 61784 38221 61840
rect 38221 61784 38277 61840
rect 38277 61784 38281 61840
rect 38217 61780 38281 61784
rect 38217 61760 38281 61764
rect 38217 61704 38221 61760
rect 38221 61704 38277 61760
rect 38277 61704 38281 61760
rect 38217 61700 38281 61704
rect 38217 61680 38281 61684
rect 38217 61624 38221 61680
rect 38221 61624 38277 61680
rect 38277 61624 38281 61680
rect 38217 61620 38281 61624
rect 46189 62405 46253 62469
rect 52971 62405 53035 62469
rect 41888 61839 42352 62303
rect 59616 62811 59680 62815
rect 59616 62755 59620 62811
rect 59620 62755 59676 62811
rect 59676 62755 59680 62811
rect 59616 62751 59680 62755
rect 59616 62731 59680 62735
rect 59616 62675 59620 62731
rect 59620 62675 59676 62731
rect 59676 62675 59680 62731
rect 59616 62671 59680 62675
rect 59626 62418 59690 62422
rect 59626 62362 59630 62418
rect 59630 62362 59686 62418
rect 59686 62362 59690 62418
rect 59626 62358 59690 62362
rect 70925 62394 70989 62458
rect 75339 62394 75403 62458
rect 82957 62376 83021 62440
rect 89508 62376 89572 62440
rect 59626 62338 59690 62342
rect 59626 62282 59630 62338
rect 59630 62282 59686 62338
rect 59686 62282 59690 62338
rect 59626 62278 59690 62282
rect 59626 62258 59690 62262
rect 59626 62202 59630 62258
rect 59630 62202 59686 62258
rect 59686 62202 59690 62258
rect 59626 62198 59690 62202
rect 59626 62178 59690 62182
rect 59626 62122 59630 62178
rect 59630 62122 59686 62178
rect 59686 62122 59690 62178
rect 59626 62118 59690 62122
rect 59626 62098 59690 62102
rect 59626 62042 59630 62098
rect 59630 62042 59686 62098
rect 59686 62042 59690 62098
rect 59626 62038 59690 62042
rect 49372 61857 49436 61921
rect 54696 61857 54760 61921
rect 56334 61857 56398 61921
rect 58567 61857 58631 61921
rect 38217 61600 38281 61604
rect 38217 61544 38221 61600
rect 38221 61544 38277 61600
rect 38277 61544 38281 61600
rect 38217 61540 38281 61544
rect 38217 61520 38281 61524
rect 38217 61464 38221 61520
rect 38221 61464 38277 61520
rect 38277 61464 38281 61520
rect 38217 61460 38281 61464
rect 38217 61440 38281 61444
rect 38217 61384 38221 61440
rect 38221 61384 38277 61440
rect 38277 61384 38281 61440
rect 38217 61380 38281 61384
rect 27464 61341 27528 61345
rect 27464 61285 27468 61341
rect 27468 61285 27524 61341
rect 27524 61285 27528 61341
rect 27464 61281 27528 61285
rect 27544 61341 27608 61345
rect 27544 61285 27548 61341
rect 27548 61285 27604 61341
rect 27604 61285 27608 61341
rect 27544 61281 27608 61285
rect 27624 61341 27688 61345
rect 27624 61285 27628 61341
rect 27628 61285 27684 61341
rect 27684 61285 27688 61341
rect 27624 61281 27688 61285
rect 27704 61341 27768 61345
rect 27704 61285 27708 61341
rect 27708 61285 27764 61341
rect 27764 61285 27768 61341
rect 27704 61281 27768 61285
rect 27784 61341 27848 61345
rect 27784 61285 27788 61341
rect 27788 61285 27844 61341
rect 27844 61285 27848 61341
rect 27784 61281 27848 61285
rect 27864 61341 27928 61345
rect 27864 61285 27868 61341
rect 27868 61285 27924 61341
rect 27924 61285 27928 61341
rect 27864 61281 27928 61285
rect 30025 61359 30089 61363
rect 30025 61303 30029 61359
rect 30029 61303 30085 61359
rect 30085 61303 30089 61359
rect 30025 61299 30089 61303
rect 30025 61279 30089 61283
rect 30025 61223 30029 61279
rect 30029 61223 30085 61279
rect 30085 61223 30089 61279
rect 30025 61219 30089 61223
rect 30025 61199 30089 61203
rect 30025 61143 30029 61199
rect 30029 61143 30085 61199
rect 30085 61143 30089 61199
rect 30025 61139 30089 61143
rect 30025 61119 30089 61123
rect 30025 61063 30029 61119
rect 30029 61063 30085 61119
rect 30085 61063 30089 61119
rect 30025 61059 30089 61063
rect 30025 61039 30089 61043
rect 30025 60983 30029 61039
rect 30029 60983 30085 61039
rect 30085 60983 30089 61039
rect 30025 60979 30089 60983
rect 30025 60959 30089 60963
rect 30025 60903 30029 60959
rect 30029 60903 30085 60959
rect 30085 60903 30089 60959
rect 30025 60899 30089 60903
rect 30025 60879 30089 60883
rect 30025 60823 30029 60879
rect 30029 60823 30085 60879
rect 30085 60823 30089 60879
rect 30025 60819 30089 60823
rect 30025 60799 30089 60803
rect 30025 60743 30029 60799
rect 30029 60743 30085 60799
rect 30085 60743 30089 60799
rect 30025 60739 30089 60743
rect 30025 60719 30089 60723
rect 30025 60663 30029 60719
rect 30029 60663 30085 60719
rect 30085 60663 30089 60719
rect 30025 60659 30089 60663
rect 30025 60639 30089 60643
rect 30025 60583 30029 60639
rect 30029 60583 30085 60639
rect 30085 60583 30089 60639
rect 30025 60579 30089 60583
rect 30025 60559 30089 60563
rect 30025 60503 30029 60559
rect 30029 60503 30085 60559
rect 30085 60503 30089 60559
rect 30025 60499 30089 60503
rect 38217 61360 38281 61364
rect 38217 61304 38221 61360
rect 38221 61304 38277 61360
rect 38277 61304 38281 61360
rect 38217 61300 38281 61304
rect 48614 61329 48678 61393
rect 54279 61329 54343 61393
rect 56334 61328 56398 61392
rect 38217 61280 38281 61284
rect 38217 61224 38221 61280
rect 38221 61224 38277 61280
rect 38277 61224 38281 61280
rect 38217 61220 38281 61224
rect 38217 61200 38281 61204
rect 38217 61144 38221 61200
rect 38221 61144 38277 61200
rect 38277 61144 38281 61200
rect 38217 61140 38281 61144
rect 71680 61819 71744 61883
rect 75885 61819 75949 61883
rect 83500 61796 83564 61860
rect 88918 61796 88982 61860
rect 59090 61328 59154 61392
rect 38217 61120 38281 61124
rect 38217 61064 38221 61120
rect 38221 61064 38277 61120
rect 38277 61064 38281 61120
rect 38217 61060 38281 61064
rect 38217 61040 38281 61044
rect 38217 60984 38221 61040
rect 38221 60984 38277 61040
rect 38277 60984 38281 61040
rect 38217 60980 38281 60984
rect 38217 60960 38281 60964
rect 38217 60904 38221 60960
rect 38221 60904 38277 60960
rect 38277 60904 38281 60960
rect 38217 60900 38281 60904
rect 38217 60880 38281 60884
rect 38217 60824 38221 60880
rect 38221 60824 38277 60880
rect 38277 60824 38281 60880
rect 38217 60820 38281 60824
rect 38217 60800 38281 60804
rect 38217 60744 38221 60800
rect 38221 60744 38277 60800
rect 38277 60744 38281 60800
rect 38217 60740 38281 60744
rect 38217 60720 38281 60724
rect 38217 60664 38221 60720
rect 38221 60664 38277 60720
rect 38277 60664 38281 60720
rect 38217 60660 38281 60664
rect 38217 60640 38281 60644
rect 38217 60584 38221 60640
rect 38221 60584 38277 60640
rect 38277 60584 38281 60640
rect 38217 60580 38281 60584
rect 38217 60560 38281 60564
rect 38217 60504 38221 60560
rect 38221 60504 38277 60560
rect 38277 60504 38281 60560
rect 38217 60500 38281 60504
rect 38217 60480 38281 60484
rect 38217 60424 38221 60480
rect 38221 60424 38277 60480
rect 38277 60424 38281 60480
rect 38217 60420 38281 60424
rect 38217 60400 38281 60404
rect 38217 60344 38221 60400
rect 38221 60344 38277 60400
rect 38277 60344 38281 60400
rect 38217 60340 38281 60344
rect 72324 61268 72388 61332
rect 76431 61268 76495 61332
rect 87850 61187 87914 61251
rect 88325 61187 88389 61251
rect 59262 61153 59326 61157
rect 59262 61097 59266 61153
rect 59266 61097 59322 61153
rect 59322 61097 59326 61153
rect 59262 61093 59326 61097
rect 59262 61073 59326 61077
rect 59262 61017 59266 61073
rect 59266 61017 59322 61073
rect 59322 61017 59326 61073
rect 59262 61013 59326 61017
rect 59262 60993 59326 60997
rect 59262 60937 59266 60993
rect 59266 60937 59322 60993
rect 59322 60937 59326 60993
rect 59262 60933 59326 60937
rect 73084 60686 73148 60750
rect 76976 60686 77040 60750
rect 59263 60669 59327 60673
rect 59263 60613 59267 60669
rect 59267 60613 59323 60669
rect 59323 60613 59327 60669
rect 59263 60609 59327 60613
rect 59263 60589 59327 60593
rect 59263 60533 59267 60589
rect 59267 60533 59323 60589
rect 59323 60533 59327 60589
rect 59263 60529 59327 60533
rect 59263 60509 59327 60513
rect 59263 60453 59267 60509
rect 59267 60453 59323 60509
rect 59323 60453 59327 60509
rect 59263 60449 59327 60453
rect 59263 60429 59327 60433
rect 59263 60373 59267 60429
rect 59267 60373 59323 60429
rect 59323 60373 59327 60429
rect 59263 60369 59327 60373
rect 38217 60320 38281 60324
rect 38217 60264 38221 60320
rect 38221 60264 38277 60320
rect 38277 60264 38281 60320
rect 38217 60260 38281 60264
rect 59263 60349 59327 60353
rect 59263 60293 59267 60349
rect 59267 60293 59323 60349
rect 59323 60293 59327 60349
rect 59263 60289 59327 60293
rect 30025 60142 30089 60146
rect 30025 60086 30029 60142
rect 30029 60086 30085 60142
rect 30085 60086 30089 60142
rect 30025 60082 30089 60086
rect 38217 60240 38281 60244
rect 38217 60184 38221 60240
rect 38221 60184 38277 60240
rect 38277 60184 38281 60240
rect 38217 60180 38281 60184
rect 30025 60062 30089 60066
rect 30025 60006 30029 60062
rect 30029 60006 30085 60062
rect 30085 60006 30089 60062
rect 30025 60002 30089 60006
rect 30025 59982 30089 59986
rect 30025 59926 30029 59982
rect 30029 59926 30085 59982
rect 30085 59926 30089 59982
rect 30025 59922 30089 59926
rect 87316 60551 87380 60615
rect 87678 60551 87742 60615
rect 60678 60112 60742 60116
rect 60678 60056 60682 60112
rect 60682 60056 60738 60112
rect 60738 60056 60742 60112
rect 60678 60052 60742 60056
rect 60758 60112 60822 60116
rect 60758 60056 60762 60112
rect 60762 60056 60818 60112
rect 60818 60056 60822 60112
rect 60758 60052 60822 60056
rect 60838 60112 60902 60116
rect 60838 60056 60842 60112
rect 60842 60056 60898 60112
rect 60898 60056 60902 60112
rect 60838 60052 60902 60056
rect 62185 60111 62249 60115
rect 62265 60111 62329 60115
rect 62345 60111 62409 60115
rect 62185 60055 62205 60111
rect 62205 60055 62229 60111
rect 62229 60055 62249 60111
rect 62265 60055 62285 60111
rect 62285 60055 62309 60111
rect 62309 60055 62329 60111
rect 62345 60055 62365 60111
rect 62365 60055 62389 60111
rect 62389 60055 62409 60111
rect 62185 60051 62249 60055
rect 62265 60051 62329 60055
rect 62345 60051 62409 60055
rect 30025 59902 30089 59906
rect 30025 59846 30029 59902
rect 30029 59846 30085 59902
rect 30085 59846 30089 59902
rect 30025 59842 30089 59846
rect 47886 59899 47950 59963
rect 30025 59822 30089 59826
rect 30025 59766 30029 59822
rect 30029 59766 30085 59822
rect 30085 59766 30089 59822
rect 30025 59762 30089 59766
rect 30025 59742 30089 59746
rect 30025 59686 30029 59742
rect 30029 59686 30085 59742
rect 30085 59686 30089 59742
rect 30025 59682 30089 59686
rect 62669 60112 62733 60116
rect 62669 60056 62673 60112
rect 62673 60056 62729 60112
rect 62729 60056 62733 60112
rect 62669 60052 62733 60056
rect 62749 60112 62813 60116
rect 62749 60056 62753 60112
rect 62753 60056 62809 60112
rect 62809 60056 62813 60112
rect 62749 60052 62813 60056
rect 62829 60112 62893 60116
rect 62829 60056 62833 60112
rect 62833 60056 62889 60112
rect 62889 60056 62893 60112
rect 62829 60052 62893 60056
rect 30025 59662 30089 59666
rect 30025 59606 30029 59662
rect 30029 59606 30085 59662
rect 30085 59606 30089 59662
rect 30025 59602 30089 59606
rect 30025 59582 30089 59586
rect 30025 59526 30029 59582
rect 30029 59526 30085 59582
rect 30085 59526 30089 59582
rect 30025 59522 30089 59526
rect 60242 59602 60306 59666
rect 30025 59502 30089 59506
rect 30025 59446 30029 59502
rect 30029 59446 30085 59502
rect 30085 59446 30089 59502
rect 30025 59442 30089 59446
rect 30025 59422 30089 59426
rect 30025 59366 30029 59422
rect 30029 59366 30085 59422
rect 30085 59366 30089 59422
rect 30025 59362 30089 59366
rect 64068 60104 64132 60108
rect 64148 60104 64212 60108
rect 64068 60048 64088 60104
rect 64088 60048 64112 60104
rect 64112 60048 64132 60104
rect 64148 60048 64168 60104
rect 64168 60048 64192 60104
rect 64192 60048 64212 60104
rect 64068 60044 64132 60048
rect 64148 60044 64212 60048
rect 66670 60107 66734 60111
rect 66670 60051 66674 60107
rect 66674 60051 66730 60107
rect 66730 60051 66734 60107
rect 66670 60047 66734 60051
rect 66750 60107 66814 60111
rect 66750 60051 66754 60107
rect 66754 60051 66810 60107
rect 66810 60051 66814 60107
rect 66750 60047 66814 60051
rect 66830 60107 66894 60111
rect 66830 60051 66834 60107
rect 66834 60051 66890 60107
rect 66890 60051 66894 60107
rect 66830 60047 66894 60051
rect 73815 60008 73879 60072
rect 80239 60008 80303 60072
rect 86767 59928 86831 59992
rect 87084 59928 87148 59992
rect 64624 59571 64688 59635
rect 66191 59580 66255 59644
rect 30025 59342 30089 59346
rect 30025 59286 30029 59342
rect 30029 59286 30085 59342
rect 30085 59286 30089 59342
rect 30025 59282 30089 59286
rect 47025 59309 47089 59373
rect 74506 59301 74570 59365
rect 79692 59301 79756 59365
rect 30025 59262 30089 59266
rect 30025 59206 30029 59262
rect 30029 59206 30085 59262
rect 30085 59206 30089 59262
rect 30025 59202 30089 59206
rect 86223 59216 86287 59280
rect 86501 59216 86565 59280
rect 30025 59182 30089 59186
rect 30025 59126 30029 59182
rect 30029 59126 30085 59182
rect 30085 59126 30089 59182
rect 30025 59122 30089 59126
rect 30025 59102 30089 59106
rect 30025 59046 30029 59102
rect 30029 59046 30085 59102
rect 30085 59046 30089 59102
rect 30025 59042 30089 59046
rect 30022 58704 30086 58708
rect 30022 58648 30026 58704
rect 30026 58648 30082 58704
rect 30082 58648 30086 58704
rect 30022 58644 30086 58648
rect 43699 58634 43763 58698
rect 30022 58624 30086 58628
rect 30022 58568 30026 58624
rect 30026 58568 30082 58624
rect 30082 58568 30086 58624
rect 30022 58564 30086 58568
rect 30022 58544 30086 58548
rect 30022 58488 30026 58544
rect 30026 58488 30082 58544
rect 30082 58488 30086 58544
rect 30022 58484 30086 58488
rect 75346 58541 75410 58605
rect 79150 58541 79214 58605
rect 84042 58480 84106 58544
rect 85922 58480 85986 58544
rect 30022 58464 30086 58468
rect 30022 58408 30026 58464
rect 30026 58408 30082 58464
rect 30082 58408 30086 58464
rect 30022 58404 30086 58408
rect 30022 58384 30086 58388
rect 30022 58328 30026 58384
rect 30026 58328 30082 58384
rect 30082 58328 30086 58384
rect 30022 58324 30086 58328
rect 30022 58304 30086 58308
rect 30022 58248 30026 58304
rect 30026 58248 30082 58304
rect 30082 58248 30086 58304
rect 30022 58244 30086 58248
rect 30022 58224 30086 58228
rect 30022 58168 30026 58224
rect 30026 58168 30082 58224
rect 30082 58168 30086 58224
rect 30022 58164 30086 58168
rect 52381 58153 52445 58217
rect 30022 58144 30086 58148
rect 30022 58088 30026 58144
rect 30026 58088 30082 58144
rect 30082 58088 30086 58144
rect 30022 58084 30086 58088
rect 30022 58064 30086 58068
rect 30022 58008 30026 58064
rect 30026 58008 30082 58064
rect 30082 58008 30086 58064
rect 30022 58004 30086 58008
rect 30022 57984 30086 57988
rect 30022 57928 30026 57984
rect 30026 57928 30082 57984
rect 30082 57928 30086 57984
rect 30022 57924 30086 57928
rect 30022 57904 30086 57908
rect 30022 57848 30026 57904
rect 30026 57848 30082 57904
rect 30082 57848 30086 57904
rect 30022 57844 30086 57848
rect 30022 57824 30086 57828
rect 30022 57768 30026 57824
rect 30026 57768 30082 57824
rect 30082 57768 30086 57824
rect 30022 57764 30086 57768
rect 52971 57808 53035 57872
rect 84599 57771 84663 57835
rect 85409 57771 85473 57835
rect 30022 57744 30086 57748
rect 30022 57688 30026 57744
rect 30026 57688 30082 57744
rect 30082 57688 30086 57744
rect 30022 57684 30086 57688
rect 76349 57704 76413 57768
rect 78607 57704 78671 57768
rect 30022 57664 30086 57668
rect 30022 57608 30026 57664
rect 30026 57608 30082 57664
rect 30082 57608 30086 57664
rect 30022 57604 30086 57608
rect 30022 57584 30086 57588
rect 30022 57528 30026 57584
rect 30026 57528 30082 57584
rect 30082 57528 30086 57584
rect 30022 57524 30086 57528
rect 35576 57569 35640 57573
rect 35576 57513 35580 57569
rect 35580 57513 35636 57569
rect 35636 57513 35640 57569
rect 35576 57509 35640 57513
rect 41955 57137 42019 57201
rect 30017 56882 30081 56886
rect 30017 56826 30021 56882
rect 30021 56826 30077 56882
rect 30077 56826 30081 56882
rect 30017 56822 30081 56826
rect 30017 56802 30081 56806
rect 30017 56746 30021 56802
rect 30021 56746 30077 56802
rect 30077 56746 30081 56802
rect 30017 56742 30081 56746
rect 30017 56722 30081 56726
rect 30017 56666 30021 56722
rect 30021 56666 30077 56722
rect 30077 56666 30081 56722
rect 30017 56662 30081 56666
rect 30017 56642 30081 56646
rect 30017 56586 30021 56642
rect 30021 56586 30077 56642
rect 30077 56586 30081 56642
rect 30017 56582 30081 56586
rect 30017 56562 30081 56566
rect 30017 56506 30021 56562
rect 30021 56506 30077 56562
rect 30077 56506 30081 56562
rect 30017 56502 30081 56506
rect 30017 56482 30081 56486
rect 30017 56426 30021 56482
rect 30021 56426 30077 56482
rect 30077 56426 30081 56482
rect 30017 56422 30081 56426
rect 65059 55829 65123 55833
rect 65059 55773 65063 55829
rect 65063 55773 65119 55829
rect 65119 55773 65123 55829
rect 65059 55769 65123 55773
rect 68441 55349 68505 55413
rect 70925 55349 70989 55413
rect 61448 54450 61512 54454
rect 61448 54394 61452 54450
rect 61452 54394 61508 54450
rect 61508 54394 61512 54450
rect 61448 54390 61512 54394
rect 65422 54455 65486 54459
rect 65422 54399 65426 54455
rect 65426 54399 65482 54455
rect 65482 54399 65486 54455
rect 65422 54395 65486 54399
rect 69060 54730 69124 54794
rect 71680 54730 71744 54794
rect 60420 54323 60484 54327
rect 60420 54267 60424 54323
rect 60424 54267 60480 54323
rect 60480 54267 60484 54323
rect 60420 54263 60484 54267
rect 53176 53710 53240 53774
rect 51815 53287 51879 53351
rect 73815 53770 73879 53774
rect 73815 53714 73819 53770
rect 73819 53714 73875 53770
rect 73875 53714 73879 53770
rect 73815 53710 73879 53714
rect 74506 53347 74570 53351
rect 74506 53291 74510 53347
rect 74510 53291 74566 53347
rect 74566 53291 74570 53347
rect 74506 53287 74570 53291
rect 67727 52762 67791 52826
rect 69060 52762 69124 52826
rect 41399 52081 41463 52085
rect 41399 52025 41403 52081
rect 41403 52025 41459 52081
rect 41459 52025 41463 52081
rect 41399 52021 41463 52025
rect 41399 52001 41463 52005
rect 41399 51945 41403 52001
rect 41403 51945 41459 52001
rect 41459 51945 41463 52001
rect 41399 51941 41463 51945
rect 41399 51921 41463 51925
rect 41399 51865 41403 51921
rect 41403 51865 41459 51921
rect 41459 51865 41463 51921
rect 41399 51861 41463 51865
rect 41399 51841 41463 51845
rect 41399 51785 41403 51841
rect 41403 51785 41459 51841
rect 41459 51785 41463 51841
rect 41399 51781 41463 51785
rect 41399 51761 41463 51765
rect 41399 51705 41403 51761
rect 41403 51705 41459 51761
rect 41459 51705 41463 51761
rect 41399 51701 41463 51705
rect 44709 52083 44773 52087
rect 44709 52027 44713 52083
rect 44713 52027 44769 52083
rect 44769 52027 44773 52083
rect 44709 52023 44773 52027
rect 44709 52003 44773 52007
rect 44709 51947 44713 52003
rect 44713 51947 44769 52003
rect 44769 51947 44773 52003
rect 44709 51943 44773 51947
rect 44709 51923 44773 51927
rect 44709 51867 44713 51923
rect 44713 51867 44769 51923
rect 44769 51867 44773 51923
rect 44709 51863 44773 51867
rect 44709 51843 44773 51847
rect 44709 51787 44713 51843
rect 44713 51787 44769 51843
rect 44769 51787 44773 51843
rect 44709 51783 44773 51787
rect 44709 51763 44773 51767
rect 44709 51707 44713 51763
rect 44713 51707 44769 51763
rect 44769 51707 44773 51763
rect 44709 51703 44773 51707
rect 39491 51630 39555 51634
rect 39491 51574 39495 51630
rect 39495 51574 39551 51630
rect 39551 51574 39555 51630
rect 39491 51570 39555 51574
rect 51815 51550 51879 51554
rect 51815 51494 51819 51550
rect 51819 51494 51875 51550
rect 51875 51494 51879 51550
rect 51815 51490 51879 51494
rect 44716 51442 44780 51446
rect 44716 51386 44720 51442
rect 44720 51386 44776 51442
rect 44776 51386 44780 51442
rect 44716 51382 44780 51386
rect 44716 51362 44780 51366
rect 44716 51306 44720 51362
rect 44720 51306 44776 51362
rect 44776 51306 44780 51362
rect 44716 51302 44780 51306
rect 44716 51282 44780 51286
rect 44716 51226 44720 51282
rect 44720 51226 44776 51282
rect 44776 51226 44780 51282
rect 44716 51222 44780 51226
rect 53176 50873 53240 50877
rect 53176 50817 53180 50873
rect 53180 50817 53236 50873
rect 53236 50817 53240 50873
rect 53176 50813 53240 50817
rect 18939 50612 19003 50616
rect 18939 50556 18943 50612
rect 18943 50556 18999 50612
rect 18999 50556 19003 50612
rect 18939 50552 19003 50556
rect 19019 50612 19083 50616
rect 19019 50556 19023 50612
rect 19023 50556 19079 50612
rect 19079 50556 19083 50612
rect 19019 50552 19083 50556
rect 19099 50612 19163 50616
rect 19099 50556 19103 50612
rect 19103 50556 19159 50612
rect 19159 50556 19163 50612
rect 19099 50552 19163 50556
rect 19179 50612 19243 50616
rect 19179 50556 19183 50612
rect 19183 50556 19239 50612
rect 19239 50556 19243 50612
rect 19179 50552 19243 50556
rect 19259 50612 19323 50616
rect 19259 50556 19263 50612
rect 19263 50556 19319 50612
rect 19319 50556 19323 50612
rect 19259 50552 19323 50556
rect 19339 50612 19403 50616
rect 19339 50556 19343 50612
rect 19343 50556 19399 50612
rect 19399 50556 19403 50612
rect 19339 50552 19403 50556
rect 19419 50612 19483 50616
rect 19419 50556 19423 50612
rect 19423 50556 19479 50612
rect 19479 50556 19483 50612
rect 19419 50552 19483 50556
rect 19499 50612 19563 50616
rect 19499 50556 19503 50612
rect 19503 50556 19559 50612
rect 19559 50556 19563 50612
rect 19499 50552 19563 50556
rect 19579 50612 19643 50616
rect 19579 50556 19583 50612
rect 19583 50556 19639 50612
rect 19639 50556 19643 50612
rect 19579 50552 19643 50556
rect 19659 50612 19723 50616
rect 19659 50556 19663 50612
rect 19663 50556 19719 50612
rect 19719 50556 19723 50612
rect 19659 50552 19723 50556
rect 19739 50612 19803 50616
rect 19739 50556 19743 50612
rect 19743 50556 19799 50612
rect 19799 50556 19803 50612
rect 19739 50552 19803 50556
rect 19819 50612 19883 50616
rect 19819 50556 19823 50612
rect 19823 50556 19879 50612
rect 19879 50556 19883 50612
rect 19819 50552 19883 50556
rect 19899 50612 19963 50616
rect 19899 50556 19903 50612
rect 19903 50556 19959 50612
rect 19959 50556 19963 50612
rect 19899 50552 19963 50556
rect 19979 50612 20043 50616
rect 19979 50556 19983 50612
rect 19983 50556 20039 50612
rect 20039 50556 20043 50612
rect 19979 50552 20043 50556
rect 20059 50612 20123 50616
rect 20059 50556 20063 50612
rect 20063 50556 20119 50612
rect 20119 50556 20123 50612
rect 20059 50552 20123 50556
rect 20139 50612 20203 50616
rect 20139 50556 20143 50612
rect 20143 50556 20199 50612
rect 20199 50556 20203 50612
rect 20139 50552 20203 50556
rect 20219 50612 20283 50616
rect 20219 50556 20223 50612
rect 20223 50556 20279 50612
rect 20279 50556 20283 50612
rect 20219 50552 20283 50556
rect 20299 50612 20363 50616
rect 20299 50556 20303 50612
rect 20303 50556 20359 50612
rect 20359 50556 20363 50612
rect 20299 50552 20363 50556
rect 20379 50612 20443 50616
rect 20379 50556 20383 50612
rect 20383 50556 20439 50612
rect 20439 50556 20443 50612
rect 20379 50552 20443 50556
rect 20459 50612 20523 50616
rect 20459 50556 20463 50612
rect 20463 50556 20519 50612
rect 20519 50556 20523 50612
rect 20459 50552 20523 50556
rect 20539 50612 20603 50616
rect 20539 50556 20543 50612
rect 20543 50556 20599 50612
rect 20599 50556 20603 50612
rect 20539 50552 20603 50556
rect 20619 50612 20683 50616
rect 20619 50556 20623 50612
rect 20623 50556 20679 50612
rect 20679 50556 20683 50612
rect 20619 50552 20683 50556
rect 20699 50612 20763 50616
rect 20699 50556 20703 50612
rect 20703 50556 20759 50612
rect 20759 50556 20763 50612
rect 20699 50552 20763 50556
rect 20779 50612 20843 50616
rect 20779 50556 20783 50612
rect 20783 50556 20839 50612
rect 20839 50556 20843 50612
rect 20779 50552 20843 50556
rect 20859 50612 20923 50616
rect 20859 50556 20863 50612
rect 20863 50556 20919 50612
rect 20919 50556 20923 50612
rect 20859 50552 20923 50556
rect 20939 50612 21003 50616
rect 20939 50556 20943 50612
rect 20943 50556 20999 50612
rect 20999 50556 21003 50612
rect 20939 50552 21003 50556
rect 21019 50612 21083 50616
rect 21019 50556 21023 50612
rect 21023 50556 21079 50612
rect 21079 50556 21083 50612
rect 21019 50552 21083 50556
rect 21099 50612 21163 50616
rect 21099 50556 21103 50612
rect 21103 50556 21159 50612
rect 21159 50556 21163 50612
rect 21099 50552 21163 50556
rect 21179 50612 21243 50616
rect 21179 50556 21183 50612
rect 21183 50556 21239 50612
rect 21239 50556 21243 50612
rect 21179 50552 21243 50556
rect 21259 50612 21323 50616
rect 21259 50556 21263 50612
rect 21263 50556 21319 50612
rect 21319 50556 21323 50612
rect 21259 50552 21323 50556
rect 21339 50612 21403 50616
rect 21339 50556 21343 50612
rect 21343 50556 21399 50612
rect 21399 50556 21403 50612
rect 21339 50552 21403 50556
rect 21419 50612 21483 50616
rect 21419 50556 21423 50612
rect 21423 50556 21479 50612
rect 21479 50556 21483 50612
rect 21419 50552 21483 50556
rect 21499 50612 21563 50616
rect 21499 50556 21503 50612
rect 21503 50556 21559 50612
rect 21559 50556 21563 50612
rect 21499 50552 21563 50556
rect 21579 50612 21643 50616
rect 21579 50556 21583 50612
rect 21583 50556 21639 50612
rect 21639 50556 21643 50612
rect 21579 50552 21643 50556
rect 21659 50612 21723 50616
rect 21659 50556 21663 50612
rect 21663 50556 21719 50612
rect 21719 50556 21723 50612
rect 21659 50552 21723 50556
rect 21739 50612 21803 50616
rect 21739 50556 21743 50612
rect 21743 50556 21799 50612
rect 21799 50556 21803 50612
rect 21739 50552 21803 50556
rect 21819 50612 21883 50616
rect 21819 50556 21823 50612
rect 21823 50556 21879 50612
rect 21879 50556 21883 50612
rect 21819 50552 21883 50556
rect 21899 50612 21963 50616
rect 21899 50556 21903 50612
rect 21903 50556 21959 50612
rect 21959 50556 21963 50612
rect 21899 50552 21963 50556
rect 21979 50612 22043 50616
rect 21979 50556 21983 50612
rect 21983 50556 22039 50612
rect 22039 50556 22043 50612
rect 21979 50552 22043 50556
rect 22059 50612 22123 50616
rect 22059 50556 22063 50612
rect 22063 50556 22119 50612
rect 22119 50556 22123 50612
rect 22059 50552 22123 50556
rect 22139 50612 22203 50616
rect 22139 50556 22143 50612
rect 22143 50556 22199 50612
rect 22199 50556 22203 50612
rect 22139 50552 22203 50556
rect 39491 50401 39555 50405
rect 39491 50345 39495 50401
rect 39495 50345 39551 50401
rect 39551 50345 39555 50401
rect 39491 50341 39555 50345
rect 44713 50481 44777 50485
rect 44713 50425 44717 50481
rect 44717 50425 44773 50481
rect 44773 50425 44777 50481
rect 44713 50421 44777 50425
rect 44713 50401 44777 50405
rect 44713 50345 44717 50401
rect 44717 50345 44773 50401
rect 44773 50345 44777 50401
rect 44713 50341 44777 50345
rect 41381 50292 41445 50296
rect 41381 50236 41385 50292
rect 41385 50236 41441 50292
rect 41441 50236 41445 50292
rect 41381 50232 41445 50236
rect 41381 50212 41445 50216
rect 41381 50156 41385 50212
rect 41385 50156 41441 50212
rect 41441 50156 41445 50212
rect 41381 50152 41445 50156
rect 41381 50132 41445 50136
rect 41381 50076 41385 50132
rect 41385 50076 41441 50132
rect 41441 50076 41445 50132
rect 41381 50072 41445 50076
rect 44713 50321 44777 50325
rect 44713 50265 44717 50321
rect 44717 50265 44773 50321
rect 44773 50265 44777 50321
rect 44713 50261 44777 50265
rect 68441 50308 68505 50372
rect 68931 50308 68995 50372
rect 44713 50241 44777 50245
rect 44713 50185 44717 50241
rect 44717 50185 44773 50241
rect 44773 50185 44777 50241
rect 44713 50181 44777 50185
rect 44713 50161 44777 50165
rect 44713 50105 44717 50161
rect 44717 50105 44773 50161
rect 44773 50105 44777 50161
rect 44713 50101 44777 50105
rect 70944 49967 71008 50031
rect 82973 49967 83037 50031
rect 38010 49597 38234 49821
rect 31653 49498 31717 49502
rect 31653 49442 31657 49498
rect 31657 49442 31713 49498
rect 31713 49442 31717 49498
rect 31653 49438 31717 49442
rect 31653 49418 31717 49422
rect 31653 49362 31657 49418
rect 31657 49362 31713 49418
rect 31713 49362 31717 49418
rect 31653 49358 31717 49362
rect 31653 49338 31717 49342
rect 31653 49282 31657 49338
rect 31657 49282 31713 49338
rect 31713 49282 31717 49338
rect 31653 49278 31717 49282
rect 31653 49258 31717 49262
rect 31653 49202 31657 49258
rect 31657 49202 31713 49258
rect 31713 49202 31717 49258
rect 31653 49198 31717 49202
rect 45770 49622 45834 49686
rect 70360 49556 70424 49620
rect 83557 49556 83621 49620
rect 31653 48959 31717 48963
rect 31653 48903 31657 48959
rect 31657 48903 31713 48959
rect 31713 48903 31717 48959
rect 31653 48899 31717 48903
rect 39491 48988 39555 48992
rect 39491 48932 39495 48988
rect 39495 48932 39551 48988
rect 39551 48932 39555 48988
rect 39491 48928 39555 48932
rect 31653 48879 31717 48883
rect 31653 48823 31657 48879
rect 31657 48823 31713 48879
rect 31713 48823 31717 48879
rect 31653 48819 31717 48823
rect 45117 48830 45181 48894
rect 64695 48806 64759 48870
rect 72324 48806 72388 48870
rect 31653 48799 31717 48803
rect 31653 48743 31657 48799
rect 31657 48743 31713 48799
rect 31713 48743 31717 48799
rect 31653 48739 31717 48743
rect 44701 48715 44765 48719
rect 44701 48659 44705 48715
rect 44705 48659 44761 48715
rect 44761 48659 44765 48715
rect 44701 48655 44765 48659
rect 44701 48635 44765 48639
rect 44701 48579 44705 48635
rect 44705 48579 44761 48635
rect 44761 48579 44765 48635
rect 44701 48575 44765 48579
rect 44701 48555 44765 48559
rect 44701 48499 44705 48555
rect 44705 48499 44761 48555
rect 44761 48499 44765 48555
rect 44701 48495 44765 48499
rect 62811 48600 62875 48604
rect 62811 48544 62815 48600
rect 62815 48544 62871 48600
rect 62871 48544 62875 48600
rect 62811 48540 62875 48544
rect 64360 48551 64424 48615
rect 62811 48520 62875 48524
rect 62811 48464 62815 48520
rect 62815 48464 62871 48520
rect 62871 48464 62875 48520
rect 62811 48460 62875 48464
rect 65223 48488 65287 48552
rect 73084 48488 73148 48552
rect 62811 48440 62875 48444
rect 62811 48384 62815 48440
rect 62815 48384 62871 48440
rect 62871 48384 62875 48440
rect 62811 48380 62875 48384
rect 62811 48360 62875 48364
rect 62811 48304 62815 48360
rect 62815 48304 62871 48360
rect 62871 48304 62875 48360
rect 62811 48300 62875 48304
rect 44705 48251 44769 48255
rect 44705 48195 44709 48251
rect 44709 48195 44765 48251
rect 44765 48195 44769 48251
rect 44705 48191 44769 48195
rect 62811 48280 62875 48284
rect 62811 48224 62815 48280
rect 62815 48224 62871 48280
rect 62871 48224 62875 48280
rect 62811 48220 62875 48224
rect 44705 48171 44769 48175
rect 44705 48115 44709 48171
rect 44709 48115 44765 48171
rect 44765 48115 44769 48171
rect 44705 48111 44769 48115
rect 68174 48160 68238 48224
rect 44705 48091 44769 48095
rect 44705 48035 44709 48091
rect 44709 48035 44765 48091
rect 44765 48035 44769 48091
rect 44705 48031 44769 48035
rect 45770 47845 45834 47909
rect 64360 47845 64424 47909
rect 76349 47845 76413 47909
rect 39491 47759 39555 47763
rect 39491 47703 39495 47759
rect 39495 47703 39551 47759
rect 39551 47703 39555 47759
rect 39491 47699 39555 47703
rect 18945 47604 19009 47608
rect 18945 47548 18949 47604
rect 18949 47548 19005 47604
rect 19005 47548 19009 47604
rect 18945 47544 19009 47548
rect 19025 47604 19089 47608
rect 19025 47548 19029 47604
rect 19029 47548 19085 47604
rect 19085 47548 19089 47604
rect 19025 47544 19089 47548
rect 19105 47604 19169 47608
rect 19105 47548 19109 47604
rect 19109 47548 19165 47604
rect 19165 47548 19169 47604
rect 19105 47544 19169 47548
rect 19185 47604 19249 47608
rect 19185 47548 19189 47604
rect 19189 47548 19245 47604
rect 19245 47548 19249 47604
rect 19185 47544 19249 47548
rect 19265 47604 19329 47608
rect 19265 47548 19269 47604
rect 19269 47548 19325 47604
rect 19325 47548 19329 47604
rect 19265 47544 19329 47548
rect 19345 47604 19409 47608
rect 19345 47548 19349 47604
rect 19349 47548 19405 47604
rect 19405 47548 19409 47604
rect 19345 47544 19409 47548
rect 19425 47604 19489 47608
rect 19425 47548 19429 47604
rect 19429 47548 19485 47604
rect 19485 47548 19489 47604
rect 19425 47544 19489 47548
rect 19505 47604 19569 47608
rect 19505 47548 19509 47604
rect 19509 47548 19565 47604
rect 19565 47548 19569 47604
rect 19505 47544 19569 47548
rect 19585 47604 19649 47608
rect 19585 47548 19589 47604
rect 19589 47548 19645 47604
rect 19645 47548 19649 47604
rect 19585 47544 19649 47548
rect 19665 47604 19729 47608
rect 19665 47548 19669 47604
rect 19669 47548 19725 47604
rect 19725 47548 19729 47604
rect 19665 47544 19729 47548
rect 19745 47604 19809 47608
rect 19745 47548 19749 47604
rect 19749 47548 19805 47604
rect 19805 47548 19809 47604
rect 19745 47544 19809 47548
rect 19825 47604 19889 47608
rect 19825 47548 19829 47604
rect 19829 47548 19885 47604
rect 19885 47548 19889 47604
rect 19825 47544 19889 47548
rect 19905 47604 19969 47608
rect 19905 47548 19909 47604
rect 19909 47548 19965 47604
rect 19965 47548 19969 47604
rect 19905 47544 19969 47548
rect 19985 47604 20049 47608
rect 19985 47548 19989 47604
rect 19989 47548 20045 47604
rect 20045 47548 20049 47604
rect 19985 47544 20049 47548
rect 20065 47604 20129 47608
rect 20065 47548 20069 47604
rect 20069 47548 20125 47604
rect 20125 47548 20129 47604
rect 20065 47544 20129 47548
rect 20145 47604 20209 47608
rect 20145 47548 20149 47604
rect 20149 47548 20205 47604
rect 20205 47548 20209 47604
rect 20145 47544 20209 47548
rect 20225 47604 20289 47608
rect 20225 47548 20229 47604
rect 20229 47548 20285 47604
rect 20285 47548 20289 47604
rect 20225 47544 20289 47548
rect 20305 47604 20369 47608
rect 20305 47548 20309 47604
rect 20309 47548 20365 47604
rect 20365 47548 20369 47604
rect 20305 47544 20369 47548
rect 20385 47604 20449 47608
rect 20385 47548 20389 47604
rect 20389 47548 20445 47604
rect 20445 47548 20449 47604
rect 20385 47544 20449 47548
rect 20465 47604 20529 47608
rect 20465 47548 20469 47604
rect 20469 47548 20525 47604
rect 20525 47548 20529 47604
rect 20465 47544 20529 47548
rect 20545 47604 20609 47608
rect 20545 47548 20549 47604
rect 20549 47548 20605 47604
rect 20605 47548 20609 47604
rect 20545 47544 20609 47548
rect 20625 47604 20689 47608
rect 20625 47548 20629 47604
rect 20629 47548 20685 47604
rect 20685 47548 20689 47604
rect 20625 47544 20689 47548
rect 20705 47604 20769 47608
rect 20705 47548 20709 47604
rect 20709 47548 20765 47604
rect 20765 47548 20769 47604
rect 20705 47544 20769 47548
rect 20785 47604 20849 47608
rect 20785 47548 20789 47604
rect 20789 47548 20845 47604
rect 20845 47548 20849 47604
rect 20785 47544 20849 47548
rect 20865 47604 20929 47608
rect 20865 47548 20869 47604
rect 20869 47548 20925 47604
rect 20925 47548 20929 47604
rect 20865 47544 20929 47548
rect 20945 47604 21009 47608
rect 20945 47548 20949 47604
rect 20949 47548 21005 47604
rect 21005 47548 21009 47604
rect 20945 47544 21009 47548
rect 21025 47604 21089 47608
rect 21025 47548 21029 47604
rect 21029 47548 21085 47604
rect 21085 47548 21089 47604
rect 21025 47544 21089 47548
rect 21105 47604 21169 47608
rect 21105 47548 21109 47604
rect 21109 47548 21165 47604
rect 21165 47548 21169 47604
rect 21105 47544 21169 47548
rect 21185 47604 21249 47608
rect 21185 47548 21189 47604
rect 21189 47548 21245 47604
rect 21245 47548 21249 47604
rect 21185 47544 21249 47548
rect 21265 47604 21329 47608
rect 21265 47548 21269 47604
rect 21269 47548 21325 47604
rect 21325 47548 21329 47604
rect 21265 47544 21329 47548
rect 21345 47604 21409 47608
rect 21345 47548 21349 47604
rect 21349 47548 21405 47604
rect 21405 47548 21409 47604
rect 21345 47544 21409 47548
rect 21425 47604 21489 47608
rect 21425 47548 21429 47604
rect 21429 47548 21485 47604
rect 21485 47548 21489 47604
rect 21425 47544 21489 47548
rect 21505 47604 21569 47608
rect 21505 47548 21509 47604
rect 21509 47548 21565 47604
rect 21565 47548 21569 47604
rect 21505 47544 21569 47548
rect 21585 47604 21649 47608
rect 21585 47548 21589 47604
rect 21589 47548 21645 47604
rect 21645 47548 21649 47604
rect 21585 47544 21649 47548
rect 21665 47604 21729 47608
rect 21665 47548 21669 47604
rect 21669 47548 21725 47604
rect 21725 47548 21729 47604
rect 21665 47544 21729 47548
rect 21745 47604 21809 47608
rect 21745 47548 21749 47604
rect 21749 47548 21805 47604
rect 21805 47548 21809 47604
rect 21745 47544 21809 47548
rect 21825 47604 21889 47608
rect 21825 47548 21829 47604
rect 21829 47548 21885 47604
rect 21885 47548 21889 47604
rect 21825 47544 21889 47548
rect 21905 47604 21969 47608
rect 21905 47548 21909 47604
rect 21909 47548 21965 47604
rect 21965 47548 21969 47604
rect 21905 47544 21969 47548
rect 21985 47604 22049 47608
rect 21985 47548 21989 47604
rect 21989 47548 22045 47604
rect 22045 47548 22049 47604
rect 21985 47544 22049 47548
rect 22065 47604 22129 47608
rect 22065 47548 22069 47604
rect 22069 47548 22125 47604
rect 22125 47548 22129 47604
rect 22065 47544 22129 47548
rect 22145 47604 22209 47608
rect 22145 47548 22149 47604
rect 22149 47548 22205 47604
rect 22205 47548 22209 47604
rect 22145 47544 22209 47548
rect 41370 47651 41434 47655
rect 41370 47595 41374 47651
rect 41374 47595 41430 47651
rect 41430 47595 41434 47651
rect 41370 47591 41434 47595
rect 41370 47571 41434 47575
rect 41370 47515 41374 47571
rect 41374 47515 41430 47571
rect 41430 47515 41434 47571
rect 41370 47511 41434 47515
rect 41370 47491 41434 47495
rect 41370 47435 41374 47491
rect 41374 47435 41430 47491
rect 41430 47435 41434 47491
rect 41370 47431 41434 47435
rect 45117 47476 45181 47540
rect 75346 47476 75410 47540
rect 44708 47277 44772 47281
rect 44708 47221 44712 47277
rect 44712 47221 44768 47277
rect 44768 47221 44772 47277
rect 44708 47217 44772 47221
rect 65887 47351 65951 47355
rect 65887 47295 65891 47351
rect 65891 47295 65947 47351
rect 65947 47295 65951 47351
rect 65887 47291 65951 47295
rect 65967 47351 66031 47355
rect 65967 47295 65971 47351
rect 65971 47295 66027 47351
rect 66027 47295 66031 47351
rect 65967 47291 66031 47295
rect 99985 48169 100049 48173
rect 99985 48113 99989 48169
rect 99989 48113 100045 48169
rect 100045 48113 100049 48169
rect 99985 48109 100049 48113
rect 100065 48169 100129 48173
rect 100065 48113 100069 48169
rect 100069 48113 100125 48169
rect 100125 48113 100129 48169
rect 100065 48109 100129 48113
rect 100145 48169 100209 48173
rect 100145 48113 100149 48169
rect 100149 48113 100205 48169
rect 100205 48113 100209 48169
rect 100145 48109 100209 48113
rect 100225 48169 100289 48173
rect 100225 48113 100229 48169
rect 100229 48113 100285 48169
rect 100285 48113 100289 48169
rect 100225 48109 100289 48113
rect 100305 48169 100369 48173
rect 100305 48113 100309 48169
rect 100309 48113 100365 48169
rect 100365 48113 100369 48169
rect 100305 48109 100369 48113
rect 100385 48169 100449 48173
rect 100385 48113 100389 48169
rect 100389 48113 100445 48169
rect 100445 48113 100449 48169
rect 100385 48109 100449 48113
rect 100465 48169 100529 48173
rect 100465 48113 100469 48169
rect 100469 48113 100525 48169
rect 100525 48113 100529 48169
rect 100465 48109 100529 48113
rect 100545 48169 100609 48173
rect 100545 48113 100549 48169
rect 100549 48113 100605 48169
rect 100605 48113 100609 48169
rect 100545 48109 100609 48113
rect 100625 48169 100689 48173
rect 100625 48113 100629 48169
rect 100629 48113 100685 48169
rect 100685 48113 100689 48169
rect 100625 48109 100689 48113
rect 100705 48169 100769 48173
rect 100705 48113 100709 48169
rect 100709 48113 100765 48169
rect 100765 48113 100769 48169
rect 100705 48109 100769 48113
rect 100785 48169 100849 48173
rect 100785 48113 100789 48169
rect 100789 48113 100845 48169
rect 100845 48113 100849 48169
rect 100785 48109 100849 48113
rect 100865 48169 100929 48173
rect 100865 48113 100869 48169
rect 100869 48113 100925 48169
rect 100925 48113 100929 48169
rect 100865 48109 100929 48113
rect 100945 48169 101009 48173
rect 100945 48113 100949 48169
rect 100949 48113 101005 48169
rect 101005 48113 101009 48169
rect 100945 48109 101009 48113
rect 101025 48169 101089 48173
rect 101025 48113 101029 48169
rect 101029 48113 101085 48169
rect 101085 48113 101089 48169
rect 101025 48109 101089 48113
rect 101105 48169 101169 48173
rect 101105 48113 101109 48169
rect 101109 48113 101165 48169
rect 101165 48113 101169 48169
rect 101105 48109 101169 48113
rect 101185 48169 101249 48173
rect 101185 48113 101189 48169
rect 101189 48113 101245 48169
rect 101245 48113 101249 48169
rect 101185 48109 101249 48113
rect 101265 48169 101329 48173
rect 101265 48113 101269 48169
rect 101269 48113 101325 48169
rect 101325 48113 101329 48169
rect 101265 48109 101329 48113
rect 101345 48169 101409 48173
rect 101345 48113 101349 48169
rect 101349 48113 101405 48169
rect 101405 48113 101409 48169
rect 101345 48109 101409 48113
rect 101425 48169 101489 48173
rect 101425 48113 101429 48169
rect 101429 48113 101485 48169
rect 101485 48113 101489 48169
rect 101425 48109 101489 48113
rect 101505 48169 101569 48173
rect 101505 48113 101509 48169
rect 101509 48113 101565 48169
rect 101565 48113 101569 48169
rect 101505 48109 101569 48113
rect 101585 48169 101649 48173
rect 101585 48113 101589 48169
rect 101589 48113 101645 48169
rect 101645 48113 101649 48169
rect 101585 48109 101649 48113
rect 101665 48169 101729 48173
rect 101665 48113 101669 48169
rect 101669 48113 101725 48169
rect 101725 48113 101729 48169
rect 101665 48109 101729 48113
rect 101745 48169 101809 48173
rect 101745 48113 101749 48169
rect 101749 48113 101805 48169
rect 101805 48113 101809 48169
rect 101745 48109 101809 48113
rect 101825 48169 101889 48173
rect 101825 48113 101829 48169
rect 101829 48113 101885 48169
rect 101885 48113 101889 48169
rect 101825 48109 101889 48113
rect 101905 48169 101969 48173
rect 101905 48113 101909 48169
rect 101909 48113 101965 48169
rect 101965 48113 101969 48169
rect 101905 48109 101969 48113
rect 101985 48169 102049 48173
rect 101985 48113 101989 48169
rect 101989 48113 102045 48169
rect 102045 48113 102049 48169
rect 101985 48109 102049 48113
rect 102065 48169 102129 48173
rect 102065 48113 102069 48169
rect 102069 48113 102125 48169
rect 102125 48113 102129 48169
rect 102065 48109 102129 48113
rect 102145 48169 102209 48173
rect 102145 48113 102149 48169
rect 102149 48113 102205 48169
rect 102205 48113 102209 48169
rect 102145 48109 102209 48113
rect 102225 48169 102289 48173
rect 102225 48113 102229 48169
rect 102229 48113 102285 48169
rect 102285 48113 102289 48169
rect 102225 48109 102289 48113
rect 102305 48169 102369 48173
rect 102305 48113 102309 48169
rect 102309 48113 102365 48169
rect 102365 48113 102369 48169
rect 102305 48109 102369 48113
rect 102385 48169 102449 48173
rect 102385 48113 102389 48169
rect 102389 48113 102445 48169
rect 102445 48113 102449 48169
rect 102385 48109 102449 48113
rect 102465 48169 102529 48173
rect 102465 48113 102469 48169
rect 102469 48113 102525 48169
rect 102525 48113 102529 48169
rect 102465 48109 102529 48113
rect 102545 48169 102609 48173
rect 102545 48113 102549 48169
rect 102549 48113 102605 48169
rect 102605 48113 102609 48169
rect 102545 48109 102609 48113
rect 102625 48169 102689 48173
rect 102625 48113 102629 48169
rect 102629 48113 102685 48169
rect 102685 48113 102689 48169
rect 102625 48109 102689 48113
rect 102705 48169 102769 48173
rect 102705 48113 102709 48169
rect 102709 48113 102765 48169
rect 102765 48113 102769 48169
rect 102705 48109 102769 48113
rect 102785 48169 102849 48173
rect 102785 48113 102789 48169
rect 102789 48113 102845 48169
rect 102845 48113 102849 48169
rect 102785 48109 102849 48113
rect 102865 48169 102929 48173
rect 102865 48113 102869 48169
rect 102869 48113 102925 48169
rect 102925 48113 102929 48169
rect 102865 48109 102929 48113
rect 102945 48169 103009 48173
rect 102945 48113 102949 48169
rect 102949 48113 103005 48169
rect 103005 48113 103009 48169
rect 102945 48109 103009 48113
rect 103025 48169 103089 48173
rect 103025 48113 103029 48169
rect 103029 48113 103085 48169
rect 103085 48113 103089 48169
rect 103025 48109 103089 48113
rect 103105 48169 103169 48173
rect 103105 48113 103109 48169
rect 103109 48113 103165 48169
rect 103165 48113 103169 48169
rect 103105 48109 103169 48113
rect 103185 48169 103249 48173
rect 103185 48113 103189 48169
rect 103189 48113 103245 48169
rect 103245 48113 103249 48169
rect 103185 48109 103249 48113
rect 93160 48036 93224 48040
rect 93160 47980 93164 48036
rect 93164 47980 93220 48036
rect 93220 47980 93224 48036
rect 93160 47976 93224 47980
rect 92246 47884 92310 47888
rect 92246 47828 92250 47884
rect 92250 47828 92306 47884
rect 92306 47828 92310 47884
rect 92246 47824 92310 47828
rect 94917 47601 94981 47605
rect 94917 47545 94921 47601
rect 94921 47545 94977 47601
rect 94977 47545 94981 47601
rect 94917 47541 94981 47545
rect 96445 47677 96449 47697
rect 96449 47677 96505 47697
rect 96505 47677 96509 47697
rect 96445 47653 96509 47677
rect 96445 47633 96449 47653
rect 96449 47633 96505 47653
rect 96505 47633 96509 47653
rect 96445 47597 96449 47617
rect 96449 47597 96505 47617
rect 96505 47597 96509 47617
rect 96445 47573 96509 47597
rect 96445 47553 96449 47573
rect 96449 47553 96505 47573
rect 96505 47553 96509 47573
rect 44708 47197 44772 47201
rect 44708 47141 44712 47197
rect 44712 47141 44768 47197
rect 44768 47141 44772 47197
rect 44708 47137 44772 47141
rect 44708 47117 44772 47121
rect 44708 47061 44712 47117
rect 44712 47061 44768 47117
rect 44768 47061 44772 47117
rect 44708 47057 44772 47061
rect 44708 47037 44772 47041
rect 44708 46981 44712 47037
rect 44712 46981 44768 47037
rect 44768 46981 44772 47037
rect 44708 46977 44772 46981
rect 44708 46957 44772 46961
rect 44708 46901 44712 46957
rect 44712 46901 44768 46957
rect 44768 46901 44772 46957
rect 44708 46897 44772 46901
rect 61913 46949 62297 47173
rect 69682 47168 69746 47232
rect 84205 47168 84269 47232
rect 94924 47200 94988 47204
rect 94924 47144 94928 47200
rect 94928 47144 94984 47200
rect 94984 47144 94988 47200
rect 94924 47140 94988 47144
rect 62812 47021 62876 47085
rect 94924 47120 94988 47124
rect 94924 47064 94928 47120
rect 94928 47064 94984 47120
rect 94984 47064 94988 47120
rect 94924 47060 94988 47064
rect 94924 47040 94988 47044
rect 94924 46984 94928 47040
rect 94928 46984 94984 47040
rect 94984 46984 94988 47040
rect 94924 46980 94988 46984
rect 96440 47206 96504 47210
rect 96440 47150 96444 47206
rect 96444 47150 96500 47206
rect 96500 47150 96504 47206
rect 96440 47146 96504 47150
rect 96440 47126 96504 47130
rect 96440 47070 96444 47126
rect 96444 47070 96500 47126
rect 96500 47070 96504 47126
rect 96440 47066 96504 47070
rect 96440 47046 96504 47050
rect 96440 46990 96444 47046
rect 96444 46990 96500 47046
rect 96500 46990 96504 47046
rect 96440 46986 96504 46990
rect 68570 46873 68634 46937
rect 68931 46874 68995 46938
rect 40495 46682 40559 46746
rect 65223 46682 65287 46746
rect 44705 46641 44769 46645
rect 44705 46585 44709 46641
rect 44709 46585 44765 46641
rect 44765 46585 44769 46641
rect 44705 46581 44769 46585
rect 44705 46561 44769 46565
rect 44705 46505 44709 46561
rect 44709 46505 44765 46561
rect 44765 46505 44769 46561
rect 44705 46501 44769 46505
rect 44705 46481 44769 46485
rect 44705 46425 44709 46481
rect 44709 46425 44765 46481
rect 44765 46425 44769 46481
rect 44705 46421 44769 46425
rect 64695 46231 64759 46295
rect 94017 46607 94241 46831
rect 96445 46351 96449 46371
rect 96449 46351 96505 46371
rect 96505 46351 96509 46371
rect 96445 46327 96509 46351
rect 96445 46307 96449 46327
rect 96449 46307 96505 46327
rect 96505 46307 96509 46327
rect 94923 46265 94987 46269
rect 94923 46209 94927 46265
rect 94927 46209 94983 46265
rect 94983 46209 94987 46265
rect 94923 46205 94987 46209
rect 96445 46271 96449 46291
rect 96449 46271 96505 46291
rect 96505 46271 96509 46291
rect 96445 46247 96509 46271
rect 96445 46227 96449 46247
rect 96449 46227 96505 46247
rect 96505 46227 96509 46247
rect 94918 45812 94982 45816
rect 94918 45756 94922 45812
rect 94922 45756 94978 45812
rect 94978 45756 94982 45812
rect 94918 45752 94982 45756
rect 69166 45613 69230 45677
rect 84751 45613 84815 45677
rect 94918 45732 94982 45736
rect 94918 45676 94922 45732
rect 94922 45676 94978 45732
rect 94978 45676 94982 45732
rect 94918 45672 94982 45676
rect 96446 45840 96510 45844
rect 96446 45784 96450 45840
rect 96450 45784 96506 45840
rect 96506 45784 96510 45840
rect 96446 45780 96510 45784
rect 96446 45760 96510 45764
rect 96446 45704 96450 45760
rect 96450 45704 96506 45760
rect 96506 45704 96510 45760
rect 96446 45700 96510 45704
rect 92246 45603 92310 45607
rect 92246 45547 92250 45603
rect 92250 45547 92306 45603
rect 92306 45547 92310 45603
rect 92246 45543 92310 45547
rect 96446 45680 96510 45684
rect 96446 45624 96450 45680
rect 96450 45624 96506 45680
rect 96506 45624 96510 45680
rect 96446 45620 96510 45624
rect 92571 45397 92635 45401
rect 92571 45341 92575 45397
rect 92575 45341 92631 45397
rect 92631 45341 92635 45397
rect 92571 45337 92635 45341
rect 99983 45173 100047 45177
rect 99983 45117 99987 45173
rect 99987 45117 100043 45173
rect 100043 45117 100047 45173
rect 99983 45113 100047 45117
rect 100063 45173 100127 45177
rect 100063 45117 100067 45173
rect 100067 45117 100123 45173
rect 100123 45117 100127 45173
rect 100063 45113 100127 45117
rect 100143 45173 100207 45177
rect 100143 45117 100147 45173
rect 100147 45117 100203 45173
rect 100203 45117 100207 45173
rect 100143 45113 100207 45117
rect 100223 45173 100287 45177
rect 100223 45117 100227 45173
rect 100227 45117 100283 45173
rect 100283 45117 100287 45173
rect 100223 45113 100287 45117
rect 100303 45173 100367 45177
rect 100303 45117 100307 45173
rect 100307 45117 100363 45173
rect 100363 45117 100367 45173
rect 100303 45113 100367 45117
rect 100383 45173 100447 45177
rect 100383 45117 100387 45173
rect 100387 45117 100443 45173
rect 100443 45117 100447 45173
rect 100383 45113 100447 45117
rect 100463 45173 100527 45177
rect 100463 45117 100467 45173
rect 100467 45117 100523 45173
rect 100523 45117 100527 45173
rect 100463 45113 100527 45117
rect 100543 45173 100607 45177
rect 100543 45117 100547 45173
rect 100547 45117 100603 45173
rect 100603 45117 100607 45173
rect 100543 45113 100607 45117
rect 100623 45173 100687 45177
rect 100623 45117 100627 45173
rect 100627 45117 100683 45173
rect 100683 45117 100687 45173
rect 100623 45113 100687 45117
rect 100703 45173 100767 45177
rect 100703 45117 100707 45173
rect 100707 45117 100763 45173
rect 100763 45117 100767 45173
rect 100703 45113 100767 45117
rect 100783 45173 100847 45177
rect 100783 45117 100787 45173
rect 100787 45117 100843 45173
rect 100843 45117 100847 45173
rect 100783 45113 100847 45117
rect 100863 45173 100927 45177
rect 100863 45117 100867 45173
rect 100867 45117 100923 45173
rect 100923 45117 100927 45173
rect 100863 45113 100927 45117
rect 100943 45173 101007 45177
rect 100943 45117 100947 45173
rect 100947 45117 101003 45173
rect 101003 45117 101007 45173
rect 100943 45113 101007 45117
rect 101023 45173 101087 45177
rect 101023 45117 101027 45173
rect 101027 45117 101083 45173
rect 101083 45117 101087 45173
rect 101023 45113 101087 45117
rect 101103 45173 101167 45177
rect 101103 45117 101107 45173
rect 101107 45117 101163 45173
rect 101163 45117 101167 45173
rect 101103 45113 101167 45117
rect 101183 45173 101247 45177
rect 101183 45117 101187 45173
rect 101187 45117 101243 45173
rect 101243 45117 101247 45173
rect 101183 45113 101247 45117
rect 101263 45173 101327 45177
rect 101263 45117 101267 45173
rect 101267 45117 101323 45173
rect 101323 45117 101327 45173
rect 101263 45113 101327 45117
rect 101343 45173 101407 45177
rect 101343 45117 101347 45173
rect 101347 45117 101403 45173
rect 101403 45117 101407 45173
rect 101343 45113 101407 45117
rect 101423 45173 101487 45177
rect 101423 45117 101427 45173
rect 101427 45117 101483 45173
rect 101483 45117 101487 45173
rect 101423 45113 101487 45117
rect 101503 45173 101567 45177
rect 101503 45117 101507 45173
rect 101507 45117 101563 45173
rect 101563 45117 101567 45173
rect 101503 45113 101567 45117
rect 101583 45173 101647 45177
rect 101583 45117 101587 45173
rect 101587 45117 101643 45173
rect 101643 45117 101647 45173
rect 101583 45113 101647 45117
rect 101663 45173 101727 45177
rect 101663 45117 101667 45173
rect 101667 45117 101723 45173
rect 101723 45117 101727 45173
rect 101663 45113 101727 45117
rect 101743 45173 101807 45177
rect 101743 45117 101747 45173
rect 101747 45117 101803 45173
rect 101803 45117 101807 45173
rect 101743 45113 101807 45117
rect 101823 45173 101887 45177
rect 101823 45117 101827 45173
rect 101827 45117 101883 45173
rect 101883 45117 101887 45173
rect 101823 45113 101887 45117
rect 101903 45173 101967 45177
rect 101903 45117 101907 45173
rect 101907 45117 101963 45173
rect 101963 45117 101967 45173
rect 101903 45113 101967 45117
rect 101983 45173 102047 45177
rect 101983 45117 101987 45173
rect 101987 45117 102043 45173
rect 102043 45117 102047 45173
rect 101983 45113 102047 45117
rect 102063 45173 102127 45177
rect 102063 45117 102067 45173
rect 102067 45117 102123 45173
rect 102123 45117 102127 45173
rect 102063 45113 102127 45117
rect 102143 45173 102207 45177
rect 102143 45117 102147 45173
rect 102147 45117 102203 45173
rect 102203 45117 102207 45173
rect 102143 45113 102207 45117
rect 102223 45173 102287 45177
rect 102223 45117 102227 45173
rect 102227 45117 102283 45173
rect 102283 45117 102287 45173
rect 102223 45113 102287 45117
rect 102303 45173 102367 45177
rect 102303 45117 102307 45173
rect 102307 45117 102363 45173
rect 102363 45117 102367 45173
rect 102303 45113 102367 45117
rect 102383 45173 102447 45177
rect 102383 45117 102387 45173
rect 102387 45117 102443 45173
rect 102443 45117 102447 45173
rect 102383 45113 102447 45117
rect 102463 45173 102527 45177
rect 102463 45117 102467 45173
rect 102467 45117 102523 45173
rect 102523 45117 102527 45173
rect 102463 45113 102527 45117
rect 102543 45173 102607 45177
rect 102543 45117 102547 45173
rect 102547 45117 102603 45173
rect 102603 45117 102607 45173
rect 102543 45113 102607 45117
rect 102623 45173 102687 45177
rect 102623 45117 102627 45173
rect 102627 45117 102683 45173
rect 102683 45117 102687 45173
rect 102623 45113 102687 45117
rect 102703 45173 102767 45177
rect 102703 45117 102707 45173
rect 102707 45117 102763 45173
rect 102763 45117 102767 45173
rect 102703 45113 102767 45117
rect 102783 45173 102847 45177
rect 102783 45117 102787 45173
rect 102787 45117 102843 45173
rect 102843 45117 102847 45173
rect 102783 45113 102847 45117
rect 102863 45173 102927 45177
rect 102863 45117 102867 45173
rect 102867 45117 102923 45173
rect 102923 45117 102927 45173
rect 102863 45113 102927 45117
rect 102943 45173 103007 45177
rect 102943 45117 102947 45173
rect 102947 45117 103003 45173
rect 103003 45117 103007 45173
rect 102943 45113 103007 45117
rect 103023 45173 103087 45177
rect 103023 45117 103027 45173
rect 103027 45117 103083 45173
rect 103083 45117 103087 45173
rect 103023 45113 103087 45117
rect 103103 45173 103167 45177
rect 103103 45117 103107 45173
rect 103107 45117 103163 45173
rect 103163 45117 103167 45173
rect 103103 45113 103167 45117
rect 103183 45173 103247 45177
rect 103183 45117 103187 45173
rect 103187 45117 103243 45173
rect 103243 45117 103247 45173
rect 103183 45113 103247 45117
rect 18947 43076 19011 43080
rect 18947 43020 18951 43076
rect 18951 43020 19007 43076
rect 19007 43020 19011 43076
rect 18947 43016 19011 43020
rect 19027 43076 19091 43080
rect 19027 43020 19031 43076
rect 19031 43020 19087 43076
rect 19087 43020 19091 43076
rect 19027 43016 19091 43020
rect 19107 43076 19171 43080
rect 19107 43020 19111 43076
rect 19111 43020 19167 43076
rect 19167 43020 19171 43076
rect 19107 43016 19171 43020
rect 19187 43076 19251 43080
rect 19187 43020 19191 43076
rect 19191 43020 19247 43076
rect 19247 43020 19251 43076
rect 19187 43016 19251 43020
rect 19267 43076 19331 43080
rect 19267 43020 19271 43076
rect 19271 43020 19327 43076
rect 19327 43020 19331 43076
rect 19267 43016 19331 43020
rect 19347 43076 19411 43080
rect 19347 43020 19351 43076
rect 19351 43020 19407 43076
rect 19407 43020 19411 43076
rect 19347 43016 19411 43020
rect 19427 43076 19491 43080
rect 19427 43020 19431 43076
rect 19431 43020 19487 43076
rect 19487 43020 19491 43076
rect 19427 43016 19491 43020
rect 19507 43076 19571 43080
rect 19507 43020 19511 43076
rect 19511 43020 19567 43076
rect 19567 43020 19571 43076
rect 19507 43016 19571 43020
rect 19587 43076 19651 43080
rect 19587 43020 19591 43076
rect 19591 43020 19647 43076
rect 19647 43020 19651 43076
rect 19587 43016 19651 43020
rect 19667 43076 19731 43080
rect 19667 43020 19671 43076
rect 19671 43020 19727 43076
rect 19727 43020 19731 43076
rect 19667 43016 19731 43020
rect 19747 43076 19811 43080
rect 19747 43020 19751 43076
rect 19751 43020 19807 43076
rect 19807 43020 19811 43076
rect 19747 43016 19811 43020
rect 19827 43076 19891 43080
rect 19827 43020 19831 43076
rect 19831 43020 19887 43076
rect 19887 43020 19891 43076
rect 19827 43016 19891 43020
rect 19907 43076 19971 43080
rect 19907 43020 19911 43076
rect 19911 43020 19967 43076
rect 19967 43020 19971 43076
rect 19907 43016 19971 43020
rect 19987 43076 20051 43080
rect 19987 43020 19991 43076
rect 19991 43020 20047 43076
rect 20047 43020 20051 43076
rect 19987 43016 20051 43020
rect 20067 43076 20131 43080
rect 20067 43020 20071 43076
rect 20071 43020 20127 43076
rect 20127 43020 20131 43076
rect 20067 43016 20131 43020
rect 20147 43076 20211 43080
rect 20147 43020 20151 43076
rect 20151 43020 20207 43076
rect 20207 43020 20211 43076
rect 20147 43016 20211 43020
rect 20227 43076 20291 43080
rect 20227 43020 20231 43076
rect 20231 43020 20287 43076
rect 20287 43020 20291 43076
rect 20227 43016 20291 43020
rect 20307 43076 20371 43080
rect 20307 43020 20311 43076
rect 20311 43020 20367 43076
rect 20367 43020 20371 43076
rect 20307 43016 20371 43020
rect 20387 43076 20451 43080
rect 20387 43020 20391 43076
rect 20391 43020 20447 43076
rect 20447 43020 20451 43076
rect 20387 43016 20451 43020
rect 20467 43076 20531 43080
rect 20467 43020 20471 43076
rect 20471 43020 20527 43076
rect 20527 43020 20531 43076
rect 20467 43016 20531 43020
rect 20547 43076 20611 43080
rect 20547 43020 20551 43076
rect 20551 43020 20607 43076
rect 20607 43020 20611 43076
rect 20547 43016 20611 43020
rect 20627 43076 20691 43080
rect 20627 43020 20631 43076
rect 20631 43020 20687 43076
rect 20687 43020 20691 43076
rect 20627 43016 20691 43020
rect 20707 43076 20771 43080
rect 20707 43020 20711 43076
rect 20711 43020 20767 43076
rect 20767 43020 20771 43076
rect 20707 43016 20771 43020
rect 20787 43076 20851 43080
rect 20787 43020 20791 43076
rect 20791 43020 20847 43076
rect 20847 43020 20851 43076
rect 20787 43016 20851 43020
rect 20867 43076 20931 43080
rect 20867 43020 20871 43076
rect 20871 43020 20927 43076
rect 20927 43020 20931 43076
rect 20867 43016 20931 43020
rect 20947 43076 21011 43080
rect 20947 43020 20951 43076
rect 20951 43020 21007 43076
rect 21007 43020 21011 43076
rect 20947 43016 21011 43020
rect 21027 43076 21091 43080
rect 21027 43020 21031 43076
rect 21031 43020 21087 43076
rect 21087 43020 21091 43076
rect 21027 43016 21091 43020
rect 21107 43076 21171 43080
rect 21107 43020 21111 43076
rect 21111 43020 21167 43076
rect 21167 43020 21171 43076
rect 21107 43016 21171 43020
rect 21187 43076 21251 43080
rect 21187 43020 21191 43076
rect 21191 43020 21247 43076
rect 21247 43020 21251 43076
rect 21187 43016 21251 43020
rect 21267 43076 21331 43080
rect 21267 43020 21271 43076
rect 21271 43020 21327 43076
rect 21327 43020 21331 43076
rect 21267 43016 21331 43020
rect 21347 43076 21411 43080
rect 21347 43020 21351 43076
rect 21351 43020 21407 43076
rect 21407 43020 21411 43076
rect 21347 43016 21411 43020
rect 21427 43076 21491 43080
rect 21427 43020 21431 43076
rect 21431 43020 21487 43076
rect 21487 43020 21491 43076
rect 21427 43016 21491 43020
rect 21507 43076 21571 43080
rect 21507 43020 21511 43076
rect 21511 43020 21567 43076
rect 21567 43020 21571 43076
rect 21507 43016 21571 43020
rect 21587 43076 21651 43080
rect 21587 43020 21591 43076
rect 21591 43020 21647 43076
rect 21647 43020 21651 43076
rect 21587 43016 21651 43020
rect 21667 43076 21731 43080
rect 21667 43020 21671 43076
rect 21671 43020 21727 43076
rect 21727 43020 21731 43076
rect 21667 43016 21731 43020
rect 21747 43076 21811 43080
rect 21747 43020 21751 43076
rect 21751 43020 21807 43076
rect 21807 43020 21811 43076
rect 21747 43016 21811 43020
rect 21827 43076 21891 43080
rect 21827 43020 21831 43076
rect 21831 43020 21887 43076
rect 21887 43020 21891 43076
rect 21827 43016 21891 43020
rect 21907 43076 21971 43080
rect 21907 43020 21911 43076
rect 21911 43020 21967 43076
rect 21967 43020 21971 43076
rect 21907 43016 21971 43020
rect 21987 43076 22051 43080
rect 21987 43020 21991 43076
rect 21991 43020 22047 43076
rect 22047 43020 22051 43076
rect 21987 43016 22051 43020
rect 22067 43076 22131 43080
rect 22067 43020 22071 43076
rect 22071 43020 22127 43076
rect 22127 43020 22131 43076
rect 22067 43016 22131 43020
rect 22147 43076 22211 43080
rect 22147 43020 22151 43076
rect 22151 43020 22207 43076
rect 22207 43020 22211 43076
rect 22147 43016 22211 43020
rect 18949 40081 19013 40085
rect 18949 40025 18953 40081
rect 18953 40025 19009 40081
rect 19009 40025 19013 40081
rect 18949 40021 19013 40025
rect 19029 40081 19093 40085
rect 19029 40025 19033 40081
rect 19033 40025 19089 40081
rect 19089 40025 19093 40081
rect 19029 40021 19093 40025
rect 19109 40081 19173 40085
rect 19109 40025 19113 40081
rect 19113 40025 19169 40081
rect 19169 40025 19173 40081
rect 19109 40021 19173 40025
rect 19189 40081 19253 40085
rect 19189 40025 19193 40081
rect 19193 40025 19249 40081
rect 19249 40025 19253 40081
rect 19189 40021 19253 40025
rect 19269 40081 19333 40085
rect 19269 40025 19273 40081
rect 19273 40025 19329 40081
rect 19329 40025 19333 40081
rect 19269 40021 19333 40025
rect 19349 40081 19413 40085
rect 19349 40025 19353 40081
rect 19353 40025 19409 40081
rect 19409 40025 19413 40081
rect 19349 40021 19413 40025
rect 19429 40081 19493 40085
rect 19429 40025 19433 40081
rect 19433 40025 19489 40081
rect 19489 40025 19493 40081
rect 19429 40021 19493 40025
rect 19509 40081 19573 40085
rect 19509 40025 19513 40081
rect 19513 40025 19569 40081
rect 19569 40025 19573 40081
rect 19509 40021 19573 40025
rect 19589 40081 19653 40085
rect 19589 40025 19593 40081
rect 19593 40025 19649 40081
rect 19649 40025 19653 40081
rect 19589 40021 19653 40025
rect 19669 40081 19733 40085
rect 19669 40025 19673 40081
rect 19673 40025 19729 40081
rect 19729 40025 19733 40081
rect 19669 40021 19733 40025
rect 19749 40081 19813 40085
rect 19749 40025 19753 40081
rect 19753 40025 19809 40081
rect 19809 40025 19813 40081
rect 19749 40021 19813 40025
rect 19829 40081 19893 40085
rect 19829 40025 19833 40081
rect 19833 40025 19889 40081
rect 19889 40025 19893 40081
rect 19829 40021 19893 40025
rect 19909 40081 19973 40085
rect 19909 40025 19913 40081
rect 19913 40025 19969 40081
rect 19969 40025 19973 40081
rect 19909 40021 19973 40025
rect 19989 40081 20053 40085
rect 19989 40025 19993 40081
rect 19993 40025 20049 40081
rect 20049 40025 20053 40081
rect 19989 40021 20053 40025
rect 20069 40081 20133 40085
rect 20069 40025 20073 40081
rect 20073 40025 20129 40081
rect 20129 40025 20133 40081
rect 20069 40021 20133 40025
rect 20149 40081 20213 40085
rect 20149 40025 20153 40081
rect 20153 40025 20209 40081
rect 20209 40025 20213 40081
rect 20149 40021 20213 40025
rect 20229 40081 20293 40085
rect 20229 40025 20233 40081
rect 20233 40025 20289 40081
rect 20289 40025 20293 40081
rect 20229 40021 20293 40025
rect 20309 40081 20373 40085
rect 20309 40025 20313 40081
rect 20313 40025 20369 40081
rect 20369 40025 20373 40081
rect 20309 40021 20373 40025
rect 20389 40081 20453 40085
rect 20389 40025 20393 40081
rect 20393 40025 20449 40081
rect 20449 40025 20453 40081
rect 20389 40021 20453 40025
rect 20469 40081 20533 40085
rect 20469 40025 20473 40081
rect 20473 40025 20529 40081
rect 20529 40025 20533 40081
rect 20469 40021 20533 40025
rect 20549 40081 20613 40085
rect 20549 40025 20553 40081
rect 20553 40025 20609 40081
rect 20609 40025 20613 40081
rect 20549 40021 20613 40025
rect 20629 40081 20693 40085
rect 20629 40025 20633 40081
rect 20633 40025 20689 40081
rect 20689 40025 20693 40081
rect 20629 40021 20693 40025
rect 20709 40081 20773 40085
rect 20709 40025 20713 40081
rect 20713 40025 20769 40081
rect 20769 40025 20773 40081
rect 20709 40021 20773 40025
rect 20789 40081 20853 40085
rect 20789 40025 20793 40081
rect 20793 40025 20849 40081
rect 20849 40025 20853 40081
rect 20789 40021 20853 40025
rect 20869 40081 20933 40085
rect 20869 40025 20873 40081
rect 20873 40025 20929 40081
rect 20929 40025 20933 40081
rect 20869 40021 20933 40025
rect 20949 40081 21013 40085
rect 20949 40025 20953 40081
rect 20953 40025 21009 40081
rect 21009 40025 21013 40081
rect 20949 40021 21013 40025
rect 21029 40081 21093 40085
rect 21029 40025 21033 40081
rect 21033 40025 21089 40081
rect 21089 40025 21093 40081
rect 21029 40021 21093 40025
rect 21109 40081 21173 40085
rect 21109 40025 21113 40081
rect 21113 40025 21169 40081
rect 21169 40025 21173 40081
rect 21109 40021 21173 40025
rect 21189 40081 21253 40085
rect 21189 40025 21193 40081
rect 21193 40025 21249 40081
rect 21249 40025 21253 40081
rect 21189 40021 21253 40025
rect 21269 40081 21333 40085
rect 21269 40025 21273 40081
rect 21273 40025 21329 40081
rect 21329 40025 21333 40081
rect 21269 40021 21333 40025
rect 21349 40081 21413 40085
rect 21349 40025 21353 40081
rect 21353 40025 21409 40081
rect 21409 40025 21413 40081
rect 21349 40021 21413 40025
rect 21429 40081 21493 40085
rect 21429 40025 21433 40081
rect 21433 40025 21489 40081
rect 21489 40025 21493 40081
rect 21429 40021 21493 40025
rect 21509 40081 21573 40085
rect 21509 40025 21513 40081
rect 21513 40025 21569 40081
rect 21569 40025 21573 40081
rect 21509 40021 21573 40025
rect 21589 40081 21653 40085
rect 21589 40025 21593 40081
rect 21593 40025 21649 40081
rect 21649 40025 21653 40081
rect 21589 40021 21653 40025
rect 21669 40081 21733 40085
rect 21669 40025 21673 40081
rect 21673 40025 21729 40081
rect 21729 40025 21733 40081
rect 21669 40021 21733 40025
rect 21749 40081 21813 40085
rect 21749 40025 21753 40081
rect 21753 40025 21809 40081
rect 21809 40025 21813 40081
rect 21749 40021 21813 40025
rect 21829 40081 21893 40085
rect 21829 40025 21833 40081
rect 21833 40025 21889 40081
rect 21889 40025 21893 40081
rect 21829 40021 21893 40025
rect 21909 40081 21973 40085
rect 21909 40025 21913 40081
rect 21913 40025 21969 40081
rect 21969 40025 21973 40081
rect 21909 40021 21973 40025
rect 21989 40081 22053 40085
rect 21989 40025 21993 40081
rect 21993 40025 22049 40081
rect 22049 40025 22053 40081
rect 21989 40021 22053 40025
rect 22069 40081 22133 40085
rect 22069 40025 22073 40081
rect 22073 40025 22129 40081
rect 22129 40025 22133 40081
rect 22069 40021 22133 40025
rect 22149 40081 22213 40085
rect 22149 40025 22153 40081
rect 22153 40025 22209 40081
rect 22209 40025 22213 40081
rect 22149 40021 22213 40025
rect 70030 44985 70094 45049
rect 31642 41904 31706 41908
rect 31642 41848 31646 41904
rect 31646 41848 31702 41904
rect 31702 41848 31706 41904
rect 31642 41844 31706 41848
rect 31642 41824 31706 41828
rect 31642 41768 31646 41824
rect 31646 41768 31702 41824
rect 31702 41768 31706 41824
rect 31642 41764 31706 41768
rect 31642 41744 31706 41748
rect 31642 41688 31646 41744
rect 31646 41688 31702 41744
rect 31702 41688 31706 41744
rect 31642 41684 31706 41688
rect 31648 41416 31712 41420
rect 31648 41360 31652 41416
rect 31652 41360 31708 41416
rect 31708 41360 31712 41416
rect 31648 41356 31712 41360
rect 31648 41336 31712 41340
rect 31648 41280 31652 41336
rect 31652 41280 31708 41336
rect 31708 41280 31712 41336
rect 31648 41276 31712 41280
rect 31648 41256 31712 41260
rect 31648 41200 31652 41256
rect 31652 41200 31708 41256
rect 31708 41200 31712 41256
rect 31648 41196 31712 41200
rect 40495 44609 40559 44673
rect 68174 44292 68238 44356
rect 46678 41175 46742 41179
rect 46678 41119 46682 41175
rect 46682 41119 46738 41175
rect 46738 41119 46742 41175
rect 46678 41115 46742 41119
rect 42942 39388 43006 39392
rect 42942 39332 42946 39388
rect 42946 39332 43002 39388
rect 43002 39332 43006 39388
rect 42942 39328 43006 39332
rect 31581 38431 31645 38435
rect 31581 38375 31585 38431
rect 31585 38375 31641 38431
rect 31641 38375 31645 38431
rect 31581 38371 31645 38375
rect 31581 38351 31645 38355
rect 31581 38295 31585 38351
rect 31585 38295 31641 38351
rect 31641 38295 31645 38351
rect 31581 38291 31645 38295
rect 31581 38271 31645 38275
rect 31581 38215 31585 38271
rect 31585 38215 31641 38271
rect 31641 38215 31645 38271
rect 31581 38211 31645 38215
rect 38871 38091 38935 38095
rect 38871 38035 38875 38091
rect 38875 38035 38931 38091
rect 38931 38035 38935 38091
rect 38871 38031 38935 38035
rect 31580 37937 31644 37941
rect 31580 37881 31584 37937
rect 31584 37881 31640 37937
rect 31640 37881 31644 37937
rect 31580 37877 31644 37881
rect 31580 37857 31644 37861
rect 31580 37801 31584 37857
rect 31584 37801 31640 37857
rect 31640 37801 31644 37857
rect 31580 37797 31644 37801
rect 31580 37777 31644 37781
rect 31580 37721 31584 37777
rect 31584 37721 31640 37777
rect 31640 37721 31644 37777
rect 31580 37717 31644 37721
rect 46124 34241 46188 34245
rect 46124 34185 46128 34241
rect 46128 34185 46184 34241
rect 46184 34185 46188 34241
rect 46124 34181 46188 34185
rect 68570 43761 68634 43825
rect 54279 43471 54343 43535
rect 51815 43001 51879 43065
rect 53176 43001 53240 43065
rect 51308 39726 51372 39730
rect 51308 39670 51312 39726
rect 51312 39670 51368 39726
rect 51368 39670 51372 39726
rect 51308 39666 51372 39670
rect 52195 38431 52259 38435
rect 52195 38375 52199 38431
rect 52199 38375 52255 38431
rect 52255 38375 52259 38431
rect 52195 38371 52259 38375
rect 52195 38351 52259 38355
rect 52195 38295 52199 38351
rect 52199 38295 52255 38351
rect 52255 38295 52259 38351
rect 52195 38291 52259 38295
rect 50932 34845 50996 34849
rect 50932 34789 50936 34845
rect 50936 34789 50992 34845
rect 50992 34789 50996 34845
rect 50932 34785 50996 34789
rect 51012 34845 51076 34849
rect 51012 34789 51016 34845
rect 51016 34789 51072 34845
rect 51072 34789 51076 34845
rect 51012 34785 51076 34789
rect 51092 34845 51156 34849
rect 51092 34789 51096 34845
rect 51096 34789 51152 34845
rect 51152 34789 51156 34845
rect 51092 34785 51156 34789
rect 50934 33602 50998 33606
rect 50934 33546 50938 33602
rect 50938 33546 50994 33602
rect 50994 33546 50998 33602
rect 50934 33542 50998 33546
rect 51014 33602 51078 33606
rect 51014 33546 51018 33602
rect 51018 33546 51074 33602
rect 51074 33546 51078 33602
rect 51014 33542 51078 33546
rect 51094 33602 51158 33606
rect 51094 33546 51098 33602
rect 51098 33546 51154 33602
rect 51154 33546 51158 33602
rect 51094 33542 51158 33546
rect 71781 43345 71845 43349
rect 71781 43289 71785 43345
rect 71785 43289 71841 43345
rect 71841 43289 71845 43345
rect 71781 43285 71845 43289
rect 80783 43400 80847 43404
rect 80783 43344 80787 43400
rect 80787 43344 80843 43400
rect 80843 43344 80847 43400
rect 80783 43340 80847 43344
rect 54696 43170 54760 43234
rect 61967 43190 62271 43194
rect 61967 43054 61971 43190
rect 61971 43054 62267 43190
rect 62267 43054 62271 43190
rect 61967 43050 62271 43054
rect 67326 43076 67390 43080
rect 67326 43020 67330 43076
rect 67330 43020 67386 43076
rect 67386 43020 67390 43076
rect 67326 43016 67390 43020
rect 78065 43080 78129 43084
rect 78065 43024 78069 43080
rect 78069 43024 78125 43080
rect 78125 43024 78129 43080
rect 78065 43020 78129 43024
rect 55590 42868 55654 42932
rect 55961 42609 56025 42673
rect 65374 42736 65438 42740
rect 65374 42680 65378 42736
rect 65378 42680 65434 42736
rect 65434 42680 65438 42736
rect 65374 42676 65438 42680
rect 70024 42646 70088 42710
rect 71209 42529 71273 42593
rect 82708 42529 82772 42593
rect 56414 42270 56478 42334
rect 56810 41989 56874 42053
rect 53922 41654 54306 41878
rect 71462 41721 71526 41785
rect 82455 41722 82519 41786
rect 58075 41483 58139 41547
rect 71783 41560 71847 41564
rect 71783 41504 71787 41560
rect 71787 41504 71843 41560
rect 71843 41504 71847 41560
rect 71783 41500 71847 41504
rect 80783 41570 80847 41574
rect 80783 41514 80787 41570
rect 80787 41514 80843 41570
rect 80843 41514 80847 41570
rect 80783 41510 80847 41514
rect 61389 41307 61453 41311
rect 61389 41251 61393 41307
rect 61393 41251 61449 41307
rect 61449 41251 61453 41307
rect 61389 41247 61453 41251
rect 63321 41307 63385 41311
rect 63321 41251 63325 41307
rect 63325 41251 63381 41307
rect 63381 41251 63385 41307
rect 63321 41247 63385 41251
rect 70050 41041 70114 41105
rect 57357 40432 68221 40436
rect 57357 40296 57361 40432
rect 57361 40296 68217 40432
rect 68217 40296 68221 40432
rect 57357 40292 68221 40296
rect 53585 40163 53649 40227
rect 53166 39412 53230 39476
rect 53959 38988 54023 38992
rect 53959 38932 53963 38988
rect 53963 38932 54019 38988
rect 54019 38932 54023 38988
rect 53959 38928 54023 38932
rect 53959 38908 54023 38912
rect 53959 38852 53963 38908
rect 53963 38852 54019 38908
rect 54019 38852 54023 38908
rect 53959 38848 54023 38852
rect 53959 38828 54023 38832
rect 53959 38772 53963 38828
rect 53963 38772 54019 38828
rect 54019 38772 54023 38828
rect 53959 38768 54023 38772
rect 53585 38602 53649 38666
rect 53909 32665 53973 32729
rect 40345 31625 40409 31629
rect 40345 31569 40349 31625
rect 40349 31569 40405 31625
rect 40405 31569 40409 31625
rect 40345 31565 40409 31569
rect 55295 37139 55359 37143
rect 55295 37083 55299 37139
rect 55299 37083 55355 37139
rect 55355 37083 55359 37139
rect 55295 37079 55359 37083
rect 55295 37059 55359 37063
rect 55295 37003 55299 37059
rect 55299 37003 55355 37059
rect 55355 37003 55359 37059
rect 55295 36999 55359 37003
rect 55295 36979 55359 36983
rect 55295 36923 55299 36979
rect 55299 36923 55355 36979
rect 55355 36923 55359 36979
rect 55295 36919 55359 36923
rect 55295 36899 55359 36903
rect 55295 36843 55299 36899
rect 55299 36843 55355 36899
rect 55355 36843 55359 36899
rect 55295 36839 55359 36843
rect 55295 36819 55359 36823
rect 55295 36763 55299 36819
rect 55299 36763 55355 36819
rect 55355 36763 55359 36819
rect 55295 36759 55359 36763
rect 55336 35544 55400 35548
rect 55336 35488 55340 35544
rect 55340 35488 55396 35544
rect 55396 35488 55400 35544
rect 55336 35484 55400 35488
rect 55336 35464 55400 35468
rect 55336 35408 55340 35464
rect 55340 35408 55396 35464
rect 55396 35408 55400 35464
rect 55336 35404 55400 35408
rect 55336 35384 55400 35388
rect 55336 35328 55340 35384
rect 55340 35328 55396 35384
rect 55396 35328 55400 35384
rect 55336 35324 55400 35328
rect 55336 35304 55400 35308
rect 55336 35248 55340 35304
rect 55340 35248 55396 35304
rect 55396 35248 55400 35304
rect 55336 35244 55400 35248
rect 55336 35224 55400 35228
rect 55336 35168 55340 35224
rect 55340 35168 55396 35224
rect 55396 35168 55400 35224
rect 55336 35164 55400 35168
rect 49919 31253 50303 31257
rect 49919 31037 50303 31253
rect 49919 31033 50303 31037
rect 31578 30668 31642 30672
rect 31578 30612 31582 30668
rect 31582 30612 31638 30668
rect 31638 30612 31642 30668
rect 31578 30608 31642 30612
rect 31578 30588 31642 30592
rect 31578 30532 31582 30588
rect 31582 30532 31638 30588
rect 31638 30532 31642 30588
rect 31578 30528 31642 30532
rect 31578 30508 31642 30512
rect 31578 30452 31582 30508
rect 31582 30452 31638 30508
rect 31638 30452 31642 30508
rect 31578 30448 31642 30452
rect 53910 30607 53974 30671
rect 38843 30321 38907 30325
rect 38843 30265 38847 30321
rect 38847 30265 38903 30321
rect 38903 30265 38907 30321
rect 38843 30261 38907 30265
rect 31577 30181 31641 30185
rect 31577 30125 31581 30181
rect 31581 30125 31637 30181
rect 31637 30125 31641 30181
rect 31577 30121 31641 30125
rect 31577 30101 31641 30105
rect 31577 30045 31581 30101
rect 31581 30045 31637 30101
rect 31637 30045 31641 30101
rect 31577 30041 31641 30045
rect 31577 30021 31641 30025
rect 31577 29965 31581 30021
rect 31581 29965 31637 30021
rect 31637 29965 31641 30021
rect 31577 29961 31641 29965
rect 52188 30146 52252 30150
rect 52188 30090 52192 30146
rect 52192 30090 52248 30146
rect 52248 30090 52252 30146
rect 52188 30086 52252 30090
rect 52188 30066 52252 30070
rect 52188 30010 52192 30066
rect 52192 30010 52248 30066
rect 52248 30010 52252 30066
rect 52188 30006 52252 30010
rect 53166 30000 53230 30064
rect 53910 29566 53974 29570
rect 53910 29510 53914 29566
rect 53914 29510 53970 29566
rect 53970 29510 53974 29566
rect 53910 29506 53974 29510
rect 53910 29486 53974 29490
rect 53910 29430 53914 29486
rect 53914 29430 53970 29486
rect 53970 29430 53974 29486
rect 53910 29426 53974 29430
rect 53910 29406 53974 29410
rect 53910 29350 53914 29406
rect 53914 29350 53970 29406
rect 53970 29350 53974 29406
rect 53910 29346 53974 29350
rect 53585 29191 53649 29255
rect 55335 33941 55399 33945
rect 55335 33885 55339 33941
rect 55339 33885 55395 33941
rect 55395 33885 55399 33941
rect 55335 33881 55399 33885
rect 55335 33861 55399 33865
rect 55335 33805 55339 33861
rect 55339 33805 55395 33861
rect 55395 33805 55399 33861
rect 55335 33801 55399 33805
rect 55335 33781 55399 33785
rect 55335 33725 55339 33781
rect 55339 33725 55395 33781
rect 55395 33725 55399 33781
rect 55335 33721 55399 33725
rect 55335 33701 55399 33705
rect 55335 33645 55339 33701
rect 55339 33645 55395 33701
rect 55395 33645 55399 33701
rect 55335 33641 55399 33645
rect 55335 33621 55399 33625
rect 55335 33565 55339 33621
rect 55339 33565 55395 33621
rect 55395 33565 55399 33621
rect 55335 33561 55399 33565
rect 71780 39729 71844 39733
rect 71780 39673 71784 39729
rect 71784 39673 71840 39729
rect 71840 39673 71844 39729
rect 71780 39669 71844 39673
rect 80780 39806 80844 39810
rect 80780 39750 80784 39806
rect 80784 39750 80840 39806
rect 80840 39750 80844 39806
rect 80780 39746 80844 39750
rect 78022 39514 78086 39518
rect 78022 39458 78026 39514
rect 78026 39458 78082 39514
rect 78082 39458 78086 39514
rect 78022 39454 78086 39458
rect 70067 39186 70131 39250
rect 71779 37983 71843 37987
rect 71779 37927 71783 37983
rect 71783 37927 71839 37983
rect 71839 37927 71843 37983
rect 71779 37923 71843 37927
rect 80780 38015 80844 38019
rect 80780 37959 80784 38015
rect 80784 37959 80840 38015
rect 80840 37959 80844 38015
rect 80780 37955 80844 37959
rect 70097 37486 70161 37550
rect 71209 37129 71273 37193
rect 71462 36321 71526 36385
rect 71796 36198 71860 36202
rect 71796 36142 71800 36198
rect 71800 36142 71856 36198
rect 71856 36142 71860 36198
rect 71796 36138 71860 36142
rect 80785 36208 80849 36212
rect 80785 36152 80789 36208
rect 80789 36152 80845 36208
rect 80845 36152 80849 36208
rect 80785 36148 80849 36152
rect 78079 35924 78143 35928
rect 78079 35868 78083 35924
rect 78083 35868 78139 35924
rect 78139 35868 78143 35924
rect 78079 35864 78143 35868
rect 70095 35634 70159 35698
rect 63592 34536 68296 34540
rect 63592 34400 63596 34536
rect 63596 34400 68292 34536
rect 68292 34400 68296 34536
rect 63592 34396 68296 34400
rect 71785 34401 71849 34405
rect 71785 34345 71789 34401
rect 71789 34345 71845 34401
rect 71845 34345 71849 34401
rect 71785 34341 71849 34345
rect 80785 34398 80849 34402
rect 80785 34342 80789 34398
rect 80789 34342 80845 34398
rect 80845 34342 80849 34398
rect 80785 34338 80849 34342
rect 93160 33172 93224 33176
rect 93160 33116 93164 33172
rect 93164 33116 93220 33172
rect 93220 33116 93224 33172
rect 93160 33112 93224 33116
rect 55338 32340 55402 32344
rect 55338 32284 55342 32340
rect 55342 32284 55398 32340
rect 55398 32284 55402 32340
rect 55338 32280 55402 32284
rect 55338 32260 55402 32264
rect 55338 32204 55342 32260
rect 55342 32204 55398 32260
rect 55398 32204 55402 32260
rect 55338 32200 55402 32204
rect 55338 32180 55402 32184
rect 55338 32124 55342 32180
rect 55342 32124 55398 32180
rect 55398 32124 55402 32180
rect 55338 32120 55402 32124
rect 55338 32100 55402 32104
rect 55338 32044 55342 32100
rect 55342 32044 55398 32100
rect 55398 32044 55402 32100
rect 55338 32040 55402 32044
rect 55338 32020 55402 32024
rect 55338 31964 55342 32020
rect 55342 31964 55398 32020
rect 55398 31964 55402 32020
rect 55338 31960 55402 31964
rect 94001 32584 94225 32808
rect 92583 32549 92647 32553
rect 92583 32493 92587 32549
rect 92587 32493 92643 32549
rect 92643 32493 92647 32549
rect 92583 32489 92647 32493
rect 93725 32487 93789 32491
rect 93725 32431 93729 32487
rect 93729 32431 93785 32487
rect 93785 32431 93789 32487
rect 93725 32427 93789 32431
rect 92122 31241 92186 31245
rect 92122 31185 92126 31241
rect 92126 31185 92182 31241
rect 92182 31185 92186 31241
rect 95670 31559 95734 31563
rect 95670 31503 95674 31559
rect 95674 31503 95730 31559
rect 95730 31503 95734 31559
rect 95670 31499 95734 31503
rect 95670 31479 95734 31483
rect 95670 31423 95674 31479
rect 95674 31423 95730 31479
rect 95730 31423 95734 31479
rect 95670 31419 95734 31423
rect 94081 31291 94145 31355
rect 92122 31181 92186 31185
rect 97189 31572 97253 31576
rect 97189 31516 97193 31572
rect 97193 31516 97249 31572
rect 97249 31516 97253 31572
rect 97189 31512 97253 31516
rect 97189 31492 97253 31496
rect 97189 31436 97193 31492
rect 97193 31436 97249 31492
rect 97249 31436 97253 31492
rect 97189 31432 97253 31436
rect 97934 30960 98318 31184
rect 99724 31237 99788 31241
rect 99724 31181 99728 31237
rect 99728 31181 99784 31237
rect 99784 31181 99788 31237
rect 99724 31177 99788 31181
rect 99804 31237 99868 31241
rect 99804 31181 99808 31237
rect 99808 31181 99864 31237
rect 99864 31181 99868 31237
rect 99804 31177 99868 31181
rect 99884 31237 99948 31241
rect 99884 31181 99888 31237
rect 99888 31181 99944 31237
rect 99944 31181 99948 31237
rect 99884 31177 99948 31181
rect 99964 31237 100028 31241
rect 99964 31181 99968 31237
rect 99968 31181 100024 31237
rect 100024 31181 100028 31237
rect 99964 31177 100028 31181
rect 100044 31237 100108 31241
rect 100044 31181 100048 31237
rect 100048 31181 100104 31237
rect 100104 31181 100108 31237
rect 100044 31177 100108 31181
rect 100124 31237 100188 31241
rect 100124 31181 100128 31237
rect 100128 31181 100184 31237
rect 100184 31181 100188 31237
rect 100124 31177 100188 31181
rect 100204 31237 100268 31241
rect 100204 31181 100208 31237
rect 100208 31181 100264 31237
rect 100264 31181 100268 31237
rect 100204 31177 100268 31181
rect 100284 31237 100348 31241
rect 100284 31181 100288 31237
rect 100288 31181 100344 31237
rect 100344 31181 100348 31237
rect 100284 31177 100348 31181
rect 100364 31237 100428 31241
rect 100364 31181 100368 31237
rect 100368 31181 100424 31237
rect 100424 31181 100428 31237
rect 100364 31177 100428 31181
rect 100444 31237 100508 31241
rect 100444 31181 100448 31237
rect 100448 31181 100504 31237
rect 100504 31181 100508 31237
rect 100444 31177 100508 31181
rect 100524 31237 100588 31241
rect 100524 31181 100528 31237
rect 100528 31181 100584 31237
rect 100584 31181 100588 31237
rect 100524 31177 100588 31181
rect 100604 31237 100668 31241
rect 100604 31181 100608 31237
rect 100608 31181 100664 31237
rect 100664 31181 100668 31237
rect 100604 31177 100668 31181
rect 100684 31237 100748 31241
rect 100684 31181 100688 31237
rect 100688 31181 100744 31237
rect 100744 31181 100748 31237
rect 100684 31177 100748 31181
rect 100764 31237 100828 31241
rect 100764 31181 100768 31237
rect 100768 31181 100824 31237
rect 100824 31181 100828 31237
rect 100764 31177 100828 31181
rect 100844 31237 100908 31241
rect 100844 31181 100848 31237
rect 100848 31181 100904 31237
rect 100904 31181 100908 31237
rect 100844 31177 100908 31181
rect 100924 31237 100988 31241
rect 100924 31181 100928 31237
rect 100928 31181 100984 31237
rect 100984 31181 100988 31237
rect 100924 31177 100988 31181
rect 101004 31237 101068 31241
rect 101004 31181 101008 31237
rect 101008 31181 101064 31237
rect 101064 31181 101068 31237
rect 101004 31177 101068 31181
rect 101084 31237 101148 31241
rect 101084 31181 101088 31237
rect 101088 31181 101144 31237
rect 101144 31181 101148 31237
rect 101084 31177 101148 31181
rect 101164 31237 101228 31241
rect 101164 31181 101168 31237
rect 101168 31181 101224 31237
rect 101224 31181 101228 31237
rect 101164 31177 101228 31181
rect 101244 31237 101308 31241
rect 101244 31181 101248 31237
rect 101248 31181 101304 31237
rect 101304 31181 101308 31237
rect 101244 31177 101308 31181
rect 101324 31237 101388 31241
rect 101324 31181 101328 31237
rect 101328 31181 101384 31237
rect 101384 31181 101388 31237
rect 101324 31177 101388 31181
rect 101404 31237 101468 31241
rect 101404 31181 101408 31237
rect 101408 31181 101464 31237
rect 101464 31181 101468 31237
rect 101404 31177 101468 31181
rect 101484 31237 101548 31241
rect 101484 31181 101488 31237
rect 101488 31181 101544 31237
rect 101544 31181 101548 31237
rect 101484 31177 101548 31181
rect 101564 31237 101628 31241
rect 101564 31181 101568 31237
rect 101568 31181 101624 31237
rect 101624 31181 101628 31237
rect 101564 31177 101628 31181
rect 101644 31237 101708 31241
rect 101644 31181 101648 31237
rect 101648 31181 101704 31237
rect 101704 31181 101708 31237
rect 101644 31177 101708 31181
rect 101724 31237 101788 31241
rect 101724 31181 101728 31237
rect 101728 31181 101784 31237
rect 101784 31181 101788 31237
rect 101724 31177 101788 31181
rect 101804 31237 101868 31241
rect 101804 31181 101808 31237
rect 101808 31181 101864 31237
rect 101864 31181 101868 31237
rect 101804 31177 101868 31181
rect 101884 31237 101948 31241
rect 101884 31181 101888 31237
rect 101888 31181 101944 31237
rect 101944 31181 101948 31237
rect 101884 31177 101948 31181
rect 101964 31237 102028 31241
rect 101964 31181 101968 31237
rect 101968 31181 102024 31237
rect 102024 31181 102028 31237
rect 101964 31177 102028 31181
rect 102044 31237 102108 31241
rect 102044 31181 102048 31237
rect 102048 31181 102104 31237
rect 102104 31181 102108 31237
rect 102044 31177 102108 31181
rect 102124 31237 102188 31241
rect 102124 31181 102128 31237
rect 102128 31181 102184 31237
rect 102184 31181 102188 31237
rect 102124 31177 102188 31181
rect 102204 31237 102268 31241
rect 102204 31181 102208 31237
rect 102208 31181 102264 31237
rect 102264 31181 102268 31237
rect 102204 31177 102268 31181
rect 102284 31237 102348 31241
rect 102284 31181 102288 31237
rect 102288 31181 102344 31237
rect 102344 31181 102348 31237
rect 102284 31177 102348 31181
rect 102364 31237 102428 31241
rect 102364 31181 102368 31237
rect 102368 31181 102424 31237
rect 102424 31181 102428 31237
rect 102364 31177 102428 31181
rect 102444 31237 102508 31241
rect 102444 31181 102448 31237
rect 102448 31181 102504 31237
rect 102504 31181 102508 31237
rect 102444 31177 102508 31181
rect 102524 31237 102588 31241
rect 102524 31181 102528 31237
rect 102528 31181 102584 31237
rect 102584 31181 102588 31237
rect 102524 31177 102588 31181
rect 102604 31237 102668 31241
rect 102604 31181 102608 31237
rect 102608 31181 102664 31237
rect 102664 31181 102668 31237
rect 102604 31177 102668 31181
rect 102684 31237 102748 31241
rect 102684 31181 102688 31237
rect 102688 31181 102744 31237
rect 102744 31181 102748 31237
rect 102684 31177 102748 31181
rect 102764 31237 102828 31241
rect 102764 31181 102768 31237
rect 102768 31181 102824 31237
rect 102824 31181 102828 31237
rect 102764 31177 102828 31181
rect 102844 31237 102908 31241
rect 102844 31181 102848 31237
rect 102848 31181 102904 31237
rect 102904 31181 102908 31237
rect 102844 31177 102908 31181
rect 102924 31237 102988 31241
rect 102924 31181 102928 31237
rect 102928 31181 102984 31237
rect 102984 31181 102988 31237
rect 102924 31177 102988 31181
rect 92121 29903 92185 29907
rect 92121 29847 92125 29903
rect 92125 29847 92181 29903
rect 92181 29847 92185 29903
rect 92121 29843 92185 29847
rect 94081 30267 94145 30271
rect 94081 30211 94085 30267
rect 94085 30211 94141 30267
rect 94141 30211 94145 30267
rect 94081 30207 94145 30211
rect 95665 30228 95729 30232
rect 95665 30172 95669 30228
rect 95669 30172 95725 30228
rect 95725 30172 95729 30228
rect 95665 30168 95729 30172
rect 95665 30148 95729 30152
rect 95665 30092 95669 30148
rect 95669 30092 95725 30148
rect 95725 30092 95729 30148
rect 95665 30088 95729 30092
rect 97194 30225 97258 30229
rect 97194 30169 97198 30225
rect 97198 30169 97254 30225
rect 97254 30169 97258 30225
rect 97194 30165 97258 30169
rect 97194 30145 97258 30149
rect 97194 30089 97198 30145
rect 97198 30089 97254 30145
rect 97254 30089 97258 30145
rect 97194 30085 97258 30089
rect 94081 29119 94145 29183
rect 95664 28875 95728 28879
rect 95664 28819 95668 28875
rect 95668 28819 95724 28875
rect 95724 28819 95728 28875
rect 95664 28815 95728 28819
rect 95664 28795 95728 28799
rect 95664 28739 95668 28795
rect 95668 28739 95724 28795
rect 95724 28739 95728 28795
rect 95664 28735 95728 28739
rect 92129 28510 92193 28514
rect 92129 28454 92133 28510
rect 92133 28454 92189 28510
rect 92189 28454 92193 28510
rect 92129 28450 92193 28454
rect 94082 28091 94146 28095
rect 94082 28035 94086 28091
rect 94086 28035 94142 28091
rect 94142 28035 94146 28091
rect 94082 28031 94146 28035
rect 97194 28853 97258 28857
rect 97194 28797 97198 28853
rect 97198 28797 97254 28853
rect 97254 28797 97258 28853
rect 97194 28793 97258 28797
rect 97194 28773 97258 28777
rect 97194 28717 97198 28773
rect 97198 28717 97254 28773
rect 97254 28717 97258 28773
rect 97194 28713 97258 28717
rect 97932 28057 98316 28281
rect 99701 28238 99765 28242
rect 99701 28182 99705 28238
rect 99705 28182 99761 28238
rect 99761 28182 99765 28238
rect 99701 28178 99765 28182
rect 99781 28238 99845 28242
rect 99781 28182 99785 28238
rect 99785 28182 99841 28238
rect 99841 28182 99845 28238
rect 99781 28178 99845 28182
rect 99861 28238 99925 28242
rect 99861 28182 99865 28238
rect 99865 28182 99921 28238
rect 99921 28182 99925 28238
rect 99861 28178 99925 28182
rect 99941 28238 100005 28242
rect 99941 28182 99945 28238
rect 99945 28182 100001 28238
rect 100001 28182 100005 28238
rect 99941 28178 100005 28182
rect 100021 28238 100085 28242
rect 100021 28182 100025 28238
rect 100025 28182 100081 28238
rect 100081 28182 100085 28238
rect 100021 28178 100085 28182
rect 100101 28238 100165 28242
rect 100101 28182 100105 28238
rect 100105 28182 100161 28238
rect 100161 28182 100165 28238
rect 100101 28178 100165 28182
rect 100181 28238 100245 28242
rect 100181 28182 100185 28238
rect 100185 28182 100241 28238
rect 100241 28182 100245 28238
rect 100181 28178 100245 28182
rect 100261 28238 100325 28242
rect 100261 28182 100265 28238
rect 100265 28182 100321 28238
rect 100321 28182 100325 28238
rect 100261 28178 100325 28182
rect 100341 28238 100405 28242
rect 100341 28182 100345 28238
rect 100345 28182 100401 28238
rect 100401 28182 100405 28238
rect 100341 28178 100405 28182
rect 100421 28238 100485 28242
rect 100421 28182 100425 28238
rect 100425 28182 100481 28238
rect 100481 28182 100485 28238
rect 100421 28178 100485 28182
rect 100501 28238 100565 28242
rect 100501 28182 100505 28238
rect 100505 28182 100561 28238
rect 100561 28182 100565 28238
rect 100501 28178 100565 28182
rect 100581 28238 100645 28242
rect 100581 28182 100585 28238
rect 100585 28182 100641 28238
rect 100641 28182 100645 28238
rect 100581 28178 100645 28182
rect 100661 28238 100725 28242
rect 100661 28182 100665 28238
rect 100665 28182 100721 28238
rect 100721 28182 100725 28238
rect 100661 28178 100725 28182
rect 100741 28238 100805 28242
rect 100741 28182 100745 28238
rect 100745 28182 100801 28238
rect 100801 28182 100805 28238
rect 100741 28178 100805 28182
rect 100821 28238 100885 28242
rect 100821 28182 100825 28238
rect 100825 28182 100881 28238
rect 100881 28182 100885 28238
rect 100821 28178 100885 28182
rect 100901 28238 100965 28242
rect 100901 28182 100905 28238
rect 100905 28182 100961 28238
rect 100961 28182 100965 28238
rect 100901 28178 100965 28182
rect 100981 28238 101045 28242
rect 100981 28182 100985 28238
rect 100985 28182 101041 28238
rect 101041 28182 101045 28238
rect 100981 28178 101045 28182
rect 101061 28238 101125 28242
rect 101061 28182 101065 28238
rect 101065 28182 101121 28238
rect 101121 28182 101125 28238
rect 101061 28178 101125 28182
rect 101141 28238 101205 28242
rect 101141 28182 101145 28238
rect 101145 28182 101201 28238
rect 101201 28182 101205 28238
rect 101141 28178 101205 28182
rect 101221 28238 101285 28242
rect 101221 28182 101225 28238
rect 101225 28182 101281 28238
rect 101281 28182 101285 28238
rect 101221 28178 101285 28182
rect 101301 28238 101365 28242
rect 101301 28182 101305 28238
rect 101305 28182 101361 28238
rect 101361 28182 101365 28238
rect 101301 28178 101365 28182
rect 101381 28238 101445 28242
rect 101381 28182 101385 28238
rect 101385 28182 101441 28238
rect 101441 28182 101445 28238
rect 101381 28178 101445 28182
rect 101461 28238 101525 28242
rect 101461 28182 101465 28238
rect 101465 28182 101521 28238
rect 101521 28182 101525 28238
rect 101461 28178 101525 28182
rect 101541 28238 101605 28242
rect 101541 28182 101545 28238
rect 101545 28182 101601 28238
rect 101601 28182 101605 28238
rect 101541 28178 101605 28182
rect 101621 28238 101685 28242
rect 101621 28182 101625 28238
rect 101625 28182 101681 28238
rect 101681 28182 101685 28238
rect 101621 28178 101685 28182
rect 101701 28238 101765 28242
rect 101701 28182 101705 28238
rect 101705 28182 101761 28238
rect 101761 28182 101765 28238
rect 101701 28178 101765 28182
rect 101781 28238 101845 28242
rect 101781 28182 101785 28238
rect 101785 28182 101841 28238
rect 101841 28182 101845 28238
rect 101781 28178 101845 28182
rect 101861 28238 101925 28242
rect 101861 28182 101865 28238
rect 101865 28182 101921 28238
rect 101921 28182 101925 28238
rect 101861 28178 101925 28182
rect 101941 28238 102005 28242
rect 101941 28182 101945 28238
rect 101945 28182 102001 28238
rect 102001 28182 102005 28238
rect 101941 28178 102005 28182
rect 102021 28238 102085 28242
rect 102021 28182 102025 28238
rect 102025 28182 102081 28238
rect 102081 28182 102085 28238
rect 102021 28178 102085 28182
rect 102101 28238 102165 28242
rect 102101 28182 102105 28238
rect 102105 28182 102161 28238
rect 102161 28182 102165 28238
rect 102101 28178 102165 28182
rect 102181 28238 102245 28242
rect 102181 28182 102185 28238
rect 102185 28182 102241 28238
rect 102241 28182 102245 28238
rect 102181 28178 102245 28182
rect 102261 28238 102325 28242
rect 102261 28182 102265 28238
rect 102265 28182 102321 28238
rect 102321 28182 102325 28238
rect 102261 28178 102325 28182
rect 102341 28238 102405 28242
rect 102341 28182 102345 28238
rect 102345 28182 102401 28238
rect 102401 28182 102405 28238
rect 102341 28178 102405 28182
rect 102421 28238 102485 28242
rect 102421 28182 102425 28238
rect 102425 28182 102481 28238
rect 102481 28182 102485 28238
rect 102421 28178 102485 28182
rect 102501 28238 102565 28242
rect 102501 28182 102505 28238
rect 102505 28182 102561 28238
rect 102561 28182 102565 28238
rect 102501 28178 102565 28182
rect 102581 28238 102645 28242
rect 102581 28182 102585 28238
rect 102585 28182 102641 28238
rect 102641 28182 102645 28238
rect 102581 28178 102645 28182
rect 102661 28238 102725 28242
rect 102661 28182 102665 28238
rect 102665 28182 102721 28238
rect 102721 28182 102725 28238
rect 102661 28178 102725 28182
rect 102741 28238 102805 28242
rect 102741 28182 102745 28238
rect 102745 28182 102801 28238
rect 102801 28182 102805 28238
rect 102741 28178 102805 28182
rect 102821 28238 102885 28242
rect 102821 28182 102825 28238
rect 102825 28182 102881 28238
rect 102881 28182 102885 28238
rect 102821 28178 102885 28182
rect 102901 28238 102965 28242
rect 102901 28182 102905 28238
rect 102905 28182 102961 28238
rect 102961 28182 102965 28238
rect 102901 28178 102965 28182
rect 102981 28238 103045 28242
rect 102981 28182 102985 28238
rect 102985 28182 103041 28238
rect 103041 28182 103045 28238
rect 102981 28178 103045 28182
rect 92125 27140 92189 27144
rect 92125 27084 92129 27140
rect 92129 27084 92185 27140
rect 92185 27084 92189 27140
rect 95667 27475 95731 27479
rect 95667 27419 95671 27475
rect 95671 27419 95727 27475
rect 95727 27419 95731 27475
rect 95667 27415 95731 27419
rect 95667 27395 95731 27399
rect 95667 27339 95671 27395
rect 95671 27339 95727 27395
rect 95727 27339 95731 27395
rect 95667 27335 95731 27339
rect 97191 27469 97255 27473
rect 97191 27413 97195 27469
rect 97195 27413 97251 27469
rect 97251 27413 97255 27469
rect 97191 27409 97255 27413
rect 97191 27389 97255 27393
rect 97191 27333 97195 27389
rect 97195 27333 97251 27389
rect 97251 27333 97255 27389
rect 97191 27329 97255 27333
rect 92125 27080 92189 27084
rect 93160 26232 93224 26236
rect 93160 26176 93164 26232
rect 93164 26176 93220 26232
rect 93220 26176 93224 26232
rect 93160 26172 93224 26176
rect 94001 25644 94225 25868
rect 92583 25609 92647 25613
rect 92583 25553 92587 25609
rect 92587 25553 92643 25609
rect 92643 25553 92647 25609
rect 92583 25549 92647 25553
rect 93725 25547 93789 25551
rect 93725 25491 93729 25547
rect 93729 25491 93785 25547
rect 93785 25491 93789 25547
rect 93725 25487 93789 25491
rect 57416 24239 78200 24243
rect 57416 24103 57420 24239
rect 57420 24103 78196 24239
rect 78196 24103 78200 24239
rect 57416 24099 78200 24103
rect 92122 24301 92186 24305
rect 92122 24245 92126 24301
rect 92126 24245 92182 24301
rect 92182 24245 92186 24301
rect 95670 24619 95734 24623
rect 95670 24563 95674 24619
rect 95674 24563 95730 24619
rect 95730 24563 95734 24619
rect 95670 24559 95734 24563
rect 95670 24539 95734 24543
rect 95670 24483 95674 24539
rect 95674 24483 95730 24539
rect 95730 24483 95734 24539
rect 95670 24479 95734 24483
rect 94081 24351 94145 24415
rect 92122 24241 92186 24245
rect 97189 24632 97253 24636
rect 97189 24576 97193 24632
rect 97193 24576 97249 24632
rect 97249 24576 97253 24632
rect 97189 24572 97253 24576
rect 97189 24552 97253 24556
rect 97189 24496 97193 24552
rect 97193 24496 97249 24552
rect 97249 24496 97253 24552
rect 97189 24492 97253 24496
rect 97934 24020 98318 24244
rect 99726 24304 99790 24308
rect 99726 24248 99730 24304
rect 99730 24248 99786 24304
rect 99786 24248 99790 24304
rect 99726 24244 99790 24248
rect 99806 24304 99870 24308
rect 99806 24248 99810 24304
rect 99810 24248 99866 24304
rect 99866 24248 99870 24304
rect 99806 24244 99870 24248
rect 99886 24304 99950 24308
rect 99886 24248 99890 24304
rect 99890 24248 99946 24304
rect 99946 24248 99950 24304
rect 99886 24244 99950 24248
rect 99966 24304 100030 24308
rect 99966 24248 99970 24304
rect 99970 24248 100026 24304
rect 100026 24248 100030 24304
rect 99966 24244 100030 24248
rect 100046 24304 100110 24308
rect 100046 24248 100050 24304
rect 100050 24248 100106 24304
rect 100106 24248 100110 24304
rect 100046 24244 100110 24248
rect 100126 24304 100190 24308
rect 100126 24248 100130 24304
rect 100130 24248 100186 24304
rect 100186 24248 100190 24304
rect 100126 24244 100190 24248
rect 100206 24304 100270 24308
rect 100206 24248 100210 24304
rect 100210 24248 100266 24304
rect 100266 24248 100270 24304
rect 100206 24244 100270 24248
rect 100286 24304 100350 24308
rect 100286 24248 100290 24304
rect 100290 24248 100346 24304
rect 100346 24248 100350 24304
rect 100286 24244 100350 24248
rect 100366 24304 100430 24308
rect 100366 24248 100370 24304
rect 100370 24248 100426 24304
rect 100426 24248 100430 24304
rect 100366 24244 100430 24248
rect 100446 24304 100510 24308
rect 100446 24248 100450 24304
rect 100450 24248 100506 24304
rect 100506 24248 100510 24304
rect 100446 24244 100510 24248
rect 100526 24304 100590 24308
rect 100526 24248 100530 24304
rect 100530 24248 100586 24304
rect 100586 24248 100590 24304
rect 100526 24244 100590 24248
rect 100606 24304 100670 24308
rect 100606 24248 100610 24304
rect 100610 24248 100666 24304
rect 100666 24248 100670 24304
rect 100606 24244 100670 24248
rect 100686 24304 100750 24308
rect 100686 24248 100690 24304
rect 100690 24248 100746 24304
rect 100746 24248 100750 24304
rect 100686 24244 100750 24248
rect 100766 24304 100830 24308
rect 100766 24248 100770 24304
rect 100770 24248 100826 24304
rect 100826 24248 100830 24304
rect 100766 24244 100830 24248
rect 100846 24304 100910 24308
rect 100846 24248 100850 24304
rect 100850 24248 100906 24304
rect 100906 24248 100910 24304
rect 100846 24244 100910 24248
rect 100926 24304 100990 24308
rect 100926 24248 100930 24304
rect 100930 24248 100986 24304
rect 100986 24248 100990 24304
rect 100926 24244 100990 24248
rect 101006 24304 101070 24308
rect 101006 24248 101010 24304
rect 101010 24248 101066 24304
rect 101066 24248 101070 24304
rect 101006 24244 101070 24248
rect 101086 24304 101150 24308
rect 101086 24248 101090 24304
rect 101090 24248 101146 24304
rect 101146 24248 101150 24304
rect 101086 24244 101150 24248
rect 101166 24304 101230 24308
rect 101166 24248 101170 24304
rect 101170 24248 101226 24304
rect 101226 24248 101230 24304
rect 101166 24244 101230 24248
rect 101246 24304 101310 24308
rect 101246 24248 101250 24304
rect 101250 24248 101306 24304
rect 101306 24248 101310 24304
rect 101246 24244 101310 24248
rect 101326 24304 101390 24308
rect 101326 24248 101330 24304
rect 101330 24248 101386 24304
rect 101386 24248 101390 24304
rect 101326 24244 101390 24248
rect 101406 24304 101470 24308
rect 101406 24248 101410 24304
rect 101410 24248 101466 24304
rect 101466 24248 101470 24304
rect 101406 24244 101470 24248
rect 101486 24304 101550 24308
rect 101486 24248 101490 24304
rect 101490 24248 101546 24304
rect 101546 24248 101550 24304
rect 101486 24244 101550 24248
rect 101566 24304 101630 24308
rect 101566 24248 101570 24304
rect 101570 24248 101626 24304
rect 101626 24248 101630 24304
rect 101566 24244 101630 24248
rect 101646 24304 101710 24308
rect 101646 24248 101650 24304
rect 101650 24248 101706 24304
rect 101706 24248 101710 24304
rect 101646 24244 101710 24248
rect 101726 24304 101790 24308
rect 101726 24248 101730 24304
rect 101730 24248 101786 24304
rect 101786 24248 101790 24304
rect 101726 24244 101790 24248
rect 101806 24304 101870 24308
rect 101806 24248 101810 24304
rect 101810 24248 101866 24304
rect 101866 24248 101870 24304
rect 101806 24244 101870 24248
rect 101886 24304 101950 24308
rect 101886 24248 101890 24304
rect 101890 24248 101946 24304
rect 101946 24248 101950 24304
rect 101886 24244 101950 24248
rect 101966 24304 102030 24308
rect 101966 24248 101970 24304
rect 101970 24248 102026 24304
rect 102026 24248 102030 24304
rect 101966 24244 102030 24248
rect 102046 24304 102110 24308
rect 102046 24248 102050 24304
rect 102050 24248 102106 24304
rect 102106 24248 102110 24304
rect 102046 24244 102110 24248
rect 102126 24304 102190 24308
rect 102126 24248 102130 24304
rect 102130 24248 102186 24304
rect 102186 24248 102190 24304
rect 102126 24244 102190 24248
rect 102206 24304 102270 24308
rect 102206 24248 102210 24304
rect 102210 24248 102266 24304
rect 102266 24248 102270 24304
rect 102206 24244 102270 24248
rect 102286 24304 102350 24308
rect 102286 24248 102290 24304
rect 102290 24248 102346 24304
rect 102346 24248 102350 24304
rect 102286 24244 102350 24248
rect 102366 24304 102430 24308
rect 102366 24248 102370 24304
rect 102370 24248 102426 24304
rect 102426 24248 102430 24304
rect 102366 24244 102430 24248
rect 102446 24304 102510 24308
rect 102446 24248 102450 24304
rect 102450 24248 102506 24304
rect 102506 24248 102510 24304
rect 102446 24244 102510 24248
rect 102526 24304 102590 24308
rect 102526 24248 102530 24304
rect 102530 24248 102586 24304
rect 102586 24248 102590 24304
rect 102526 24244 102590 24248
rect 102606 24304 102670 24308
rect 102606 24248 102610 24304
rect 102610 24248 102666 24304
rect 102666 24248 102670 24304
rect 102606 24244 102670 24248
rect 102686 24304 102750 24308
rect 102686 24248 102690 24304
rect 102690 24248 102746 24304
rect 102746 24248 102750 24304
rect 102686 24244 102750 24248
rect 102766 24304 102830 24308
rect 102766 24248 102770 24304
rect 102770 24248 102826 24304
rect 102826 24248 102830 24304
rect 102766 24244 102830 24248
rect 102846 24304 102910 24308
rect 102846 24248 102850 24304
rect 102850 24248 102906 24304
rect 102906 24248 102910 24304
rect 102846 24244 102910 24248
rect 102926 24304 102990 24308
rect 102926 24248 102930 24304
rect 102930 24248 102986 24304
rect 102986 24248 102990 24304
rect 102926 24244 102990 24248
rect 92121 22963 92185 22967
rect 92121 22907 92125 22963
rect 92125 22907 92181 22963
rect 92181 22907 92185 22963
rect 92121 22903 92185 22907
rect 94081 23327 94145 23331
rect 94081 23271 94085 23327
rect 94085 23271 94141 23327
rect 94141 23271 94145 23327
rect 94081 23267 94145 23271
rect 95665 23288 95729 23292
rect 95665 23232 95669 23288
rect 95669 23232 95725 23288
rect 95725 23232 95729 23288
rect 95665 23228 95729 23232
rect 95665 23208 95729 23212
rect 95665 23152 95669 23208
rect 95669 23152 95725 23208
rect 95725 23152 95729 23208
rect 95665 23148 95729 23152
rect 97194 23285 97258 23289
rect 97194 23229 97198 23285
rect 97198 23229 97254 23285
rect 97254 23229 97258 23285
rect 97194 23225 97258 23229
rect 97194 23205 97258 23209
rect 97194 23149 97198 23205
rect 97198 23149 97254 23205
rect 97254 23149 97258 23205
rect 97194 23145 97258 23149
rect 94081 22179 94145 22243
rect 95664 21935 95728 21939
rect 95664 21879 95668 21935
rect 95668 21879 95724 21935
rect 95724 21879 95728 21935
rect 95664 21875 95728 21879
rect 95664 21855 95728 21859
rect 95664 21799 95668 21855
rect 95668 21799 95724 21855
rect 95724 21799 95728 21855
rect 95664 21795 95728 21799
rect 92129 21570 92193 21574
rect 92129 21514 92133 21570
rect 92133 21514 92189 21570
rect 92189 21514 92193 21570
rect 92129 21510 92193 21514
rect 94082 21151 94146 21155
rect 94082 21095 94086 21151
rect 94086 21095 94142 21151
rect 94142 21095 94146 21151
rect 94082 21091 94146 21095
rect 97194 21913 97258 21917
rect 97194 21857 97198 21913
rect 97198 21857 97254 21913
rect 97254 21857 97258 21913
rect 97194 21853 97258 21857
rect 97194 21833 97258 21837
rect 97194 21777 97198 21833
rect 97198 21777 97254 21833
rect 97254 21777 97258 21833
rect 97194 21773 97258 21777
rect 97932 21117 98316 21341
rect 99682 21298 99746 21302
rect 99682 21242 99686 21298
rect 99686 21242 99742 21298
rect 99742 21242 99746 21298
rect 99682 21238 99746 21242
rect 99762 21298 99826 21302
rect 99762 21242 99766 21298
rect 99766 21242 99822 21298
rect 99822 21242 99826 21298
rect 99762 21238 99826 21242
rect 99842 21298 99906 21302
rect 99842 21242 99846 21298
rect 99846 21242 99902 21298
rect 99902 21242 99906 21298
rect 99842 21238 99906 21242
rect 99922 21298 99986 21302
rect 99922 21242 99926 21298
rect 99926 21242 99982 21298
rect 99982 21242 99986 21298
rect 99922 21238 99986 21242
rect 100002 21298 100066 21302
rect 100002 21242 100006 21298
rect 100006 21242 100062 21298
rect 100062 21242 100066 21298
rect 100002 21238 100066 21242
rect 100082 21298 100146 21302
rect 100082 21242 100086 21298
rect 100086 21242 100142 21298
rect 100142 21242 100146 21298
rect 100082 21238 100146 21242
rect 100162 21298 100226 21302
rect 100162 21242 100166 21298
rect 100166 21242 100222 21298
rect 100222 21242 100226 21298
rect 100162 21238 100226 21242
rect 100242 21298 100306 21302
rect 100242 21242 100246 21298
rect 100246 21242 100302 21298
rect 100302 21242 100306 21298
rect 100242 21238 100306 21242
rect 100322 21298 100386 21302
rect 100322 21242 100326 21298
rect 100326 21242 100382 21298
rect 100382 21242 100386 21298
rect 100322 21238 100386 21242
rect 100402 21298 100466 21302
rect 100402 21242 100406 21298
rect 100406 21242 100462 21298
rect 100462 21242 100466 21298
rect 100402 21238 100466 21242
rect 100482 21298 100546 21302
rect 100482 21242 100486 21298
rect 100486 21242 100542 21298
rect 100542 21242 100546 21298
rect 100482 21238 100546 21242
rect 100562 21298 100626 21302
rect 100562 21242 100566 21298
rect 100566 21242 100622 21298
rect 100622 21242 100626 21298
rect 100562 21238 100626 21242
rect 100642 21298 100706 21302
rect 100642 21242 100646 21298
rect 100646 21242 100702 21298
rect 100702 21242 100706 21298
rect 100642 21238 100706 21242
rect 100722 21298 100786 21302
rect 100722 21242 100726 21298
rect 100726 21242 100782 21298
rect 100782 21242 100786 21298
rect 100722 21238 100786 21242
rect 100802 21298 100866 21302
rect 100802 21242 100806 21298
rect 100806 21242 100862 21298
rect 100862 21242 100866 21298
rect 100802 21238 100866 21242
rect 100882 21298 100946 21302
rect 100882 21242 100886 21298
rect 100886 21242 100942 21298
rect 100942 21242 100946 21298
rect 100882 21238 100946 21242
rect 100962 21298 101026 21302
rect 100962 21242 100966 21298
rect 100966 21242 101022 21298
rect 101022 21242 101026 21298
rect 100962 21238 101026 21242
rect 101042 21298 101106 21302
rect 101042 21242 101046 21298
rect 101046 21242 101102 21298
rect 101102 21242 101106 21298
rect 101042 21238 101106 21242
rect 101122 21298 101186 21302
rect 101122 21242 101126 21298
rect 101126 21242 101182 21298
rect 101182 21242 101186 21298
rect 101122 21238 101186 21242
rect 101202 21298 101266 21302
rect 101202 21242 101206 21298
rect 101206 21242 101262 21298
rect 101262 21242 101266 21298
rect 101202 21238 101266 21242
rect 101282 21298 101346 21302
rect 101282 21242 101286 21298
rect 101286 21242 101342 21298
rect 101342 21242 101346 21298
rect 101282 21238 101346 21242
rect 101362 21298 101426 21302
rect 101362 21242 101366 21298
rect 101366 21242 101422 21298
rect 101422 21242 101426 21298
rect 101362 21238 101426 21242
rect 101442 21298 101506 21302
rect 101442 21242 101446 21298
rect 101446 21242 101502 21298
rect 101502 21242 101506 21298
rect 101442 21238 101506 21242
rect 101522 21298 101586 21302
rect 101522 21242 101526 21298
rect 101526 21242 101582 21298
rect 101582 21242 101586 21298
rect 101522 21238 101586 21242
rect 101602 21298 101666 21302
rect 101602 21242 101606 21298
rect 101606 21242 101662 21298
rect 101662 21242 101666 21298
rect 101602 21238 101666 21242
rect 101682 21298 101746 21302
rect 101682 21242 101686 21298
rect 101686 21242 101742 21298
rect 101742 21242 101746 21298
rect 101682 21238 101746 21242
rect 101762 21298 101826 21302
rect 101762 21242 101766 21298
rect 101766 21242 101822 21298
rect 101822 21242 101826 21298
rect 101762 21238 101826 21242
rect 101842 21298 101906 21302
rect 101842 21242 101846 21298
rect 101846 21242 101902 21298
rect 101902 21242 101906 21298
rect 101842 21238 101906 21242
rect 101922 21298 101986 21302
rect 101922 21242 101926 21298
rect 101926 21242 101982 21298
rect 101982 21242 101986 21298
rect 101922 21238 101986 21242
rect 102002 21298 102066 21302
rect 102002 21242 102006 21298
rect 102006 21242 102062 21298
rect 102062 21242 102066 21298
rect 102002 21238 102066 21242
rect 102082 21298 102146 21302
rect 102082 21242 102086 21298
rect 102086 21242 102142 21298
rect 102142 21242 102146 21298
rect 102082 21238 102146 21242
rect 102162 21298 102226 21302
rect 102162 21242 102166 21298
rect 102166 21242 102222 21298
rect 102222 21242 102226 21298
rect 102162 21238 102226 21242
rect 102242 21298 102306 21302
rect 102242 21242 102246 21298
rect 102246 21242 102302 21298
rect 102302 21242 102306 21298
rect 102242 21238 102306 21242
rect 102322 21298 102386 21302
rect 102322 21242 102326 21298
rect 102326 21242 102382 21298
rect 102382 21242 102386 21298
rect 102322 21238 102386 21242
rect 102402 21298 102466 21302
rect 102402 21242 102406 21298
rect 102406 21242 102462 21298
rect 102462 21242 102466 21298
rect 102402 21238 102466 21242
rect 102482 21298 102546 21302
rect 102482 21242 102486 21298
rect 102486 21242 102542 21298
rect 102542 21242 102546 21298
rect 102482 21238 102546 21242
rect 102562 21298 102626 21302
rect 102562 21242 102566 21298
rect 102566 21242 102622 21298
rect 102622 21242 102626 21298
rect 102562 21238 102626 21242
rect 102642 21298 102706 21302
rect 102642 21242 102646 21298
rect 102646 21242 102702 21298
rect 102702 21242 102706 21298
rect 102642 21238 102706 21242
rect 102722 21298 102786 21302
rect 102722 21242 102726 21298
rect 102726 21242 102782 21298
rect 102782 21242 102786 21298
rect 102722 21238 102786 21242
rect 102802 21298 102866 21302
rect 102802 21242 102806 21298
rect 102806 21242 102862 21298
rect 102862 21242 102866 21298
rect 102802 21238 102866 21242
rect 102882 21298 102946 21302
rect 102882 21242 102886 21298
rect 102886 21242 102942 21298
rect 102942 21242 102946 21298
rect 102882 21238 102946 21242
rect 102962 21298 103026 21302
rect 102962 21242 102966 21298
rect 102966 21242 103022 21298
rect 103022 21242 103026 21298
rect 102962 21238 103026 21242
rect 78296 20449 78360 20513
rect 92125 20200 92189 20204
rect 92125 20144 92129 20200
rect 92129 20144 92185 20200
rect 92185 20144 92189 20200
rect 95667 20535 95731 20539
rect 95667 20479 95671 20535
rect 95671 20479 95727 20535
rect 95727 20479 95731 20535
rect 95667 20475 95731 20479
rect 95667 20455 95731 20459
rect 95667 20399 95671 20455
rect 95671 20399 95727 20455
rect 95727 20399 95731 20455
rect 95667 20395 95731 20399
rect 97191 20529 97255 20533
rect 97191 20473 97195 20529
rect 97195 20473 97251 20529
rect 97251 20473 97255 20529
rect 97191 20469 97255 20473
rect 97191 20449 97255 20453
rect 97191 20393 97195 20449
rect 97195 20393 97251 20449
rect 97251 20393 97255 20449
rect 97191 20389 97255 20393
rect 92125 20140 92189 20144
rect 78296 19977 78360 20041
rect 78296 19442 78360 19506
rect 78296 18979 78360 19043
rect 53513 17174 53577 17178
rect 53513 17118 53517 17174
rect 53517 17118 53573 17174
rect 53573 17118 53577 17174
rect 53513 17114 53577 17118
rect 53513 17094 53577 17098
rect 53513 17038 53517 17094
rect 53517 17038 53573 17094
rect 53573 17038 53577 17094
rect 53513 17034 53577 17038
rect 53513 17014 53577 17018
rect 53513 16958 53517 17014
rect 53517 16958 53573 17014
rect 53573 16958 53577 17014
rect 53513 16954 53577 16958
rect 53513 16934 53577 16938
rect 53513 16878 53517 16934
rect 53517 16878 53573 16934
rect 53573 16878 53577 16934
rect 53513 16874 53577 16878
rect 53513 16854 53577 16858
rect 53513 16798 53517 16854
rect 53517 16798 53573 16854
rect 53573 16798 53577 16854
rect 53513 16794 53577 16798
rect 53513 16774 53577 16778
rect 53513 16718 53517 16774
rect 53517 16718 53573 16774
rect 53573 16718 53577 16774
rect 53513 16714 53577 16718
rect 53513 16694 53577 16698
rect 53513 16638 53517 16694
rect 53517 16638 53573 16694
rect 53573 16638 53577 16694
rect 53513 16634 53577 16638
rect 53513 16614 53577 16618
rect 53513 16558 53517 16614
rect 53517 16558 53573 16614
rect 53573 16558 53577 16614
rect 53513 16554 53577 16558
rect 53513 16534 53577 16538
rect 53513 16478 53517 16534
rect 53517 16478 53573 16534
rect 53573 16478 53577 16534
rect 53513 16474 53577 16478
rect 53513 16454 53577 16458
rect 53513 16398 53517 16454
rect 53517 16398 53573 16454
rect 53573 16398 53577 16454
rect 53513 16394 53577 16398
rect 53513 16374 53577 16378
rect 53513 16318 53517 16374
rect 53517 16318 53573 16374
rect 53573 16318 53577 16374
rect 53513 16314 53577 16318
rect 53513 16294 53577 16298
rect 53513 16238 53517 16294
rect 53517 16238 53573 16294
rect 53573 16238 53577 16294
rect 53513 16234 53577 16238
rect 53513 16214 53577 16218
rect 53513 16158 53517 16214
rect 53517 16158 53573 16214
rect 53573 16158 53577 16214
rect 53513 16154 53577 16158
rect 53513 16134 53577 16138
rect 53513 16078 53517 16134
rect 53517 16078 53573 16134
rect 53573 16078 53577 16134
rect 53513 16074 53577 16078
rect 53513 16054 53577 16058
rect 53513 15998 53517 16054
rect 53517 15998 53573 16054
rect 53573 15998 53577 16054
rect 53513 15994 53577 15998
rect 53513 15974 53577 15978
rect 53513 15918 53517 15974
rect 53517 15918 53573 15974
rect 53573 15918 53577 15974
rect 53513 15914 53577 15918
rect 53513 15894 53577 15898
rect 53513 15838 53517 15894
rect 53517 15838 53573 15894
rect 53573 15838 53577 15894
rect 53513 15834 53577 15838
rect 53513 15814 53577 15818
rect 53513 15758 53517 15814
rect 53517 15758 53573 15814
rect 53573 15758 53577 15814
rect 53513 15754 53577 15758
rect 53513 15734 53577 15738
rect 53513 15678 53517 15734
rect 53517 15678 53573 15734
rect 53573 15678 53577 15734
rect 53513 15674 53577 15678
rect 53513 15654 53577 15658
rect 53513 15598 53517 15654
rect 53517 15598 53573 15654
rect 53573 15598 53577 15654
rect 53513 15594 53577 15598
rect 53513 15574 53577 15578
rect 53513 15518 53517 15574
rect 53517 15518 53573 15574
rect 53573 15518 53577 15574
rect 53513 15514 53577 15518
rect 53513 15494 53577 15498
rect 53513 15438 53517 15494
rect 53517 15438 53573 15494
rect 53573 15438 53577 15494
rect 53513 15434 53577 15438
rect 53513 15414 53577 15418
rect 53513 15358 53517 15414
rect 53517 15358 53573 15414
rect 53573 15358 53577 15414
rect 53513 15354 53577 15358
rect 53513 15334 53577 15338
rect 53513 15278 53517 15334
rect 53517 15278 53573 15334
rect 53573 15278 53577 15334
rect 53513 15274 53577 15278
rect 53513 15254 53577 15258
rect 53513 15198 53517 15254
rect 53517 15198 53573 15254
rect 53573 15198 53577 15254
rect 53513 15194 53577 15198
rect 53513 15174 53577 15178
rect 53513 15118 53517 15174
rect 53517 15118 53573 15174
rect 53573 15118 53577 15174
rect 53513 15114 53577 15118
rect 53513 15094 53577 15098
rect 53513 15038 53517 15094
rect 53517 15038 53573 15094
rect 53573 15038 53577 15094
rect 53513 15034 53577 15038
rect 53513 15014 53577 15018
rect 53513 14958 53517 15014
rect 53517 14958 53573 15014
rect 53573 14958 53577 15014
rect 53513 14954 53577 14958
rect 53513 14934 53577 14938
rect 53513 14878 53517 14934
rect 53517 14878 53573 14934
rect 53573 14878 53577 14934
rect 53513 14874 53577 14878
rect 53513 14854 53577 14858
rect 53513 14798 53517 14854
rect 53517 14798 53573 14854
rect 53573 14798 53577 14854
rect 53513 14794 53577 14798
rect 53513 14774 53577 14778
rect 53513 14718 53517 14774
rect 53517 14718 53573 14774
rect 53573 14718 53577 14774
rect 53513 14714 53577 14718
rect 53513 14694 53577 14698
rect 53513 14638 53517 14694
rect 53517 14638 53573 14694
rect 53573 14638 53577 14694
rect 53513 14634 53577 14638
rect 53513 14614 53577 14618
rect 53513 14558 53517 14614
rect 53517 14558 53573 14614
rect 53573 14558 53577 14614
rect 53513 14554 53577 14558
rect 53513 14534 53577 14538
rect 53513 14478 53517 14534
rect 53517 14478 53573 14534
rect 53573 14478 53577 14534
rect 53513 14474 53577 14478
rect 53513 14454 53577 14458
rect 53513 14398 53517 14454
rect 53517 14398 53573 14454
rect 53573 14398 53577 14454
rect 53513 14394 53577 14398
rect 53513 14374 53577 14378
rect 53513 14318 53517 14374
rect 53517 14318 53573 14374
rect 53573 14318 53577 14374
rect 53513 14314 53577 14318
rect 53513 14294 53577 14298
rect 53513 14238 53517 14294
rect 53517 14238 53573 14294
rect 53573 14238 53577 14294
rect 53513 14234 53577 14238
rect 53513 14214 53577 14218
rect 53513 14158 53517 14214
rect 53517 14158 53573 14214
rect 53573 14158 53577 14214
rect 53513 14154 53577 14158
rect 53513 14134 53577 14138
rect 53513 14078 53517 14134
rect 53517 14078 53573 14134
rect 53573 14078 53577 14134
rect 53513 14074 53577 14078
rect 53513 14054 53577 14058
rect 53513 13998 53517 14054
rect 53517 13998 53573 14054
rect 53573 13998 53577 14054
rect 53513 13994 53577 13998
rect 53513 13974 53577 13978
rect 53513 13918 53517 13974
rect 53517 13918 53573 13974
rect 53573 13918 53577 13974
rect 53513 13914 53577 13918
rect 56519 17167 56583 17171
rect 56519 17111 56523 17167
rect 56523 17111 56579 17167
rect 56579 17111 56583 17167
rect 56519 17107 56583 17111
rect 56519 17087 56583 17091
rect 56519 17031 56523 17087
rect 56523 17031 56579 17087
rect 56579 17031 56583 17087
rect 56519 17027 56583 17031
rect 56519 17007 56583 17011
rect 56519 16951 56523 17007
rect 56523 16951 56579 17007
rect 56579 16951 56583 17007
rect 56519 16947 56583 16951
rect 56519 16927 56583 16931
rect 56519 16871 56523 16927
rect 56523 16871 56579 16927
rect 56579 16871 56583 16927
rect 56519 16867 56583 16871
rect 56519 16847 56583 16851
rect 56519 16791 56523 16847
rect 56523 16791 56579 16847
rect 56579 16791 56583 16847
rect 56519 16787 56583 16791
rect 56519 16767 56583 16771
rect 56519 16711 56523 16767
rect 56523 16711 56579 16767
rect 56579 16711 56583 16767
rect 56519 16707 56583 16711
rect 56519 16687 56583 16691
rect 56519 16631 56523 16687
rect 56523 16631 56579 16687
rect 56579 16631 56583 16687
rect 56519 16627 56583 16631
rect 56519 16607 56583 16611
rect 56519 16551 56523 16607
rect 56523 16551 56579 16607
rect 56579 16551 56583 16607
rect 56519 16547 56583 16551
rect 56519 16527 56583 16531
rect 56519 16471 56523 16527
rect 56523 16471 56579 16527
rect 56579 16471 56583 16527
rect 56519 16467 56583 16471
rect 56519 16447 56583 16451
rect 56519 16391 56523 16447
rect 56523 16391 56579 16447
rect 56579 16391 56583 16447
rect 56519 16387 56583 16391
rect 56519 16367 56583 16371
rect 56519 16311 56523 16367
rect 56523 16311 56579 16367
rect 56579 16311 56583 16367
rect 56519 16307 56583 16311
rect 56519 16287 56583 16291
rect 56519 16231 56523 16287
rect 56523 16231 56579 16287
rect 56579 16231 56583 16287
rect 56519 16227 56583 16231
rect 56519 16207 56583 16211
rect 56519 16151 56523 16207
rect 56523 16151 56579 16207
rect 56579 16151 56583 16207
rect 56519 16147 56583 16151
rect 56519 16127 56583 16131
rect 56519 16071 56523 16127
rect 56523 16071 56579 16127
rect 56579 16071 56583 16127
rect 56519 16067 56583 16071
rect 56519 16047 56583 16051
rect 56519 15991 56523 16047
rect 56523 15991 56579 16047
rect 56579 15991 56583 16047
rect 56519 15987 56583 15991
rect 56519 15967 56583 15971
rect 56519 15911 56523 15967
rect 56523 15911 56579 15967
rect 56579 15911 56583 15967
rect 56519 15907 56583 15911
rect 56519 15887 56583 15891
rect 56519 15831 56523 15887
rect 56523 15831 56579 15887
rect 56579 15831 56583 15887
rect 56519 15827 56583 15831
rect 56519 15807 56583 15811
rect 56519 15751 56523 15807
rect 56523 15751 56579 15807
rect 56579 15751 56583 15807
rect 56519 15747 56583 15751
rect 56519 15727 56583 15731
rect 56519 15671 56523 15727
rect 56523 15671 56579 15727
rect 56579 15671 56583 15727
rect 56519 15667 56583 15671
rect 56519 15647 56583 15651
rect 56519 15591 56523 15647
rect 56523 15591 56579 15647
rect 56579 15591 56583 15647
rect 56519 15587 56583 15591
rect 56519 15567 56583 15571
rect 56519 15511 56523 15567
rect 56523 15511 56579 15567
rect 56579 15511 56583 15567
rect 56519 15507 56583 15511
rect 56519 15487 56583 15491
rect 56519 15431 56523 15487
rect 56523 15431 56579 15487
rect 56579 15431 56583 15487
rect 56519 15427 56583 15431
rect 56519 15407 56583 15411
rect 56519 15351 56523 15407
rect 56523 15351 56579 15407
rect 56579 15351 56583 15407
rect 56519 15347 56583 15351
rect 56519 15327 56583 15331
rect 56519 15271 56523 15327
rect 56523 15271 56579 15327
rect 56579 15271 56583 15327
rect 56519 15267 56583 15271
rect 56519 15247 56583 15251
rect 56519 15191 56523 15247
rect 56523 15191 56579 15247
rect 56579 15191 56583 15247
rect 56519 15187 56583 15191
rect 56519 15167 56583 15171
rect 56519 15111 56523 15167
rect 56523 15111 56579 15167
rect 56579 15111 56583 15167
rect 56519 15107 56583 15111
rect 56519 15087 56583 15091
rect 56519 15031 56523 15087
rect 56523 15031 56579 15087
rect 56579 15031 56583 15087
rect 56519 15027 56583 15031
rect 56519 15007 56583 15011
rect 56519 14951 56523 15007
rect 56523 14951 56579 15007
rect 56579 14951 56583 15007
rect 56519 14947 56583 14951
rect 56519 14927 56583 14931
rect 56519 14871 56523 14927
rect 56523 14871 56579 14927
rect 56579 14871 56583 14927
rect 56519 14867 56583 14871
rect 56519 14847 56583 14851
rect 56519 14791 56523 14847
rect 56523 14791 56579 14847
rect 56579 14791 56583 14847
rect 56519 14787 56583 14791
rect 56519 14767 56583 14771
rect 56519 14711 56523 14767
rect 56523 14711 56579 14767
rect 56579 14711 56583 14767
rect 56519 14707 56583 14711
rect 56519 14687 56583 14691
rect 56519 14631 56523 14687
rect 56523 14631 56579 14687
rect 56579 14631 56583 14687
rect 56519 14627 56583 14631
rect 56519 14607 56583 14611
rect 56519 14551 56523 14607
rect 56523 14551 56579 14607
rect 56579 14551 56583 14607
rect 56519 14547 56583 14551
rect 56519 14527 56583 14531
rect 56519 14471 56523 14527
rect 56523 14471 56579 14527
rect 56579 14471 56583 14527
rect 56519 14467 56583 14471
rect 56519 14447 56583 14451
rect 56519 14391 56523 14447
rect 56523 14391 56579 14447
rect 56579 14391 56583 14447
rect 56519 14387 56583 14391
rect 56519 14367 56583 14371
rect 56519 14311 56523 14367
rect 56523 14311 56579 14367
rect 56579 14311 56583 14367
rect 56519 14307 56583 14311
rect 56519 14287 56583 14291
rect 56519 14231 56523 14287
rect 56523 14231 56579 14287
rect 56579 14231 56583 14287
rect 56519 14227 56583 14231
rect 56519 14207 56583 14211
rect 56519 14151 56523 14207
rect 56523 14151 56579 14207
rect 56579 14151 56583 14207
rect 56519 14147 56583 14151
rect 56519 14127 56583 14131
rect 56519 14071 56523 14127
rect 56523 14071 56579 14127
rect 56579 14071 56583 14127
rect 56519 14067 56583 14071
rect 56519 14047 56583 14051
rect 56519 13991 56523 14047
rect 56523 13991 56579 14047
rect 56579 13991 56583 14047
rect 56519 13987 56583 13991
rect 56519 13967 56583 13971
rect 56519 13911 56523 13967
rect 56523 13911 56579 13967
rect 56579 13911 56583 13967
rect 56519 13907 56583 13911
<< metal4 >>
rect 1 112382 120001 112464
rect 1 110546 2083 112382
rect 3919 110546 13841 112382
rect 14397 110546 21841 112382
rect 22397 110546 29841 112382
rect 30397 110546 37841 112382
rect 38397 110546 45841 112382
rect 46397 110546 53841 112382
rect 54397 110546 61841 112382
rect 62397 110546 69841 112382
rect 70397 110546 77841 112382
rect 78397 110546 85841 112382
rect 86397 110546 93841 112382
rect 94397 110546 101841 112382
rect 102397 110546 112083 112382
rect 113919 110546 120001 112382
rect 1 110464 120001 110546
rect 1 108382 120001 108464
rect 1 106546 6083 108382
rect 7919 106546 17841 108382
rect 18397 106546 25841 108382
rect 26397 106546 33841 108382
rect 34397 106546 41841 108382
rect 42397 106546 49841 108382
rect 50397 106546 57841 108382
rect 58397 106546 65841 108382
rect 66397 106546 73841 108382
rect 74397 106546 81841 108382
rect 82397 106546 89841 108382
rect 90397 106546 97841 108382
rect 98397 106546 105841 108382
rect 106397 106546 116083 108382
rect 117919 106546 120001 108382
rect 1 106464 120001 106546
rect 40164 100714 40404 100828
rect 40164 100650 40263 100714
rect 40327 100650 40404 100714
rect 40164 100634 40404 100650
rect 40164 100570 40263 100634
rect 40327 100570 40404 100634
rect 40164 100554 40404 100570
rect 40164 100490 40263 100554
rect 40327 100490 40404 100554
rect 40164 100474 40404 100490
rect 40164 100410 40263 100474
rect 40327 100410 40404 100474
rect 40164 100394 40404 100410
rect 40164 100330 40263 100394
rect 40327 100330 40404 100394
rect 40164 100314 40404 100330
rect 40164 100250 40263 100314
rect 40327 100250 40404 100314
rect 40164 100234 40404 100250
rect 40164 100170 40263 100234
rect 40327 100170 40404 100234
rect 40164 100154 40404 100170
rect 40164 100090 40263 100154
rect 40327 100090 40404 100154
rect 40164 100074 40404 100090
rect 40164 100010 40263 100074
rect 40327 100010 40404 100074
rect 40164 99994 40404 100010
rect 40164 99930 40263 99994
rect 40327 99930 40404 99994
rect 40164 99914 40404 99930
rect 40164 99850 40263 99914
rect 40327 99850 40404 99914
rect 40164 99834 40404 99850
rect 40164 99770 40263 99834
rect 40327 99770 40404 99834
rect 40164 99754 40404 99770
rect 40164 99690 40263 99754
rect 40327 99690 40404 99754
rect 40164 99674 40404 99690
rect 40164 99610 40263 99674
rect 40327 99610 40404 99674
rect 40164 99594 40404 99610
rect 40164 99530 40263 99594
rect 40327 99530 40404 99594
rect 40164 99514 40404 99530
rect 40164 99450 40263 99514
rect 40327 99450 40404 99514
rect 40164 99434 40404 99450
rect 40164 99370 40263 99434
rect 40327 99370 40404 99434
rect 40164 99354 40404 99370
rect 40164 99290 40263 99354
rect 40327 99290 40404 99354
rect 40164 99274 40404 99290
rect 43180 100720 43420 100913
rect 43180 100656 43264 100720
rect 43328 100656 43420 100720
rect 43180 100640 43420 100656
rect 43180 100576 43264 100640
rect 43328 100576 43420 100640
rect 43180 100560 43420 100576
rect 43180 100496 43264 100560
rect 43328 100496 43420 100560
rect 43180 100480 43420 100496
rect 43180 100416 43264 100480
rect 43328 100416 43420 100480
rect 43180 100400 43420 100416
rect 43180 100336 43264 100400
rect 43328 100336 43420 100400
rect 43180 100320 43420 100336
rect 43180 100256 43264 100320
rect 43328 100256 43420 100320
rect 43180 100240 43420 100256
rect 43180 100176 43264 100240
rect 43328 100176 43420 100240
rect 43180 100160 43420 100176
rect 43180 100096 43264 100160
rect 43328 100096 43420 100160
rect 43180 100080 43420 100096
rect 43180 100016 43264 100080
rect 43328 100016 43420 100080
rect 43180 100000 43420 100016
rect 43180 99936 43264 100000
rect 43328 99936 43420 100000
rect 43180 99920 43420 99936
rect 43180 99856 43264 99920
rect 43328 99856 43420 99920
rect 43180 99840 43420 99856
rect 43180 99776 43264 99840
rect 43328 99776 43420 99840
rect 43180 99760 43420 99776
rect 43180 99696 43264 99760
rect 43328 99696 43420 99760
rect 43180 99680 43420 99696
rect 43180 99616 43264 99680
rect 43328 99616 43420 99680
rect 43180 99600 43420 99616
rect 43180 99536 43264 99600
rect 43328 99536 43420 99600
rect 43180 99520 43420 99536
rect 43180 99456 43264 99520
rect 43328 99456 43420 99520
rect 43180 99440 43420 99456
rect 43180 99376 43264 99440
rect 43328 99376 43420 99440
rect 43180 99360 43420 99376
rect 43180 99296 43264 99360
rect 43328 99296 43420 99360
rect 43180 99280 43420 99296
rect 43180 99275 43264 99280
rect 40164 99210 40263 99274
rect 40327 99210 40404 99274
rect 40164 99194 40404 99210
rect 40164 99130 40263 99194
rect 40327 99130 40404 99194
rect 40164 99114 40404 99130
rect 40164 99090 40263 99114
rect 37853 99088 40263 99090
rect 37853 98852 38000 99088
rect 38236 99050 40263 99088
rect 40327 99050 40404 99114
rect 38236 99034 40404 99050
rect 41851 99273 43264 99275
rect 41851 99037 41998 99273
rect 42234 99216 43264 99273
rect 43328 99216 43420 99280
rect 42234 99200 43420 99216
rect 42234 99136 43264 99200
rect 43328 99136 43420 99200
rect 68177 100716 68417 100900
rect 68177 100652 68269 100716
rect 68333 100652 68417 100716
rect 68177 100636 68417 100652
rect 68177 100572 68269 100636
rect 68333 100572 68417 100636
rect 68177 100556 68417 100572
rect 68177 100492 68269 100556
rect 68333 100492 68417 100556
rect 68177 100476 68417 100492
rect 68177 100412 68269 100476
rect 68333 100412 68417 100476
rect 68177 100396 68417 100412
rect 68177 100332 68269 100396
rect 68333 100332 68417 100396
rect 68177 100316 68417 100332
rect 68177 100252 68269 100316
rect 68333 100252 68417 100316
rect 68177 100236 68417 100252
rect 68177 100172 68269 100236
rect 68333 100172 68417 100236
rect 68177 100156 68417 100172
rect 68177 100092 68269 100156
rect 68333 100092 68417 100156
rect 68177 100076 68417 100092
rect 68177 100012 68269 100076
rect 68333 100012 68417 100076
rect 68177 99996 68417 100012
rect 68177 99932 68269 99996
rect 68333 99932 68417 99996
rect 68177 99916 68417 99932
rect 68177 99852 68269 99916
rect 68333 99852 68417 99916
rect 68177 99836 68417 99852
rect 68177 99772 68269 99836
rect 68333 99772 68417 99836
rect 68177 99756 68417 99772
rect 68177 99692 68269 99756
rect 68333 99692 68417 99756
rect 68177 99676 68417 99692
rect 68177 99612 68269 99676
rect 68333 99612 68417 99676
rect 68177 99596 68417 99612
rect 68177 99532 68269 99596
rect 68333 99532 68417 99596
rect 68177 99516 68417 99532
rect 68177 99452 68269 99516
rect 68333 99452 68417 99516
rect 68177 99436 68417 99452
rect 68177 99372 68269 99436
rect 68333 99372 68417 99436
rect 68177 99356 68417 99372
rect 68177 99292 68269 99356
rect 68333 99292 68417 99356
rect 68177 99276 68417 99292
rect 68177 99212 68269 99276
rect 68333 99212 68417 99276
rect 68177 99196 68417 99212
rect 68177 99194 68269 99196
rect 42234 99120 43420 99136
rect 42234 99056 43264 99120
rect 43328 99056 43420 99120
rect 42234 99040 43420 99056
rect 42234 99037 43264 99040
rect 41851 99035 43264 99037
rect 38236 98970 40263 99034
rect 40327 98970 40404 99034
rect 38236 98954 40404 98970
rect 38236 98890 40263 98954
rect 40327 98890 40404 98954
rect 38236 98874 40404 98890
rect 38236 98852 40263 98874
rect 37853 98850 40263 98852
rect 40164 98810 40263 98850
rect 40327 98810 40404 98874
rect 40164 98794 40404 98810
rect 40164 98730 40263 98794
rect 40327 98730 40404 98794
rect 40164 98714 40404 98730
rect 40164 98650 40263 98714
rect 40327 98650 40404 98714
rect 40164 98634 40404 98650
rect 40164 98570 40263 98634
rect 40327 98570 40404 98634
rect 40164 98554 40404 98570
rect 40164 98490 40263 98554
rect 40327 98490 40404 98554
rect 40164 98474 40404 98490
rect 40164 98410 40263 98474
rect 40327 98410 40404 98474
rect 40164 98394 40404 98410
rect 40164 98330 40263 98394
rect 40327 98330 40404 98394
rect 40164 98314 40404 98330
rect 40164 98250 40263 98314
rect 40327 98250 40404 98314
rect 40164 98234 40404 98250
rect 40164 98170 40263 98234
rect 40327 98170 40404 98234
rect 40164 98154 40404 98170
rect 40164 98090 40263 98154
rect 40327 98090 40404 98154
rect 40164 98074 40404 98090
rect 40164 98010 40263 98074
rect 40327 98010 40404 98074
rect 40164 97994 40404 98010
rect 40164 97930 40263 97994
rect 40327 97930 40404 97994
rect 40164 97914 40404 97930
rect 40164 97850 40263 97914
rect 40327 97850 40404 97914
rect 40164 97834 40404 97850
rect 40164 97770 40263 97834
rect 40327 97770 40404 97834
rect 40164 97754 40404 97770
rect 40164 97690 40263 97754
rect 40327 97690 40404 97754
rect 40164 97674 40404 97690
rect 40164 97610 40263 97674
rect 40327 97610 40404 97674
rect 40164 97594 40404 97610
rect 40164 97530 40263 97594
rect 40327 97530 40404 97594
rect 40164 97514 40404 97530
rect 40164 97450 40263 97514
rect 40327 97450 40404 97514
rect 40164 96581 40404 97450
rect 43180 98976 43264 99035
rect 43328 98976 43420 99040
rect 43180 98960 43420 98976
rect 43180 98896 43264 98960
rect 43328 98896 43420 98960
rect 68176 99132 68269 99194
rect 68333 99194 68417 99196
rect 71177 100729 71417 100898
rect 71177 100665 71270 100729
rect 71334 100665 71417 100729
rect 71177 100649 71417 100665
rect 71177 100585 71270 100649
rect 71334 100585 71417 100649
rect 71177 100569 71417 100585
rect 71177 100505 71270 100569
rect 71334 100505 71417 100569
rect 71177 100489 71417 100505
rect 71177 100425 71270 100489
rect 71334 100425 71417 100489
rect 71177 100409 71417 100425
rect 71177 100345 71270 100409
rect 71334 100345 71417 100409
rect 71177 100329 71417 100345
rect 71177 100265 71270 100329
rect 71334 100265 71417 100329
rect 71177 100249 71417 100265
rect 71177 100185 71270 100249
rect 71334 100185 71417 100249
rect 71177 100169 71417 100185
rect 71177 100105 71270 100169
rect 71334 100105 71417 100169
rect 71177 100089 71417 100105
rect 71177 100025 71270 100089
rect 71334 100025 71417 100089
rect 71177 100009 71417 100025
rect 71177 99945 71270 100009
rect 71334 99945 71417 100009
rect 71177 99929 71417 99945
rect 71177 99865 71270 99929
rect 71334 99865 71417 99929
rect 71177 99849 71417 99865
rect 71177 99785 71270 99849
rect 71334 99785 71417 99849
rect 71177 99769 71417 99785
rect 71177 99705 71270 99769
rect 71334 99705 71417 99769
rect 71177 99689 71417 99705
rect 71177 99625 71270 99689
rect 71334 99625 71417 99689
rect 71177 99609 71417 99625
rect 71177 99545 71270 99609
rect 71334 99545 71417 99609
rect 71177 99529 71417 99545
rect 71177 99465 71270 99529
rect 71334 99465 71417 99529
rect 71177 99449 71417 99465
rect 71177 99385 71270 99449
rect 71334 99385 71417 99449
rect 71177 99369 71417 99385
rect 71177 99305 71270 99369
rect 71334 99305 71417 99369
rect 71177 99289 71417 99305
rect 71177 99225 71270 99289
rect 71334 99225 71417 99289
rect 71177 99209 71417 99225
rect 68333 99192 70382 99194
rect 68333 99132 69999 99192
rect 68176 99116 69999 99132
rect 68176 99052 68269 99116
rect 68333 99052 69999 99116
rect 68176 99036 69999 99052
rect 68176 98972 68269 99036
rect 68333 98972 69999 99036
rect 68176 98956 69999 98972
rect 70235 98956 70382 99192
rect 68176 98954 68269 98956
rect 43180 98880 43420 98896
rect 43180 98816 43264 98880
rect 43328 98816 43420 98880
rect 43180 98800 43420 98816
rect 43180 98736 43264 98800
rect 43328 98736 43420 98800
rect 43180 98720 43420 98736
rect 43180 98656 43264 98720
rect 43328 98656 43420 98720
rect 43180 98640 43420 98656
rect 43180 98576 43264 98640
rect 43328 98576 43420 98640
rect 43180 98560 43420 98576
rect 43180 98496 43264 98560
rect 43328 98496 43420 98560
rect 43180 98480 43420 98496
rect 43180 98416 43264 98480
rect 43328 98416 43420 98480
rect 43180 98400 43420 98416
rect 43180 98336 43264 98400
rect 43328 98336 43420 98400
rect 43180 98320 43420 98336
rect 43180 98256 43264 98320
rect 43328 98256 43420 98320
rect 43180 98240 43420 98256
rect 43180 98176 43264 98240
rect 43328 98176 43420 98240
rect 43180 98160 43420 98176
rect 43180 98096 43264 98160
rect 43328 98096 43420 98160
rect 43180 98080 43420 98096
rect 43180 98016 43264 98080
rect 43328 98016 43420 98080
rect 43180 98000 43420 98016
rect 43180 97936 43264 98000
rect 43328 97936 43420 98000
rect 43180 97920 43420 97936
rect 43180 97856 43264 97920
rect 43328 97856 43420 97920
rect 43180 97840 43420 97856
rect 43180 97776 43264 97840
rect 43328 97776 43420 97840
rect 43180 97760 43420 97776
rect 43180 97696 43264 97760
rect 43328 97696 43420 97760
rect 43180 97680 43420 97696
rect 43180 97616 43264 97680
rect 43328 97616 43420 97680
rect 43180 97600 43420 97616
rect 43180 97536 43264 97600
rect 43328 97536 43420 97600
rect 43180 97520 43420 97536
rect 43180 97456 43264 97520
rect 43328 97456 43420 97520
rect 43180 97264 43420 97456
rect 68177 98892 68269 98954
rect 68333 98954 70382 98956
rect 71177 99145 71270 99209
rect 71334 99186 71417 99209
rect 71334 99184 74381 99186
rect 71334 99145 73998 99184
rect 71177 99129 73998 99145
rect 71177 99065 71270 99129
rect 71334 99065 73998 99129
rect 71177 99049 73998 99065
rect 71177 98985 71270 99049
rect 71334 98985 73998 99049
rect 71177 98969 73998 98985
rect 68333 98892 68417 98954
rect 68177 98876 68417 98892
rect 68177 98812 68269 98876
rect 68333 98812 68417 98876
rect 68177 98796 68417 98812
rect 68177 98732 68269 98796
rect 68333 98732 68417 98796
rect 68177 98716 68417 98732
rect 68177 98652 68269 98716
rect 68333 98652 68417 98716
rect 68177 98636 68417 98652
rect 68177 98572 68269 98636
rect 68333 98572 68417 98636
rect 68177 98556 68417 98572
rect 68177 98492 68269 98556
rect 68333 98492 68417 98556
rect 68177 98476 68417 98492
rect 68177 98412 68269 98476
rect 68333 98412 68417 98476
rect 68177 98396 68417 98412
rect 68177 98332 68269 98396
rect 68333 98332 68417 98396
rect 68177 98316 68417 98332
rect 68177 98252 68269 98316
rect 68333 98252 68417 98316
rect 68177 98236 68417 98252
rect 68177 98172 68269 98236
rect 68333 98172 68417 98236
rect 68177 98156 68417 98172
rect 68177 98092 68269 98156
rect 68333 98092 68417 98156
rect 68177 98076 68417 98092
rect 68177 98012 68269 98076
rect 68333 98012 68417 98076
rect 68177 97996 68417 98012
rect 68177 97932 68269 97996
rect 68333 97932 68417 97996
rect 68177 97916 68417 97932
rect 68177 97852 68269 97916
rect 68333 97852 68417 97916
rect 68177 97836 68417 97852
rect 68177 97772 68269 97836
rect 68333 97772 68417 97836
rect 68177 97756 68417 97772
rect 68177 97692 68269 97756
rect 68333 97692 68417 97756
rect 68177 97676 68417 97692
rect 68177 97612 68269 97676
rect 68333 97612 68417 97676
rect 68177 97596 68417 97612
rect 68177 97532 68269 97596
rect 68333 97532 68417 97596
rect 68177 97516 68417 97532
rect 68177 97452 68269 97516
rect 68333 97452 68417 97516
rect 68177 97266 68417 97452
rect 71177 98905 71270 98969
rect 71334 98948 73998 98969
rect 74234 98948 74381 99184
rect 71334 98946 74381 98948
rect 71334 98905 71417 98946
rect 71177 98889 71417 98905
rect 71177 98825 71270 98889
rect 71334 98825 71417 98889
rect 71177 98809 71417 98825
rect 71177 98745 71270 98809
rect 71334 98745 71417 98809
rect 71177 98729 71417 98745
rect 71177 98665 71270 98729
rect 71334 98665 71417 98729
rect 71177 98649 71417 98665
rect 71177 98585 71270 98649
rect 71334 98585 71417 98649
rect 71177 98569 71417 98585
rect 71177 98505 71270 98569
rect 71334 98505 71417 98569
rect 71177 98489 71417 98505
rect 71177 98425 71270 98489
rect 71334 98425 71417 98489
rect 71177 98409 71417 98425
rect 71177 98345 71270 98409
rect 71334 98345 71417 98409
rect 71177 98329 71417 98345
rect 71177 98265 71270 98329
rect 71334 98265 71417 98329
rect 71177 98249 71417 98265
rect 71177 98185 71270 98249
rect 71334 98185 71417 98249
rect 71177 98169 71417 98185
rect 71177 98105 71270 98169
rect 71334 98105 71417 98169
rect 71177 98089 71417 98105
rect 71177 98025 71270 98089
rect 71334 98025 71417 98089
rect 71177 98009 71417 98025
rect 71177 97945 71270 98009
rect 71334 97945 71417 98009
rect 71177 97929 71417 97945
rect 71177 97865 71270 97929
rect 71334 97865 71417 97929
rect 71177 97849 71417 97865
rect 71177 97785 71270 97849
rect 71334 97785 71417 97849
rect 71177 97769 71417 97785
rect 71177 97705 71270 97769
rect 71334 97705 71417 97769
rect 71177 97689 71417 97705
rect 71177 97625 71270 97689
rect 71334 97625 71417 97689
rect 71177 97609 71417 97625
rect 71177 97545 71270 97609
rect 71334 97545 71417 97609
rect 71177 97529 71417 97545
rect 71177 97465 71270 97529
rect 71334 97465 71417 97529
rect 71177 97254 71417 97465
rect 40164 96517 43023 96581
rect 40429 95824 40495 95825
rect 40429 95760 40430 95824
rect 40494 95760 40495 95824
rect 41608 95821 41672 96517
rect 41824 95827 41890 95828
rect 40429 95759 40495 95760
rect 41607 95820 41673 95821
rect 40430 94920 40494 95759
rect 41607 95756 41608 95820
rect 41672 95756 41673 95820
rect 41824 95763 41825 95827
rect 41889 95763 41890 95827
rect 42959 95825 43023 96517
rect 41824 95762 41890 95763
rect 42958 95824 43024 95825
rect 41607 95755 41673 95756
rect 41825 95016 41889 95762
rect 42958 95760 42959 95824
rect 43023 95760 43024 95824
rect 42958 95759 43024 95760
rect 41825 95014 42382 95016
rect 41825 94920 41999 95014
rect 40430 94856 41999 94920
rect 40430 94325 40494 94856
rect 41852 94778 41999 94856
rect 42235 94778 42382 95014
rect 41852 94776 42382 94778
rect 40430 94320 40605 94325
rect 37853 94257 38429 94259
rect 37853 94021 38000 94257
rect 38236 94165 38429 94257
rect 40430 94256 40540 94320
rect 40604 94256 40605 94320
rect 41867 94308 41931 94776
rect 41866 94307 41932 94308
rect 40539 94255 40605 94256
rect 41653 94306 41719 94307
rect 41653 94242 41654 94306
rect 41718 94242 41719 94306
rect 41866 94243 41867 94307
rect 41931 94243 41932 94307
rect 41866 94242 41932 94243
rect 43030 94307 43096 94308
rect 43030 94243 43031 94307
rect 43095 94243 43096 94307
rect 43030 94242 43096 94243
rect 41653 94241 41719 94242
rect 41654 94165 41718 94241
rect 43031 94165 43095 94242
rect 38236 94101 43095 94165
rect 38236 94021 38429 94101
rect 37853 94019 38429 94021
rect 93724 93356 93790 93357
rect 93724 93292 93725 93356
rect 93789 93292 93790 93356
rect 93724 93280 93790 93292
rect 41855 92935 42385 92937
rect 41855 92829 42002 92935
rect 40517 92765 42002 92829
rect 40517 91636 40581 92765
rect 41132 92284 41196 92765
rect 41855 92699 42002 92765
rect 42238 92829 42385 92935
rect 42238 92765 42854 92829
rect 42238 92699 42385 92765
rect 41855 92697 42385 92699
rect 41672 92538 41736 92564
rect 41671 92514 41737 92538
rect 41671 92450 41672 92514
rect 41736 92450 41737 92514
rect 41671 92434 41737 92450
rect 41671 92370 41672 92434
rect 41736 92370 41737 92434
rect 41671 92354 41737 92370
rect 41671 92290 41672 92354
rect 41736 92290 41737 92354
rect 41130 92277 41205 92284
rect 41130 92213 41135 92277
rect 41199 92213 41205 92277
rect 41130 92197 41205 92213
rect 41130 92133 41135 92197
rect 41199 92133 41205 92197
rect 41671 92274 41737 92290
rect 42220 92287 42284 92697
rect 41671 92210 41672 92274
rect 41736 92210 41737 92274
rect 41671 92187 41737 92210
rect 42214 92280 42289 92287
rect 42214 92216 42219 92280
rect 42283 92216 42289 92280
rect 42214 92200 42289 92216
rect 41130 92126 41205 92133
rect 40516 91635 40582 91636
rect 40516 91571 40517 91635
rect 40581 91571 40582 91635
rect 41672 91630 41736 92187
rect 42214 92136 42219 92200
rect 42283 92136 42289 92200
rect 42214 92129 42289 92136
rect 42790 91641 42854 92765
rect 93158 92763 93226 92765
rect 93158 92699 93160 92763
rect 93224 92699 93226 92763
rect 93158 92697 93226 92699
rect 93159 92660 93225 92697
rect 92569 92103 92637 92105
rect 92569 92039 92571 92103
rect 92635 92039 92637 92103
rect 92569 92037 92637 92039
rect 42789 91640 42855 91641
rect 40516 91570 40582 91571
rect 41671 91629 41737 91630
rect 41671 91565 41672 91629
rect 41736 91565 41737 91629
rect 42789 91576 42790 91640
rect 42854 91576 42855 91640
rect 42789 91575 42855 91576
rect 41671 91564 41737 91565
rect 37849 91142 38379 91144
rect 37849 90906 37996 91142
rect 38232 91052 38379 91142
rect 41672 91052 41736 91564
rect 38232 90988 41736 91052
rect 38232 90906 38379 90988
rect 37849 90904 38379 90906
rect 43998 90792 44062 90794
rect 43997 90791 44063 90792
rect 43997 90727 43998 90791
rect 44062 90727 44063 90791
rect 43997 90726 44063 90727
rect 49020 90791 49086 90792
rect 49020 90727 49021 90791
rect 49085 90727 49086 90791
rect 49020 90726 49086 90727
rect 43998 83603 44062 90726
rect 44778 90468 44844 90469
rect 44778 90404 44779 90468
rect 44843 90404 44844 90468
rect 44778 90403 44844 90404
rect 44779 83603 44843 90403
rect 45789 90036 45853 90040
rect 45788 90035 45854 90036
rect 45788 89971 45789 90035
rect 45853 89971 45854 90035
rect 45788 89970 45854 89971
rect 45789 83603 45853 89970
rect 46558 89783 46622 89790
rect 46557 89782 46623 89783
rect 46557 89718 46558 89782
rect 46622 89718 46623 89782
rect 46557 89717 46623 89718
rect 46022 87555 46358 87580
rect 46022 87251 46038 87555
rect 46342 87251 46358 87555
rect 46022 87226 46358 87251
rect 46558 83603 46622 89717
rect 49021 89352 49085 90726
rect 49827 90468 49893 90469
rect 49827 90404 49828 90468
rect 49892 90404 49893 90468
rect 49827 90403 49893 90404
rect 49020 89351 49086 89352
rect 49020 89287 49021 89351
rect 49085 89287 49086 89351
rect 49020 89286 49086 89287
rect 49828 89099 49892 90403
rect 54420 90035 54486 90036
rect 54420 89971 54421 90035
rect 54485 89971 54486 90035
rect 54420 89970 54486 89971
rect 54421 89352 54485 89970
rect 55227 89782 55293 89783
rect 55227 89718 55228 89782
rect 55292 89718 55293 89782
rect 55227 89717 55293 89718
rect 54420 89351 54486 89352
rect 54420 89287 54421 89351
rect 54485 89287 54495 89351
rect 54420 89286 54486 89287
rect 55228 89099 55292 89717
rect 49827 89098 49893 89099
rect 49827 89034 49828 89098
rect 49892 89034 49893 89098
rect 49827 89033 49893 89034
rect 55227 89098 55293 89099
rect 55227 89034 55228 89098
rect 55292 89034 55303 89098
rect 55227 89033 55293 89034
rect 73811 88750 90426 88789
rect 73811 88686 74525 88750
rect 74589 88686 81053 88750
rect 81117 88686 88669 88750
rect 88733 88686 90426 88750
rect 73811 88670 90426 88686
rect 73811 88606 74525 88670
rect 74589 88606 81053 88670
rect 81117 88606 88669 88670
rect 88733 88606 90426 88670
rect 73811 88601 90426 88606
rect 73811 88595 85995 88601
rect 73811 88590 78001 88595
rect 73811 88526 74525 88590
rect 74589 88526 78001 88590
rect 73811 88510 78001 88526
rect 73811 88446 74525 88510
rect 74589 88446 78001 88510
rect 73811 88430 78001 88446
rect 73811 88366 74525 88430
rect 74589 88366 78001 88430
rect 73811 88359 78001 88366
rect 78237 88590 85995 88595
rect 78237 88526 81053 88590
rect 81117 88526 85995 88590
rect 78237 88510 85995 88526
rect 78237 88446 81053 88510
rect 81117 88446 85995 88510
rect 78237 88430 85995 88446
rect 78237 88366 81053 88430
rect 81117 88366 85995 88430
rect 78237 88365 85995 88366
rect 86231 88590 90426 88601
rect 86231 88526 88669 88590
rect 88733 88526 90426 88590
rect 86231 88510 90426 88526
rect 86231 88446 88669 88510
rect 88733 88446 90426 88510
rect 86231 88430 90426 88446
rect 86231 88366 88669 88430
rect 88733 88366 90426 88430
rect 86231 88365 90426 88366
rect 78237 88359 90426 88365
rect 73811 88350 90426 88359
rect 73811 88286 74525 88350
rect 74589 88286 81053 88350
rect 81117 88286 88669 88350
rect 88733 88286 90426 88350
rect 73811 88270 90426 88286
rect 73811 88206 74525 88270
rect 74589 88206 81053 88270
rect 81117 88206 88669 88270
rect 88733 88206 90426 88270
rect 73811 88169 90426 88206
rect 53853 87431 54383 87433
rect 49020 87426 49464 87427
rect 46906 87424 46972 87425
rect 47209 87424 47653 87425
rect 49020 87424 49050 87426
rect 46906 87360 46907 87424
rect 46971 87360 47239 87424
rect 47303 87360 47319 87424
rect 47383 87360 47399 87424
rect 47463 87360 47479 87424
rect 47543 87360 47559 87424
rect 47623 87362 49050 87424
rect 49114 87362 49130 87426
rect 49194 87362 49210 87426
rect 49274 87362 49290 87426
rect 49354 87362 49370 87426
rect 49434 87424 49464 87426
rect 53853 87424 54000 87431
rect 49434 87422 54000 87424
rect 49434 87362 50845 87422
rect 47623 87360 50845 87362
rect 46906 87359 46972 87360
rect 47209 87359 47653 87360
rect 50815 87358 50845 87360
rect 50909 87358 50925 87422
rect 50989 87358 51005 87422
rect 51069 87358 51085 87422
rect 51149 87358 51165 87422
rect 51229 87420 54000 87422
rect 51229 87360 52644 87420
rect 51229 87358 51259 87360
rect 50815 87357 51259 87358
rect 52614 87356 52644 87360
rect 52708 87356 52724 87420
rect 52788 87356 52804 87420
rect 52868 87356 52884 87420
rect 52948 87356 52964 87420
rect 53028 87360 54000 87420
rect 53028 87356 53058 87360
rect 52614 87355 53058 87356
rect 50154 87226 50396 87229
rect 50154 86990 50157 87226
rect 50393 86990 50396 87226
rect 53853 87195 54000 87360
rect 54236 87425 54383 87431
rect 54236 87424 54849 87425
rect 54236 87360 54435 87424
rect 54499 87360 54515 87424
rect 54579 87360 54595 87424
rect 54659 87360 54675 87424
rect 54739 87360 54755 87424
rect 54819 87420 57337 87424
rect 54819 87360 56237 87420
rect 54236 87359 54849 87360
rect 54236 87195 54383 87359
rect 56207 87356 56237 87360
rect 56301 87356 56317 87420
rect 56381 87356 56397 87420
rect 56461 87356 56477 87420
rect 56541 87356 56557 87420
rect 56621 87360 57337 87420
rect 56621 87356 56651 87360
rect 56207 87355 56651 87356
rect 53853 87193 54383 87195
rect 57850 87252 58382 87255
rect 57850 87246 57998 87252
rect 58234 87246 58382 87252
rect 57850 87022 57884 87246
rect 58348 87022 58382 87246
rect 57850 87016 57998 87022
rect 58234 87016 58382 87022
rect 57850 87013 58382 87016
rect 50154 86987 50396 86990
rect 73809 86747 90321 86789
rect 73809 86683 75070 86747
rect 75134 86683 76158 86747
rect 76222 86683 78334 86747
rect 78398 86683 79422 86747
rect 79486 86683 80510 86747
rect 80574 86683 81598 86747
rect 81662 86683 82686 86747
rect 82750 86683 83774 86747
rect 83838 86683 85950 86747
rect 86014 86683 87038 86747
rect 87102 86683 88126 86747
rect 88190 86739 90321 86747
rect 88190 86683 90384 86739
rect 73809 86667 90384 86683
rect 73809 86604 75070 86667
rect 73809 86368 74004 86604
rect 74240 86603 75070 86604
rect 75134 86603 76158 86667
rect 76222 86603 78334 86667
rect 78398 86603 79422 86667
rect 79486 86603 80510 86667
rect 80574 86603 81598 86667
rect 81662 86603 82686 86667
rect 82750 86603 83774 86667
rect 83838 86603 85950 86667
rect 86014 86603 87038 86667
rect 87102 86603 88126 86667
rect 88190 86603 90384 86667
rect 74240 86597 90384 86603
rect 74240 86587 82000 86597
rect 74240 86523 75070 86587
rect 75134 86523 76158 86587
rect 76222 86523 78334 86587
rect 78398 86523 79422 86587
rect 79486 86523 80510 86587
rect 80574 86523 81598 86587
rect 81662 86523 82000 86587
rect 74240 86507 82000 86523
rect 74240 86443 75070 86507
rect 75134 86443 76158 86507
rect 76222 86443 78334 86507
rect 78398 86443 79422 86507
rect 79486 86443 80510 86507
rect 80574 86443 81598 86507
rect 81662 86443 82000 86507
rect 74240 86427 82000 86443
rect 74240 86368 75070 86427
rect 73809 86363 75070 86368
rect 75134 86363 76158 86427
rect 76222 86363 78334 86427
rect 78398 86363 79422 86427
rect 79486 86363 80510 86427
rect 80574 86363 81598 86427
rect 81662 86363 82000 86427
rect 73809 86361 82000 86363
rect 82236 86593 90384 86597
rect 82236 86587 90003 86593
rect 82236 86523 82686 86587
rect 82750 86523 83774 86587
rect 83838 86523 85950 86587
rect 86014 86523 87038 86587
rect 87102 86523 88126 86587
rect 88190 86523 90003 86587
rect 82236 86507 90003 86523
rect 82236 86443 82686 86507
rect 82750 86443 83774 86507
rect 83838 86443 85950 86507
rect 86014 86443 87038 86507
rect 87102 86443 88126 86507
rect 88190 86443 90003 86507
rect 82236 86427 90003 86443
rect 82236 86363 82686 86427
rect 82750 86363 83774 86427
rect 83838 86363 85950 86427
rect 86014 86363 87038 86427
rect 87102 86363 88126 86427
rect 88190 86363 90003 86427
rect 82236 86361 90003 86363
rect 73809 86357 90003 86361
rect 90239 86357 90384 86593
rect 73809 86347 90384 86357
rect 73809 86283 75070 86347
rect 75134 86283 76158 86347
rect 76222 86283 78334 86347
rect 78398 86283 79422 86347
rect 79486 86283 80510 86347
rect 80574 86283 81598 86347
rect 81662 86283 82686 86347
rect 82750 86283 83774 86347
rect 83838 86283 85950 86347
rect 86014 86283 87038 86347
rect 87102 86283 88126 86347
rect 88190 86283 90384 86347
rect 73809 86267 90384 86283
rect 73809 86203 75070 86267
rect 75134 86203 76158 86267
rect 76222 86203 78334 86267
rect 78398 86203 79422 86267
rect 79486 86203 80510 86267
rect 80574 86203 81598 86267
rect 81662 86203 82686 86267
rect 82750 86203 83774 86267
rect 83838 86203 85950 86267
rect 86014 86203 87038 86267
rect 87102 86203 88126 86267
rect 88190 86211 90384 86267
rect 88190 86203 90321 86211
rect 73809 86169 90321 86203
rect 43625 83539 44062 83603
rect 37856 74710 38386 74712
rect 37856 74474 38003 74710
rect 38239 74474 38386 74710
rect 37856 74472 38386 74474
rect 29858 73846 30388 73848
rect 29858 73610 30005 73846
rect 30241 73742 30388 73846
rect 30268 73678 30284 73742
rect 30348 73678 30388 73742
rect 30241 73610 30388 73678
rect 29858 73608 30388 73610
rect 30969 73243 34390 73245
rect 30969 73200 34007 73243
rect 30969 73136 31130 73200
rect 31194 73136 31210 73200
rect 31274 73136 31290 73200
rect 31354 73136 31370 73200
rect 31434 73136 34007 73200
rect 30969 73007 34007 73136
rect 34243 73007 34390 73243
rect 30969 73005 34390 73007
rect 29932 67300 30172 67395
rect 29932 67236 30023 67300
rect 30087 67236 30172 67300
rect 29932 67220 30172 67236
rect 29932 67156 30023 67220
rect 30087 67178 30172 67220
rect 30087 67176 30385 67178
rect 29932 67140 30040 67156
rect 29932 67076 30023 67140
rect 29932 67060 30040 67076
rect 29932 66996 30023 67060
rect 29932 66980 30040 66996
rect 29932 66916 30023 66980
rect 30276 66940 30385 67176
rect 43625 67084 43689 83539
rect 43998 76413 44062 83539
rect 44401 83539 44843 83603
rect 43997 76412 44063 76413
rect 43997 76348 43998 76412
rect 44062 76348 44063 76412
rect 43997 76347 44063 76348
rect 43624 67083 43690 67084
rect 43624 67019 43625 67083
rect 43689 67019 43690 67083
rect 43624 67018 43690 67019
rect 43625 67014 43689 67018
rect 30087 66938 30385 66940
rect 30087 66916 30172 66938
rect 29932 66900 30172 66916
rect 29932 66836 30023 66900
rect 30087 66836 30172 66900
rect 29932 66159 30172 66836
rect 44401 66421 44465 83539
rect 44779 76736 44843 83539
rect 45381 83539 45853 83603
rect 44778 76735 44844 76736
rect 44778 76671 44779 76735
rect 44843 76671 44844 76735
rect 44778 76670 44844 76671
rect 45381 68628 45445 83539
rect 45789 77169 45853 83539
rect 46189 83539 46622 83603
rect 45788 77168 45854 77169
rect 45788 77104 45789 77168
rect 45853 77104 45854 77168
rect 45788 77103 45854 77104
rect 45732 71278 45798 71279
rect 45732 71214 45733 71278
rect 45797 71214 45798 71278
rect 45732 71213 45798 71214
rect 45733 68628 45797 71213
rect 45381 68564 45797 68628
rect 46189 68641 46253 83539
rect 46558 77425 46622 83539
rect 57438 84828 57734 84909
rect 50116 79351 50388 79419
rect 50116 79115 50134 79351
rect 50370 79115 50388 79351
rect 50116 79031 50388 79115
rect 50116 78795 50134 79031
rect 50370 78795 50388 79031
rect 50116 78728 50388 78795
rect 50229 78619 50293 78728
rect 50227 78618 50293 78619
rect 48536 78617 48602 78618
rect 50227 78617 50228 78618
rect 48536 78553 48537 78617
rect 48601 78554 50228 78617
rect 50292 78617 50293 78618
rect 51932 78617 51998 78618
rect 53728 78617 53794 78618
rect 55557 78617 55623 78618
rect 50292 78554 51933 78617
rect 48601 78553 51933 78554
rect 51997 78553 53729 78617
rect 53793 78553 55558 78617
rect 55622 78553 57334 78617
rect 48536 78552 48602 78553
rect 51932 78552 51998 78553
rect 53728 78552 53794 78553
rect 55557 78552 55623 78553
rect 53857 78442 54387 78444
rect 50984 78426 51228 78427
rect 47389 78425 47633 78426
rect 50984 78425 50994 78426
rect 47363 78361 47399 78425
rect 47463 78361 47479 78425
rect 47543 78361 47559 78425
rect 47623 78424 50994 78425
rect 47623 78361 49194 78424
rect 47389 78360 47633 78361
rect 49184 78360 49194 78361
rect 49258 78360 49274 78424
rect 49338 78360 49354 78424
rect 49418 78362 50994 78424
rect 51058 78362 51074 78426
rect 51138 78362 51154 78426
rect 51218 78425 51228 78426
rect 52782 78425 53026 78426
rect 53857 78425 54004 78442
rect 51218 78362 52792 78425
rect 49418 78361 52792 78362
rect 52856 78361 52872 78425
rect 52936 78361 52952 78425
rect 53016 78361 54004 78425
rect 49418 78360 49428 78361
rect 52782 78360 53026 78361
rect 49184 78359 49428 78360
rect 53857 78206 54004 78361
rect 54240 78425 54387 78442
rect 57270 78427 57334 78553
rect 54580 78426 54824 78427
rect 57269 78426 57335 78427
rect 54580 78425 54590 78426
rect 54240 78362 54590 78425
rect 54654 78362 54670 78426
rect 54734 78362 54750 78426
rect 54814 78425 54824 78426
rect 56383 78425 56627 78426
rect 54814 78362 56393 78425
rect 54240 78361 56393 78362
rect 56457 78361 56473 78425
rect 56537 78361 56553 78425
rect 56617 78361 56627 78425
rect 57269 78362 57270 78426
rect 57334 78362 57335 78426
rect 57269 78361 57335 78362
rect 54240 78206 54387 78361
rect 56383 78360 56627 78361
rect 53857 78204 54387 78206
rect 49828 78105 49894 78106
rect 49828 78041 49829 78105
rect 49893 78041 49894 78105
rect 49828 78040 49894 78041
rect 55228 78105 55294 78106
rect 55228 78041 55229 78105
rect 55293 78041 55303 78105
rect 55228 78040 55294 78041
rect 49020 77852 49086 77853
rect 49020 77788 49021 77852
rect 49085 77788 49086 77852
rect 49020 77787 49086 77788
rect 46557 77424 46623 77425
rect 46557 77360 46558 77424
rect 46622 77360 46623 77424
rect 46557 77359 46623 77360
rect 49021 76413 49085 77787
rect 49829 76736 49893 78040
rect 54420 77852 54486 77853
rect 54420 77788 54421 77852
rect 54485 77788 54495 77852
rect 54420 77787 54486 77788
rect 54421 77169 54485 77787
rect 55229 77425 55293 78040
rect 55228 77424 55294 77425
rect 55228 77360 55229 77424
rect 55293 77360 55294 77424
rect 57438 77422 57455 84828
rect 55228 77359 55294 77360
rect 54420 77168 54486 77169
rect 54420 77104 54421 77168
rect 54485 77104 54486 77168
rect 57432 77164 57455 77422
rect 57599 84147 57734 84828
rect 67270 84840 67646 84859
rect 57599 84146 57862 84147
rect 57599 84144 58380 84146
rect 57599 83908 57997 84144
rect 58233 83908 58380 84144
rect 67270 84135 67306 84840
rect 57599 83906 58380 83908
rect 65855 84133 67306 84135
rect 57599 81533 57734 83906
rect 65855 83897 66002 84133
rect 66238 83897 67306 84133
rect 65855 83895 67306 83897
rect 57599 81293 57851 81533
rect 57599 80772 57734 81293
rect 57599 80771 57762 80772
rect 57599 80769 58380 80771
rect 57599 80533 57997 80769
rect 58233 80533 58380 80769
rect 67270 80760 67306 83895
rect 57599 80531 58380 80533
rect 65854 80758 67306 80760
rect 57599 80530 57762 80531
rect 57599 77422 57734 80530
rect 65854 80522 66001 80758
rect 66237 80522 67306 80758
rect 65854 80520 67306 80522
rect 57599 77421 57765 77422
rect 57599 77394 58409 77421
rect 57599 77164 57997 77394
rect 57432 77158 57997 77164
rect 58233 77367 58409 77394
rect 67270 77385 67306 80520
rect 65854 77383 67306 77385
rect 58233 77189 58438 77367
rect 58233 77158 58409 77189
rect 57432 77126 58409 77158
rect 65854 77147 66001 77383
rect 66237 77147 67306 77383
rect 65854 77145 67306 77147
rect 54420 77103 54486 77104
rect 49828 76735 49894 76736
rect 49828 76671 49829 76735
rect 49893 76671 49894 76735
rect 49828 76670 49894 76671
rect 49020 76412 49086 76413
rect 49020 76348 49021 76412
rect 49085 76348 49086 76412
rect 49020 76347 49086 76348
rect 67270 76055 67306 77145
rect 67163 75877 67306 76055
rect 48084 75721 50387 75723
rect 48084 75485 50004 75721
rect 50240 75485 50387 75721
rect 48084 75483 50387 75485
rect 48084 75272 48324 75483
rect 48084 75265 48325 75272
rect 48084 75201 48250 75265
rect 48314 75201 48325 75265
rect 49371 75269 49437 75270
rect 49371 75205 49372 75269
rect 49436 75205 49437 75269
rect 49371 75204 49437 75205
rect 48084 75185 48325 75201
rect 48084 75121 48250 75185
rect 48314 75121 48325 75185
rect 48084 75105 48325 75121
rect 48084 75041 48250 75105
rect 48314 75041 48325 75105
rect 48084 75036 48325 75041
rect 48239 75035 48325 75036
rect 48219 74798 48317 74814
rect 48219 74734 48235 74798
rect 48299 74734 48317 74798
rect 48219 74718 48317 74734
rect 48219 74654 48235 74718
rect 48299 74654 48317 74718
rect 48219 74638 48317 74654
rect 48219 74574 48235 74638
rect 48299 74574 48317 74638
rect 48219 74558 48317 74574
rect 48219 74494 48235 74558
rect 48299 74494 48317 74558
rect 48219 74478 48317 74494
rect 48219 74414 48235 74478
rect 48299 74414 48317 74478
rect 48219 74399 48317 74414
rect 48613 74463 48679 74464
rect 48613 74399 48614 74463
rect 48678 74399 48679 74463
rect 48613 74398 48679 74399
rect 48614 74095 48678 74398
rect 48613 74094 48679 74095
rect 48613 74030 48614 74094
rect 48678 74030 48679 74094
rect 48613 74029 48679 74030
rect 46606 70655 46672 70656
rect 46606 70591 46607 70655
rect 46671 70591 46672 70655
rect 46606 70590 46672 70591
rect 46607 68641 46671 70590
rect 46189 68577 46671 68641
rect 44400 66420 44466 66421
rect 44400 66356 44401 66420
rect 44465 66356 44466 66420
rect 44400 66355 44466 66356
rect 44401 66350 44465 66355
rect 29932 66095 30023 66159
rect 30087 66095 30172 66159
rect 35618 66185 35684 66186
rect 35618 66121 35619 66185
rect 35683 66121 39414 66185
rect 35618 66120 35684 66121
rect 29932 66079 30172 66095
rect 29932 66015 30023 66079
rect 30087 66015 30172 66079
rect 29932 65999 30172 66015
rect 29932 65935 30023 65999
rect 30087 65935 30172 65999
rect 29932 65919 30172 65935
rect 29932 65855 30023 65919
rect 30087 65855 30172 65919
rect 29932 65839 30172 65855
rect 29932 65775 30023 65839
rect 30087 65775 30172 65839
rect 29932 65759 30172 65775
rect 29932 65695 30023 65759
rect 30087 65695 30172 65759
rect 29932 65679 30172 65695
rect 29932 65615 30023 65679
rect 30087 65615 30172 65679
rect 29932 65599 30172 65615
rect 29932 65535 30023 65599
rect 30087 65535 30172 65599
rect 29932 65519 30172 65535
rect 29932 65455 30023 65519
rect 30087 65455 30172 65519
rect 29932 65439 30172 65455
rect 29932 65375 30023 65439
rect 30087 65375 30172 65439
rect 29932 65359 30172 65375
rect 29932 65295 30023 65359
rect 30087 65295 30172 65359
rect 29932 65279 30172 65295
rect 29932 65215 30023 65279
rect 30087 65215 30172 65279
rect 29932 65199 30172 65215
rect 29932 65135 30023 65199
rect 30087 65135 30172 65199
rect 29932 65119 30172 65135
rect 29932 65055 30023 65119
rect 30087 65055 30172 65119
rect 29932 64633 30172 65055
rect 29932 64569 30028 64633
rect 30092 64569 30172 64633
rect 29932 64553 30172 64569
rect 29932 64489 30028 64553
rect 30092 64489 30172 64553
rect 29932 64473 30172 64489
rect 29932 64409 30028 64473
rect 30092 64409 30172 64473
rect 29932 64393 30172 64409
rect 29932 64329 30028 64393
rect 30092 64329 30172 64393
rect 29932 64313 30172 64329
rect 29932 64249 30028 64313
rect 30092 64249 30172 64313
rect 29932 64233 30172 64249
rect 29932 64169 30028 64233
rect 30092 64169 30172 64233
rect 29932 64153 30172 64169
rect 29932 64089 30028 64153
rect 30092 64089 30172 64153
rect 29932 64073 30172 64089
rect 29932 64009 30028 64073
rect 30092 64009 30172 64073
rect 29932 63993 30172 64009
rect 29932 63929 30028 63993
rect 30092 63972 30172 63993
rect 30092 63970 30395 63972
rect 29932 63913 30045 63929
rect 29932 63849 30028 63913
rect 29932 63833 30045 63849
rect 29932 63769 30028 63833
rect 29932 63753 30045 63769
rect 29932 63689 30028 63753
rect 30281 63734 30395 63970
rect 39350 63846 39414 66121
rect 39350 63782 39997 63846
rect 30092 63732 30395 63734
rect 30092 63689 30172 63732
rect 29932 63673 30172 63689
rect 29932 63609 30028 63673
rect 30092 63609 30172 63673
rect 29932 63593 30172 63609
rect 29932 63529 30028 63593
rect 30092 63529 30172 63593
rect 25281 63170 25347 63189
rect 25281 63106 25282 63170
rect 25346 63106 25347 63170
rect 25281 63090 25347 63106
rect 25281 63026 25282 63090
rect 25346 63045 25347 63090
rect 29932 63130 30172 63529
rect 29932 63066 30022 63130
rect 30086 63066 30172 63130
rect 29932 63050 30172 63066
rect 25346 63026 26149 63045
rect 25281 63010 26149 63026
rect 25281 62946 25282 63010
rect 25346 62981 26149 63010
rect 25346 62946 25347 62981
rect 25281 62930 25347 62946
rect 25281 62866 25282 62930
rect 25346 62866 25347 62930
rect 25281 62848 25347 62866
rect 25282 62631 25348 62636
rect 25282 62567 25283 62631
rect 25347 62567 25348 62631
rect 25282 62551 25348 62567
rect 21876 62518 22339 62520
rect 21876 62282 21989 62518
rect 22225 62437 22339 62518
rect 25282 62487 25283 62551
rect 25347 62487 25348 62551
rect 26085 62531 26149 62981
rect 29932 62986 30022 63050
rect 30086 62986 30172 63050
rect 29932 62970 30172 62986
rect 29932 62906 30022 62970
rect 30086 62906 30172 62970
rect 29932 62890 30172 62906
rect 29932 62826 30022 62890
rect 30086 62826 30172 62890
rect 29932 62810 30172 62826
rect 29932 62746 30022 62810
rect 30086 62746 30172 62810
rect 29932 62730 30172 62746
rect 29932 62666 30022 62730
rect 30086 62666 30172 62730
rect 29932 62650 30172 62666
rect 29932 62586 30022 62650
rect 30086 62586 30172 62650
rect 29932 62570 30172 62586
rect 25282 62471 25348 62487
rect 25282 62437 25283 62471
rect 22225 62407 25283 62437
rect 25347 62407 25348 62471
rect 22225 62391 25348 62407
rect 22225 62373 25283 62391
rect 22225 62282 22339 62373
rect 21876 62280 22339 62282
rect 25282 62327 25283 62373
rect 25347 62327 25348 62391
rect 25282 62311 25348 62327
rect 25282 62247 25283 62311
rect 25347 62247 25348 62311
rect 25888 62529 26351 62531
rect 25888 62293 26001 62529
rect 26237 62435 26351 62529
rect 29932 62506 30022 62570
rect 30086 62506 30172 62570
rect 29932 62490 30172 62506
rect 27479 62435 27945 62436
rect 26237 62371 27480 62435
rect 27544 62371 27560 62435
rect 27624 62371 27640 62435
rect 27704 62371 27720 62435
rect 27784 62371 27800 62435
rect 27864 62371 27880 62435
rect 27944 62371 27945 62435
rect 26237 62293 26351 62371
rect 27479 62370 27945 62371
rect 29932 62426 30022 62490
rect 30086 62426 30172 62490
rect 29932 62410 30172 62426
rect 25888 62291 26351 62293
rect 29932 62346 30022 62410
rect 30086 62346 30172 62410
rect 29932 62330 30172 62346
rect 25282 62231 25348 62247
rect 25282 62167 25283 62231
rect 25347 62167 25348 62231
rect 25282 62162 25348 62167
rect 29932 62266 30022 62330
rect 30086 62266 30172 62330
rect 25876 61431 26339 61433
rect 25876 61195 25989 61431
rect 26225 61345 26339 61431
rect 29932 61363 30172 62266
rect 38138 63524 38378 63711
rect 38138 63460 38217 63524
rect 38281 63460 38378 63524
rect 38138 63444 38378 63460
rect 38138 63380 38217 63444
rect 38281 63380 38378 63444
rect 38138 63364 38378 63380
rect 38138 63300 38217 63364
rect 38281 63300 38378 63364
rect 38138 63284 38378 63300
rect 38138 63220 38217 63284
rect 38281 63220 38378 63284
rect 38138 63204 38378 63220
rect 38138 63140 38217 63204
rect 38281 63140 38378 63204
rect 38138 63124 38378 63140
rect 38138 63060 38217 63124
rect 38281 63060 38378 63124
rect 38138 63044 38378 63060
rect 38138 62980 38217 63044
rect 38281 62980 38378 63044
rect 38138 62964 38378 62980
rect 38138 62900 38217 62964
rect 38281 62900 38378 62964
rect 38138 62884 38378 62900
rect 38138 62820 38217 62884
rect 38281 62820 38378 62884
rect 38138 62804 38378 62820
rect 45381 62813 45445 68564
rect 45380 62812 45446 62813
rect 43699 62805 43763 62806
rect 38138 62740 38217 62804
rect 38281 62740 38378 62804
rect 42196 62741 43763 62805
rect 45380 62748 45381 62812
rect 45445 62748 45446 62812
rect 45380 62747 45446 62748
rect 45381 62746 45445 62747
rect 38138 62724 38378 62740
rect 38138 62660 38217 62724
rect 38281 62660 38378 62724
rect 38138 62644 38378 62660
rect 38138 62580 38217 62644
rect 38281 62580 38378 62644
rect 38138 62564 38378 62580
rect 38138 62500 38217 62564
rect 38281 62500 38378 62564
rect 38138 62484 38378 62500
rect 38138 62420 38217 62484
rect 38281 62420 38378 62484
rect 38138 62404 38378 62420
rect 38138 62340 38217 62404
rect 38281 62340 38378 62404
rect 38138 62324 38378 62340
rect 38138 62260 38217 62324
rect 38281 62260 38378 62324
rect 38138 62244 38378 62260
rect 38138 62180 38217 62244
rect 38281 62180 38378 62244
rect 38138 62164 38378 62180
rect 38138 62100 38217 62164
rect 38281 62100 38378 62164
rect 38138 62084 38378 62100
rect 33902 61926 34365 62035
rect 38138 62020 38217 62084
rect 38281 62020 38378 62084
rect 38138 62004 38378 62020
rect 38138 61940 38217 62004
rect 38281 61940 38378 62004
rect 38138 61926 38378 61940
rect 33902 61924 38378 61926
rect 33902 61916 38217 61924
rect 33902 61680 34015 61916
rect 34251 61860 38217 61916
rect 38281 61860 38378 61924
rect 34251 61844 38378 61860
rect 34251 61780 38217 61844
rect 38281 61780 38378 61844
rect 41877 62303 42363 62322
rect 41877 61839 41888 62303
rect 42352 61839 42363 62303
rect 41877 61820 42363 61839
rect 34251 61764 38378 61780
rect 34251 61700 38217 61764
rect 38281 61700 38378 61764
rect 34251 61686 38378 61700
rect 34251 61680 34365 61686
rect 33902 61562 34365 61680
rect 38138 61684 38378 61686
rect 38138 61620 38217 61684
rect 38281 61620 38378 61684
rect 38138 61604 38378 61620
rect 27441 61345 27952 61346
rect 26225 61281 27464 61345
rect 27528 61281 27544 61345
rect 27608 61281 27624 61345
rect 27688 61281 27704 61345
rect 27768 61281 27784 61345
rect 27848 61281 27864 61345
rect 27928 61281 27952 61345
rect 26225 61195 26339 61281
rect 27441 61280 27952 61281
rect 29932 61299 30025 61363
rect 30089 61299 30172 61363
rect 29932 61283 30172 61299
rect 25876 61193 26339 61195
rect 29932 61219 30025 61283
rect 30089 61219 30172 61283
rect 29932 61203 30172 61219
rect 29932 61139 30025 61203
rect 30089 61139 30172 61203
rect 29932 61123 30172 61139
rect 29932 61059 30025 61123
rect 30089 61059 30172 61123
rect 29932 61043 30172 61059
rect 29932 60979 30025 61043
rect 30089 60979 30172 61043
rect 29932 60963 30172 60979
rect 29932 60899 30025 60963
rect 30089 60899 30172 60963
rect 29932 60883 30172 60899
rect 29932 60819 30025 60883
rect 30089 60819 30172 60883
rect 29932 60803 30172 60819
rect 29932 60739 30025 60803
rect 30089 60739 30172 60803
rect 29932 60723 30172 60739
rect 29932 60659 30025 60723
rect 30089 60659 30172 60723
rect 29932 60643 30172 60659
rect 29932 60579 30025 60643
rect 30089 60579 30172 60643
rect 29932 60563 30172 60579
rect 29932 60499 30025 60563
rect 30089 60499 30172 60563
rect 29932 60146 30172 60499
rect 29932 60082 30025 60146
rect 30089 60082 30172 60146
rect 29932 60066 30172 60082
rect 29932 60002 30025 60066
rect 30089 60002 30172 60066
rect 29932 59986 30172 60002
rect 29932 59922 30025 59986
rect 30089 59922 30172 59986
rect 38138 61540 38217 61604
rect 38281 61540 38378 61604
rect 38138 61524 38378 61540
rect 38138 61460 38217 61524
rect 38281 61460 38378 61524
rect 38138 61444 38378 61460
rect 38138 61380 38217 61444
rect 38281 61380 38378 61444
rect 38138 61364 38378 61380
rect 38138 61300 38217 61364
rect 38281 61300 38378 61364
rect 38138 61284 38378 61300
rect 38138 61220 38217 61284
rect 38281 61220 38378 61284
rect 38138 61204 38378 61220
rect 38138 61140 38217 61204
rect 38281 61140 38378 61204
rect 38138 61124 38378 61140
rect 38138 61060 38217 61124
rect 38281 61060 38378 61124
rect 38138 61044 38378 61060
rect 38138 60980 38217 61044
rect 38281 60980 38378 61044
rect 38138 60964 38378 60980
rect 38138 60900 38217 60964
rect 38281 60900 38378 60964
rect 38138 60884 38378 60900
rect 38138 60820 38217 60884
rect 38281 60820 38378 60884
rect 38138 60804 38378 60820
rect 38138 60740 38217 60804
rect 38281 60740 38378 60804
rect 38138 60724 38378 60740
rect 38138 60660 38217 60724
rect 38281 60660 38378 60724
rect 38138 60644 38378 60660
rect 38138 60580 38217 60644
rect 38281 60580 38378 60644
rect 38138 60564 38378 60580
rect 38138 60500 38217 60564
rect 38281 60500 38378 60564
rect 38138 60484 38378 60500
rect 38138 60420 38217 60484
rect 38281 60420 38378 60484
rect 38138 60404 38378 60420
rect 38138 60340 38217 60404
rect 38281 60340 38378 60404
rect 38138 60324 38378 60340
rect 38138 60260 38217 60324
rect 38281 60260 38378 60324
rect 38138 60244 38378 60260
rect 38138 60180 38217 60244
rect 38281 60180 38378 60244
rect 38138 59979 38378 60180
rect 39351 60351 40088 60415
rect 29932 59906 30172 59922
rect 29932 59842 30025 59906
rect 30089 59903 30172 59906
rect 30089 59901 30395 59903
rect 29932 59826 30045 59842
rect 29932 59762 30025 59826
rect 29932 59746 30045 59762
rect 29932 59682 30025 59746
rect 29932 59666 30045 59682
rect 29932 59602 30025 59666
rect 30281 59665 30395 59901
rect 30089 59663 30395 59665
rect 30089 59602 30172 59663
rect 29932 59586 30172 59602
rect 29932 59522 30025 59586
rect 30089 59522 30172 59586
rect 29932 59506 30172 59522
rect 29932 59442 30025 59506
rect 30089 59442 30172 59506
rect 29932 59426 30172 59442
rect 29932 59362 30025 59426
rect 30089 59362 30172 59426
rect 29932 59346 30172 59362
rect 29932 59282 30025 59346
rect 30089 59282 30172 59346
rect 29932 59266 30172 59282
rect 29932 59202 30025 59266
rect 30089 59202 30172 59266
rect 29932 59186 30172 59202
rect 29932 59122 30025 59186
rect 30089 59122 30172 59186
rect 29932 59106 30172 59122
rect 29932 59042 30025 59106
rect 30089 59042 30172 59106
rect 29932 58708 30172 59042
rect 29932 58644 30022 58708
rect 30086 58644 30172 58708
rect 29932 58628 30172 58644
rect 29932 58564 30022 58628
rect 30086 58564 30172 58628
rect 29932 58548 30172 58564
rect 29932 58484 30022 58548
rect 30086 58484 30172 58548
rect 29932 58468 30172 58484
rect 29932 58404 30022 58468
rect 30086 58404 30172 58468
rect 29932 58388 30172 58404
rect 29932 58324 30022 58388
rect 30086 58324 30172 58388
rect 29932 58308 30172 58324
rect 29932 58244 30022 58308
rect 30086 58244 30172 58308
rect 29932 58228 30172 58244
rect 29932 58164 30022 58228
rect 30086 58164 30172 58228
rect 29932 58148 30172 58164
rect 29932 58084 30022 58148
rect 30086 58084 30172 58148
rect 29932 58068 30172 58084
rect 29932 58004 30022 58068
rect 30086 58004 30172 58068
rect 29932 57988 30172 58004
rect 29932 57924 30022 57988
rect 30086 57924 30172 57988
rect 29932 57908 30172 57924
rect 29932 57844 30022 57908
rect 30086 57844 30172 57908
rect 29932 57828 30172 57844
rect 29932 57764 30022 57828
rect 30086 57764 30172 57828
rect 29932 57748 30172 57764
rect 29932 57684 30022 57748
rect 30086 57684 30172 57748
rect 29932 57668 30172 57684
rect 29932 57604 30022 57668
rect 30086 57604 30172 57668
rect 29932 57588 30172 57604
rect 29932 57524 30022 57588
rect 30086 57524 30172 57588
rect 29932 56886 30172 57524
rect 35575 57573 35641 57574
rect 39351 57573 39415 60351
rect 35575 57509 35576 57573
rect 35640 57509 39415 57573
rect 35575 57508 35641 57509
rect 41955 57202 42019 59368
rect 43699 58699 43763 62741
rect 46189 62470 46253 68577
rect 47885 67083 47951 67084
rect 47885 67019 47886 67083
rect 47950 67019 47951 67083
rect 47885 67018 47951 67019
rect 47024 66420 47090 66421
rect 47024 66356 47025 66420
rect 47089 66356 47090 66420
rect 47024 66355 47090 66356
rect 46188 62469 46254 62470
rect 46188 62405 46189 62469
rect 46253 62405 46254 62469
rect 46188 62404 46254 62405
rect 46189 62398 46253 62404
rect 47025 59374 47089 66355
rect 47886 59964 47950 67018
rect 48614 61394 48678 74029
rect 49372 73447 49436 75204
rect 51122 75143 51399 75146
rect 51122 75121 57233 75143
rect 51122 75079 54010 75121
rect 54246 75079 57233 75121
rect 51122 75068 53753 75079
rect 51122 74924 51434 75068
rect 53178 74935 53753 75068
rect 54537 75069 57233 75079
rect 54537 74935 55452 75069
rect 53178 74924 54010 74935
rect 51122 74885 54010 74924
rect 54246 74925 55452 74935
rect 56316 74925 57233 75069
rect 54246 74885 57233 74925
rect 51122 74867 57233 74885
rect 51122 74742 51399 74867
rect 49371 73446 49437 73447
rect 49371 73382 49372 73446
rect 49436 73382 49437 73446
rect 49371 73381 49437 73382
rect 49372 61922 49436 73381
rect 51122 71798 51182 74742
rect 51326 72813 51399 74742
rect 56956 74757 57233 74867
rect 56956 72813 57043 74757
rect 51326 72793 57043 72813
rect 51326 72557 54004 72793
rect 54240 72557 57043 72793
rect 51326 72536 57043 72557
rect 51326 71798 51399 72536
rect 51122 71710 51399 71798
rect 56956 71813 57043 72536
rect 57187 71813 57233 74757
rect 57694 74019 58392 74039
rect 57694 73783 57997 74019
rect 58233 73783 58392 74019
rect 67270 74010 67306 75877
rect 57694 73744 58392 73783
rect 65854 74008 67306 74010
rect 65854 73772 66001 74008
rect 66237 73772 67306 74008
rect 65854 73770 67306 73772
rect 56956 71737 57233 71813
rect 67270 71656 67306 73770
rect 67610 71656 67646 84840
rect 73811 84750 90426 84789
rect 73811 84686 74525 84750
rect 74589 84686 75613 84750
rect 75677 84686 76701 84750
rect 76765 84686 77789 84750
rect 77853 84686 78877 84750
rect 78941 84686 79965 84750
rect 80029 84686 81053 84750
rect 81117 84686 82141 84750
rect 82205 84686 83229 84750
rect 83293 84686 84317 84750
rect 84381 84686 85405 84750
rect 85469 84686 86493 84750
rect 86557 84686 87581 84750
rect 87645 84686 88669 84750
rect 88733 84686 90426 84750
rect 73811 84670 90426 84686
rect 73811 84606 74525 84670
rect 74589 84606 75613 84670
rect 75677 84606 76701 84670
rect 76765 84606 77789 84670
rect 77853 84606 78877 84670
rect 78941 84606 79965 84670
rect 80029 84606 81053 84670
rect 81117 84606 82141 84670
rect 82205 84606 83229 84670
rect 83293 84606 84317 84670
rect 84381 84606 85405 84670
rect 85469 84606 86493 84670
rect 86557 84606 87581 84670
rect 87645 84606 88669 84670
rect 88733 84606 90426 84670
rect 73811 84601 90426 84606
rect 73811 84595 85995 84601
rect 73811 84590 78001 84595
rect 73811 84526 74525 84590
rect 74589 84526 75613 84590
rect 75677 84526 76701 84590
rect 76765 84526 77789 84590
rect 77853 84526 78001 84590
rect 73811 84510 78001 84526
rect 73811 84446 74525 84510
rect 74589 84446 75613 84510
rect 75677 84446 76701 84510
rect 76765 84446 77789 84510
rect 77853 84446 78001 84510
rect 73811 84430 78001 84446
rect 73811 84366 74525 84430
rect 74589 84366 75613 84430
rect 75677 84366 76701 84430
rect 76765 84366 77789 84430
rect 77853 84366 78001 84430
rect 73811 84359 78001 84366
rect 78237 84590 85995 84595
rect 78237 84526 78877 84590
rect 78941 84526 79965 84590
rect 80029 84526 81053 84590
rect 81117 84526 82141 84590
rect 82205 84526 83229 84590
rect 83293 84526 84317 84590
rect 84381 84526 85405 84590
rect 85469 84526 85995 84590
rect 78237 84510 85995 84526
rect 78237 84446 78877 84510
rect 78941 84446 79965 84510
rect 80029 84446 81053 84510
rect 81117 84446 82141 84510
rect 82205 84446 83229 84510
rect 83293 84446 84317 84510
rect 84381 84446 85405 84510
rect 85469 84446 85995 84510
rect 78237 84430 85995 84446
rect 78237 84366 78877 84430
rect 78941 84366 79965 84430
rect 80029 84366 81053 84430
rect 81117 84366 82141 84430
rect 82205 84366 83229 84430
rect 83293 84366 84317 84430
rect 84381 84366 85405 84430
rect 85469 84366 85995 84430
rect 78237 84365 85995 84366
rect 86231 84590 90426 84601
rect 86231 84526 86493 84590
rect 86557 84526 87581 84590
rect 87645 84526 88669 84590
rect 88733 84526 90426 84590
rect 86231 84510 90426 84526
rect 86231 84446 86493 84510
rect 86557 84446 87581 84510
rect 87645 84446 88669 84510
rect 88733 84446 90426 84510
rect 86231 84430 90426 84446
rect 86231 84366 86493 84430
rect 86557 84366 87581 84430
rect 87645 84366 88669 84430
rect 88733 84366 90426 84430
rect 86231 84365 90426 84366
rect 78237 84359 90426 84365
rect 73811 84350 90426 84359
rect 73811 84286 74525 84350
rect 74589 84286 75613 84350
rect 75677 84286 76701 84350
rect 76765 84286 77789 84350
rect 77853 84286 78877 84350
rect 78941 84286 79965 84350
rect 80029 84286 81053 84350
rect 81117 84286 82141 84350
rect 82205 84286 83229 84350
rect 83293 84286 84317 84350
rect 84381 84286 85405 84350
rect 85469 84286 86493 84350
rect 86557 84286 87581 84350
rect 87645 84286 88669 84350
rect 88733 84286 90426 84350
rect 73811 84270 90426 84286
rect 73811 84206 74525 84270
rect 74589 84206 75613 84270
rect 75677 84206 76701 84270
rect 76765 84206 77789 84270
rect 77853 84206 78877 84270
rect 78941 84206 79965 84270
rect 80029 84206 81053 84270
rect 81117 84206 82141 84270
rect 82205 84206 83229 84270
rect 83293 84206 84317 84270
rect 84381 84206 85405 84270
rect 85469 84206 86493 84270
rect 86557 84206 87581 84270
rect 87645 84206 88669 84270
rect 88733 84206 90426 84270
rect 73811 84169 90426 84206
rect 73809 82747 90321 82789
rect 73809 82683 75070 82747
rect 75134 82683 76158 82747
rect 76222 82683 77246 82747
rect 77310 82683 78334 82747
rect 78398 82683 79422 82747
rect 79486 82683 80510 82747
rect 80574 82683 81598 82747
rect 81662 82683 82686 82747
rect 82750 82683 83774 82747
rect 83838 82683 84862 82747
rect 84926 82683 85950 82747
rect 86014 82683 87038 82747
rect 87102 82683 88126 82747
rect 88190 82739 90321 82747
rect 88190 82683 90384 82739
rect 73809 82667 90384 82683
rect 73809 82604 75070 82667
rect 73809 82368 74004 82604
rect 74240 82603 75070 82604
rect 75134 82603 76158 82667
rect 76222 82603 77246 82667
rect 77310 82603 78334 82667
rect 78398 82603 79422 82667
rect 79486 82603 80510 82667
rect 80574 82603 81598 82667
rect 81662 82603 82686 82667
rect 82750 82603 83774 82667
rect 83838 82603 84862 82667
rect 84926 82603 85950 82667
rect 86014 82603 87038 82667
rect 87102 82603 88126 82667
rect 88190 82603 90384 82667
rect 74240 82597 90384 82603
rect 74240 82587 82000 82597
rect 74240 82523 75070 82587
rect 75134 82523 76158 82587
rect 76222 82523 77246 82587
rect 77310 82523 78334 82587
rect 78398 82523 79422 82587
rect 79486 82523 80510 82587
rect 80574 82523 81598 82587
rect 81662 82523 82000 82587
rect 74240 82507 82000 82523
rect 74240 82443 75070 82507
rect 75134 82443 76158 82507
rect 76222 82443 77246 82507
rect 77310 82443 78334 82507
rect 78398 82443 79422 82507
rect 79486 82443 80510 82507
rect 80574 82443 81598 82507
rect 81662 82443 82000 82507
rect 74240 82427 82000 82443
rect 74240 82368 75070 82427
rect 73809 82363 75070 82368
rect 75134 82363 76158 82427
rect 76222 82363 77246 82427
rect 77310 82363 78334 82427
rect 78398 82363 79422 82427
rect 79486 82363 80510 82427
rect 80574 82363 81598 82427
rect 81662 82363 82000 82427
rect 73809 82361 82000 82363
rect 82236 82593 90384 82597
rect 82236 82587 90003 82593
rect 82236 82523 82686 82587
rect 82750 82523 83774 82587
rect 83838 82523 84862 82587
rect 84926 82523 85950 82587
rect 86014 82523 87038 82587
rect 87102 82523 88126 82587
rect 88190 82523 90003 82587
rect 82236 82507 90003 82523
rect 82236 82443 82686 82507
rect 82750 82443 83774 82507
rect 83838 82443 84862 82507
rect 84926 82443 85950 82507
rect 86014 82443 87038 82507
rect 87102 82443 88126 82507
rect 88190 82443 90003 82507
rect 82236 82427 90003 82443
rect 82236 82363 82686 82427
rect 82750 82363 83774 82427
rect 83838 82363 84862 82427
rect 84926 82363 85950 82427
rect 86014 82363 87038 82427
rect 87102 82363 88126 82427
rect 88190 82363 90003 82427
rect 82236 82361 90003 82363
rect 73809 82357 90003 82361
rect 90239 82357 90384 82593
rect 73809 82347 90384 82357
rect 73809 82283 75070 82347
rect 75134 82283 76158 82347
rect 76222 82283 77246 82347
rect 77310 82283 78334 82347
rect 78398 82283 79422 82347
rect 79486 82283 80510 82347
rect 80574 82283 81598 82347
rect 81662 82283 82686 82347
rect 82750 82283 83774 82347
rect 83838 82283 84862 82347
rect 84926 82283 85950 82347
rect 86014 82283 87038 82347
rect 87102 82283 88126 82347
rect 88190 82283 90384 82347
rect 73809 82267 90384 82283
rect 73809 82203 75070 82267
rect 75134 82203 76158 82267
rect 76222 82203 77246 82267
rect 77310 82203 78334 82267
rect 78398 82203 79422 82267
rect 79486 82203 80510 82267
rect 80574 82203 81598 82267
rect 81662 82203 82686 82267
rect 82750 82203 83774 82267
rect 83838 82203 84862 82267
rect 84926 82203 85950 82267
rect 86014 82203 87038 82267
rect 87102 82203 88126 82267
rect 88190 82211 90384 82267
rect 88190 82203 90321 82211
rect 73809 82169 90321 82203
rect 73811 80750 90426 80789
rect 73811 80686 74525 80750
rect 74589 80686 75613 80750
rect 75677 80686 76701 80750
rect 76765 80686 77789 80750
rect 77853 80686 78877 80750
rect 78941 80686 79965 80750
rect 80029 80686 81053 80750
rect 81117 80686 82141 80750
rect 82205 80686 83229 80750
rect 83293 80686 84317 80750
rect 84381 80686 85405 80750
rect 85469 80686 86493 80750
rect 86557 80686 87581 80750
rect 87645 80686 88669 80750
rect 88733 80686 90426 80750
rect 73811 80670 90426 80686
rect 73811 80606 74525 80670
rect 74589 80606 75613 80670
rect 75677 80606 76701 80670
rect 76765 80606 77789 80670
rect 77853 80606 78877 80670
rect 78941 80606 79965 80670
rect 80029 80606 81053 80670
rect 81117 80606 82141 80670
rect 82205 80606 83229 80670
rect 83293 80606 84317 80670
rect 84381 80606 85405 80670
rect 85469 80606 86493 80670
rect 86557 80606 87581 80670
rect 87645 80606 88669 80670
rect 88733 80606 90426 80670
rect 73811 80601 90426 80606
rect 73811 80595 85995 80601
rect 73811 80590 78001 80595
rect 73811 80526 74525 80590
rect 74589 80526 75613 80590
rect 75677 80526 76701 80590
rect 76765 80526 77789 80590
rect 77853 80526 78001 80590
rect 73811 80510 78001 80526
rect 73811 80446 74525 80510
rect 74589 80446 75613 80510
rect 75677 80446 76701 80510
rect 76765 80446 77789 80510
rect 77853 80446 78001 80510
rect 73811 80430 78001 80446
rect 73811 80366 74525 80430
rect 74589 80366 75613 80430
rect 75677 80366 76701 80430
rect 76765 80366 77789 80430
rect 77853 80366 78001 80430
rect 73811 80359 78001 80366
rect 78237 80590 85995 80595
rect 78237 80526 78877 80590
rect 78941 80526 79965 80590
rect 80029 80526 81053 80590
rect 81117 80526 82141 80590
rect 82205 80526 83229 80590
rect 83293 80526 84317 80590
rect 84381 80526 85405 80590
rect 85469 80526 85995 80590
rect 78237 80510 85995 80526
rect 78237 80446 78877 80510
rect 78941 80446 79965 80510
rect 80029 80446 81053 80510
rect 81117 80446 82141 80510
rect 82205 80446 83229 80510
rect 83293 80446 84317 80510
rect 84381 80446 85405 80510
rect 85469 80446 85995 80510
rect 78237 80430 85995 80446
rect 78237 80366 78877 80430
rect 78941 80366 79965 80430
rect 80029 80366 81053 80430
rect 81117 80366 82141 80430
rect 82205 80366 83229 80430
rect 83293 80366 84317 80430
rect 84381 80366 85405 80430
rect 85469 80366 85995 80430
rect 78237 80365 85995 80366
rect 86231 80590 90426 80601
rect 86231 80526 86493 80590
rect 86557 80526 87581 80590
rect 87645 80526 88669 80590
rect 88733 80526 90426 80590
rect 86231 80510 90426 80526
rect 86231 80446 86493 80510
rect 86557 80446 87581 80510
rect 87645 80446 88669 80510
rect 88733 80446 90426 80510
rect 86231 80430 90426 80446
rect 86231 80366 86493 80430
rect 86557 80366 87581 80430
rect 87645 80366 88669 80430
rect 88733 80366 90426 80430
rect 86231 80365 90426 80366
rect 78237 80359 90426 80365
rect 73811 80350 90426 80359
rect 73811 80286 74525 80350
rect 74589 80286 75613 80350
rect 75677 80286 76701 80350
rect 76765 80286 77789 80350
rect 77853 80286 78877 80350
rect 78941 80286 79965 80350
rect 80029 80286 81053 80350
rect 81117 80286 82141 80350
rect 82205 80286 83229 80350
rect 83293 80286 84317 80350
rect 84381 80286 85405 80350
rect 85469 80286 86493 80350
rect 86557 80286 87581 80350
rect 87645 80286 88669 80350
rect 88733 80286 90426 80350
rect 73811 80270 90426 80286
rect 73811 80206 74525 80270
rect 74589 80206 75613 80270
rect 75677 80206 76701 80270
rect 76765 80206 77789 80270
rect 77853 80206 78877 80270
rect 78941 80206 79965 80270
rect 80029 80206 81053 80270
rect 81117 80206 82141 80270
rect 82205 80206 83229 80270
rect 83293 80206 84317 80270
rect 84381 80206 85405 80270
rect 85469 80206 86493 80270
rect 86557 80206 87581 80270
rect 87645 80206 88669 80270
rect 88733 80206 90426 80270
rect 73811 80169 90426 80206
rect 73809 78747 90321 78789
rect 73809 78683 75070 78747
rect 75134 78683 76158 78747
rect 76222 78683 77246 78747
rect 77310 78683 78334 78747
rect 78398 78683 79422 78747
rect 79486 78683 80510 78747
rect 80574 78683 81598 78747
rect 81662 78683 82686 78747
rect 82750 78683 83774 78747
rect 83838 78683 84862 78747
rect 84926 78683 85950 78747
rect 86014 78683 87038 78747
rect 87102 78683 88126 78747
rect 88190 78739 90321 78747
rect 88190 78683 90384 78739
rect 73809 78667 90384 78683
rect 73809 78604 75070 78667
rect 73809 78368 74004 78604
rect 74240 78603 75070 78604
rect 75134 78603 76158 78667
rect 76222 78603 77246 78667
rect 77310 78603 78334 78667
rect 78398 78603 79422 78667
rect 79486 78603 80510 78667
rect 80574 78603 81598 78667
rect 81662 78603 82686 78667
rect 82750 78603 83774 78667
rect 83838 78603 84862 78667
rect 84926 78603 85950 78667
rect 86014 78603 87038 78667
rect 87102 78603 88126 78667
rect 88190 78603 90384 78667
rect 74240 78597 90384 78603
rect 74240 78587 82000 78597
rect 74240 78523 75070 78587
rect 75134 78523 76158 78587
rect 76222 78523 77246 78587
rect 77310 78523 78334 78587
rect 78398 78523 79422 78587
rect 79486 78523 80510 78587
rect 80574 78523 81598 78587
rect 81662 78523 82000 78587
rect 74240 78507 82000 78523
rect 74240 78443 75070 78507
rect 75134 78443 76158 78507
rect 76222 78443 77246 78507
rect 77310 78443 78334 78507
rect 78398 78443 79422 78507
rect 79486 78443 80510 78507
rect 80574 78443 81598 78507
rect 81662 78443 82000 78507
rect 74240 78427 82000 78443
rect 74240 78368 75070 78427
rect 73809 78363 75070 78368
rect 75134 78363 76158 78427
rect 76222 78363 77246 78427
rect 77310 78363 78334 78427
rect 78398 78363 79422 78427
rect 79486 78363 80510 78427
rect 80574 78363 81598 78427
rect 81662 78363 82000 78427
rect 73809 78361 82000 78363
rect 82236 78593 90384 78597
rect 82236 78587 90003 78593
rect 82236 78523 82686 78587
rect 82750 78523 83774 78587
rect 83838 78523 84862 78587
rect 84926 78523 85950 78587
rect 86014 78523 87038 78587
rect 87102 78523 88126 78587
rect 88190 78523 90003 78587
rect 82236 78507 90003 78523
rect 82236 78443 82686 78507
rect 82750 78443 83774 78507
rect 83838 78443 84862 78507
rect 84926 78443 85950 78507
rect 86014 78443 87038 78507
rect 87102 78443 88126 78507
rect 88190 78443 90003 78507
rect 82236 78427 90003 78443
rect 82236 78363 82686 78427
rect 82750 78363 83774 78427
rect 83838 78363 84862 78427
rect 84926 78363 85950 78427
rect 86014 78363 87038 78427
rect 87102 78363 88126 78427
rect 88190 78363 90003 78427
rect 82236 78361 90003 78363
rect 73809 78357 90003 78361
rect 90239 78357 90384 78593
rect 73809 78347 90384 78357
rect 73809 78283 75070 78347
rect 75134 78283 76158 78347
rect 76222 78283 77246 78347
rect 77310 78283 78334 78347
rect 78398 78283 79422 78347
rect 79486 78283 80510 78347
rect 80574 78283 81598 78347
rect 81662 78283 82686 78347
rect 82750 78283 83774 78347
rect 83838 78283 84862 78347
rect 84926 78283 85950 78347
rect 86014 78283 87038 78347
rect 87102 78283 88126 78347
rect 88190 78283 90384 78347
rect 73809 78267 90384 78283
rect 73809 78203 75070 78267
rect 75134 78203 76158 78267
rect 76222 78203 77246 78267
rect 77310 78203 78334 78267
rect 78398 78203 79422 78267
rect 79486 78203 80510 78267
rect 80574 78203 81598 78267
rect 81662 78203 82686 78267
rect 82750 78203 83774 78267
rect 83838 78203 84862 78267
rect 84926 78203 85950 78267
rect 86014 78203 87038 78267
rect 87102 78203 88126 78267
rect 88190 78211 90384 78267
rect 88190 78203 90321 78211
rect 73809 78169 90321 78203
rect 73811 76750 90426 76789
rect 73811 76686 74525 76750
rect 74589 76686 75613 76750
rect 75677 76686 76701 76750
rect 76765 76686 77789 76750
rect 77853 76686 78877 76750
rect 78941 76686 79965 76750
rect 80029 76686 81053 76750
rect 81117 76686 82141 76750
rect 82205 76686 83229 76750
rect 83293 76686 84317 76750
rect 84381 76686 85405 76750
rect 85469 76686 86493 76750
rect 86557 76686 87581 76750
rect 87645 76686 88669 76750
rect 88733 76686 90426 76750
rect 73811 76670 90426 76686
rect 73811 76606 74525 76670
rect 74589 76606 75613 76670
rect 75677 76606 76701 76670
rect 76765 76606 77789 76670
rect 77853 76606 78877 76670
rect 78941 76606 79965 76670
rect 80029 76606 81053 76670
rect 81117 76606 82141 76670
rect 82205 76606 83229 76670
rect 83293 76606 84317 76670
rect 84381 76606 85405 76670
rect 85469 76606 86493 76670
rect 86557 76606 87581 76670
rect 87645 76606 88669 76670
rect 88733 76606 90426 76670
rect 73811 76601 90426 76606
rect 73811 76595 85995 76601
rect 73811 76590 78001 76595
rect 73811 76526 74525 76590
rect 74589 76526 75613 76590
rect 75677 76526 76701 76590
rect 76765 76526 77789 76590
rect 77853 76526 78001 76590
rect 73811 76510 78001 76526
rect 73811 76446 74525 76510
rect 74589 76446 75613 76510
rect 75677 76446 76701 76510
rect 76765 76446 77789 76510
rect 77853 76446 78001 76510
rect 73811 76430 78001 76446
rect 73811 76366 74525 76430
rect 74589 76366 75613 76430
rect 75677 76366 76701 76430
rect 76765 76366 77789 76430
rect 77853 76366 78001 76430
rect 73811 76359 78001 76366
rect 78237 76590 85995 76595
rect 78237 76526 78877 76590
rect 78941 76526 79965 76590
rect 80029 76526 81053 76590
rect 81117 76526 82141 76590
rect 82205 76526 83229 76590
rect 83293 76526 84317 76590
rect 84381 76526 85405 76590
rect 85469 76526 85995 76590
rect 78237 76510 85995 76526
rect 78237 76446 78877 76510
rect 78941 76446 79965 76510
rect 80029 76446 81053 76510
rect 81117 76446 82141 76510
rect 82205 76446 83229 76510
rect 83293 76446 84317 76510
rect 84381 76446 85405 76510
rect 85469 76446 85995 76510
rect 78237 76430 85995 76446
rect 78237 76366 78877 76430
rect 78941 76366 79965 76430
rect 80029 76366 81053 76430
rect 81117 76366 82141 76430
rect 82205 76366 83229 76430
rect 83293 76366 84317 76430
rect 84381 76366 85405 76430
rect 85469 76366 85995 76430
rect 78237 76365 85995 76366
rect 86231 76590 90426 76601
rect 86231 76526 86493 76590
rect 86557 76526 87581 76590
rect 87645 76526 88669 76590
rect 88733 76526 90426 76590
rect 86231 76510 90426 76526
rect 86231 76446 86493 76510
rect 86557 76446 87581 76510
rect 87645 76446 88669 76510
rect 88733 76446 90426 76510
rect 86231 76430 90426 76446
rect 86231 76366 86493 76430
rect 86557 76366 87581 76430
rect 87645 76366 88669 76430
rect 88733 76366 90426 76430
rect 86231 76365 90426 76366
rect 78237 76359 90426 76365
rect 73811 76350 90426 76359
rect 73811 76286 74525 76350
rect 74589 76286 75613 76350
rect 75677 76286 76701 76350
rect 76765 76286 77789 76350
rect 77853 76286 78877 76350
rect 78941 76286 79965 76350
rect 80029 76286 81053 76350
rect 81117 76286 82141 76350
rect 82205 76286 83229 76350
rect 83293 76286 84317 76350
rect 84381 76286 85405 76350
rect 85469 76286 86493 76350
rect 86557 76286 87581 76350
rect 87645 76286 88669 76350
rect 88733 76286 90426 76350
rect 73811 76270 90426 76286
rect 73811 76206 74525 76270
rect 74589 76206 75613 76270
rect 75677 76206 76701 76270
rect 76765 76206 77789 76270
rect 77853 76206 78877 76270
rect 78941 76206 79965 76270
rect 80029 76206 81053 76270
rect 81117 76206 82141 76270
rect 82205 76206 83229 76270
rect 83293 76206 84317 76270
rect 84381 76206 85405 76270
rect 85469 76206 86493 76270
rect 86557 76206 87581 76270
rect 87645 76206 88669 76270
rect 88733 76206 90426 76270
rect 73811 76169 90426 76206
rect 73809 74747 90321 74789
rect 73809 74683 75070 74747
rect 75134 74683 77246 74747
rect 77310 74683 78334 74747
rect 78398 74683 80510 74747
rect 80574 74683 81598 74747
rect 81662 74683 82686 74747
rect 82750 74683 84862 74747
rect 84926 74683 85950 74747
rect 86014 74683 88126 74747
rect 88190 74739 90321 74747
rect 88190 74683 90384 74739
rect 73809 74667 90384 74683
rect 73809 74604 75070 74667
rect 73809 74368 74004 74604
rect 74240 74603 75070 74604
rect 75134 74603 77246 74667
rect 77310 74603 78334 74667
rect 78398 74603 80510 74667
rect 80574 74603 81598 74667
rect 81662 74603 82686 74667
rect 82750 74603 84862 74667
rect 84926 74603 85950 74667
rect 86014 74603 88126 74667
rect 88190 74603 90384 74667
rect 74240 74597 90384 74603
rect 74240 74587 82000 74597
rect 74240 74523 75070 74587
rect 75134 74523 77246 74587
rect 77310 74523 78334 74587
rect 78398 74523 80510 74587
rect 80574 74523 81598 74587
rect 81662 74523 82000 74587
rect 74240 74507 82000 74523
rect 74240 74443 75070 74507
rect 75134 74443 77246 74507
rect 77310 74443 78334 74507
rect 78398 74443 80510 74507
rect 80574 74443 81598 74507
rect 81662 74443 82000 74507
rect 74240 74427 82000 74443
rect 74240 74368 75070 74427
rect 73809 74363 75070 74368
rect 75134 74363 77246 74427
rect 77310 74363 78334 74427
rect 78398 74363 80510 74427
rect 80574 74363 81598 74427
rect 81662 74363 82000 74427
rect 73809 74361 82000 74363
rect 82236 74593 90384 74597
rect 82236 74587 90003 74593
rect 82236 74523 82686 74587
rect 82750 74523 84862 74587
rect 84926 74523 85950 74587
rect 86014 74523 88126 74587
rect 88190 74523 90003 74587
rect 82236 74507 90003 74523
rect 82236 74443 82686 74507
rect 82750 74443 84862 74507
rect 84926 74443 85950 74507
rect 86014 74443 88126 74507
rect 88190 74443 90003 74507
rect 82236 74427 90003 74443
rect 82236 74363 82686 74427
rect 82750 74363 84862 74427
rect 84926 74363 85950 74427
rect 86014 74363 88126 74427
rect 88190 74363 90003 74427
rect 82236 74361 90003 74363
rect 73809 74357 90003 74361
rect 90239 74357 90384 74593
rect 73809 74347 90384 74357
rect 73809 74283 75070 74347
rect 75134 74283 77246 74347
rect 77310 74283 78334 74347
rect 78398 74283 80510 74347
rect 80574 74283 81598 74347
rect 81662 74283 82686 74347
rect 82750 74283 84862 74347
rect 84926 74283 85950 74347
rect 86014 74283 88126 74347
rect 88190 74283 90384 74347
rect 73809 74267 90384 74283
rect 73809 74203 75070 74267
rect 75134 74203 77246 74267
rect 77310 74203 78334 74267
rect 78398 74203 80510 74267
rect 80574 74203 81598 74267
rect 81662 74203 82686 74267
rect 82750 74203 84862 74267
rect 84926 74203 85950 74267
rect 86014 74203 88126 74267
rect 88190 74211 90384 74267
rect 88190 74203 90321 74211
rect 73809 74169 90321 74203
rect 73811 72750 90426 72789
rect 73811 72686 74525 72750
rect 74589 72686 75613 72750
rect 75677 72686 76701 72750
rect 76765 72686 77789 72750
rect 77853 72686 78877 72750
rect 78941 72686 79965 72750
rect 80029 72686 81053 72750
rect 81117 72686 86493 72750
rect 86557 72686 87581 72750
rect 87645 72686 88669 72750
rect 88733 72686 90426 72750
rect 73811 72670 90426 72686
rect 73811 72606 74525 72670
rect 74589 72606 75613 72670
rect 75677 72606 76701 72670
rect 76765 72606 77789 72670
rect 77853 72606 78877 72670
rect 78941 72606 79965 72670
rect 80029 72606 81053 72670
rect 81117 72606 86493 72670
rect 86557 72606 87581 72670
rect 87645 72606 88669 72670
rect 88733 72606 90426 72670
rect 73811 72601 90426 72606
rect 73811 72595 85995 72601
rect 73811 72590 78001 72595
rect 73811 72526 74525 72590
rect 74589 72526 75613 72590
rect 75677 72526 76701 72590
rect 76765 72526 77789 72590
rect 77853 72526 78001 72590
rect 73811 72510 78001 72526
rect 73811 72446 74525 72510
rect 74589 72446 75613 72510
rect 75677 72446 76701 72510
rect 76765 72446 77789 72510
rect 77853 72446 78001 72510
rect 73811 72430 78001 72446
rect 73811 72366 74525 72430
rect 74589 72366 75613 72430
rect 75677 72366 76701 72430
rect 76765 72366 77789 72430
rect 77853 72366 78001 72430
rect 73811 72359 78001 72366
rect 78237 72590 85995 72595
rect 78237 72526 78877 72590
rect 78941 72526 79965 72590
rect 80029 72526 81053 72590
rect 81117 72526 85995 72590
rect 78237 72510 85995 72526
rect 78237 72446 78877 72510
rect 78941 72446 79965 72510
rect 80029 72446 81053 72510
rect 81117 72446 85995 72510
rect 78237 72430 85995 72446
rect 78237 72366 78877 72430
rect 78941 72366 79965 72430
rect 80029 72366 81053 72430
rect 81117 72366 85995 72430
rect 78237 72365 85995 72366
rect 86231 72590 90426 72601
rect 86231 72526 86493 72590
rect 86557 72526 87581 72590
rect 87645 72526 88669 72590
rect 88733 72526 90426 72590
rect 86231 72510 90426 72526
rect 86231 72446 86493 72510
rect 86557 72446 87581 72510
rect 87645 72446 88669 72510
rect 88733 72446 90426 72510
rect 86231 72430 90426 72446
rect 86231 72366 86493 72430
rect 86557 72366 87581 72430
rect 87645 72366 88669 72430
rect 88733 72366 90426 72430
rect 86231 72365 90426 72366
rect 78237 72359 90426 72365
rect 73811 72350 90426 72359
rect 73811 72286 74525 72350
rect 74589 72286 75613 72350
rect 75677 72286 76701 72350
rect 76765 72286 77789 72350
rect 77853 72286 78877 72350
rect 78941 72286 79965 72350
rect 80029 72286 81053 72350
rect 81117 72286 86493 72350
rect 86557 72286 87581 72350
rect 87645 72286 88669 72350
rect 88733 72286 90426 72350
rect 73811 72270 90426 72286
rect 73811 72206 74525 72270
rect 74589 72206 75613 72270
rect 75677 72206 76701 72270
rect 76765 72206 77789 72270
rect 77853 72206 78877 72270
rect 78941 72206 79965 72270
rect 80029 72206 81053 72270
rect 81117 72206 86493 72270
rect 86557 72206 87581 72270
rect 87645 72206 88669 72270
rect 88733 72206 90426 72270
rect 73811 72169 90426 72206
rect 67270 71638 67646 71656
rect 50682 71278 50748 71279
rect 50682 71214 50683 71278
rect 50747 71214 69124 71278
rect 50682 71213 50748 71214
rect 50682 70655 50748 70656
rect 50682 70591 50683 70655
rect 50747 70591 68505 70655
rect 50682 70590 50748 70591
rect 51122 70260 51420 70341
rect 51122 63876 51199 70260
rect 51343 69399 51420 70260
rect 67273 70131 67646 70151
rect 57424 69855 57713 69986
rect 51343 69101 51442 69399
rect 51343 68680 51420 69101
rect 51343 68623 54435 68680
rect 51343 68387 54000 68623
rect 54236 68387 54435 68623
rect 51343 68340 54435 68387
rect 57424 68351 57473 69855
rect 57617 68566 57713 69855
rect 67273 68566 67307 70131
rect 57617 68534 58466 68566
rect 57617 68351 57993 68534
rect 51343 63913 51420 68340
rect 57424 68298 57993 68351
rect 58229 68298 58466 68534
rect 57424 68277 58466 68298
rect 67181 68277 67307 68566
rect 67273 67260 67307 68277
rect 65854 67258 67307 67260
rect 65854 67022 66001 67258
rect 66237 67022 67307 67258
rect 65854 67020 67307 67022
rect 57419 65393 57659 65433
rect 51343 63906 56959 63913
rect 51343 63876 54008 63906
rect 51122 63850 54008 63876
rect 54244 63850 56959 63906
rect 51122 63770 51426 63850
rect 51381 63706 51426 63770
rect 56930 63706 56959 63850
rect 57419 63889 57454 65393
rect 57598 64890 57659 65393
rect 57856 64890 58386 64891
rect 57598 64889 58386 64890
rect 57598 64653 58003 64889
rect 58239 64653 58386 64889
rect 57598 64651 58386 64653
rect 57598 64650 58022 64651
rect 57598 63889 57659 64650
rect 57419 63832 57659 63889
rect 67273 63907 67307 67020
rect 67611 63907 67646 70131
rect 67273 63888 67646 63907
rect 51381 63670 54008 63706
rect 54244 63670 56959 63706
rect 51381 63658 56959 63670
rect 57850 63460 58380 63462
rect 57850 63224 57997 63460
rect 58233 63372 58380 63460
rect 58233 63308 59732 63372
rect 58233 63224 58380 63308
rect 57850 63222 58380 63224
rect 59606 62895 59732 63308
rect 59606 62831 59616 62895
rect 59680 62831 59732 62895
rect 59606 62815 59732 62831
rect 52380 62812 52446 62813
rect 52380 62748 52381 62812
rect 52445 62748 52446 62812
rect 52380 62747 52446 62748
rect 59606 62751 59616 62815
rect 59680 62751 59732 62815
rect 49371 61921 49437 61922
rect 49371 61857 49372 61921
rect 49436 61857 49437 61921
rect 49371 61856 49437 61857
rect 48613 61393 48679 61394
rect 48613 61329 48614 61393
rect 48678 61329 48679 61393
rect 48613 61328 48679 61329
rect 47885 59963 47951 59964
rect 47885 59899 47886 59963
rect 47950 59899 47951 59963
rect 47885 59898 47951 59899
rect 47024 59373 47090 59374
rect 47024 59309 47025 59373
rect 47089 59309 47090 59373
rect 47024 59308 47090 59309
rect 43698 58698 43764 58699
rect 43698 58634 43699 58698
rect 43763 58634 43764 58698
rect 43698 58633 43764 58634
rect 52381 58218 52445 62747
rect 59606 62735 59732 62751
rect 59606 62671 59616 62735
rect 59680 62671 59732 62735
rect 59606 62654 59732 62671
rect 52970 62469 53036 62470
rect 52970 62405 52971 62469
rect 53035 62405 53036 62469
rect 52970 62404 53036 62405
rect 59608 62422 59734 62444
rect 52380 58217 52446 58218
rect 52380 58153 52381 58217
rect 52445 58153 52446 58217
rect 52380 58152 52446 58153
rect 52971 57873 53035 62404
rect 59608 62358 59626 62422
rect 59690 62358 59734 62422
rect 59608 62342 59734 62358
rect 59608 62278 59626 62342
rect 59690 62278 59734 62342
rect 59608 62262 59734 62278
rect 59608 62198 59626 62262
rect 59690 62198 59734 62262
rect 59608 62182 59734 62198
rect 59608 62118 59626 62182
rect 59690 62118 59734 62182
rect 59608 62102 59734 62118
rect 59608 62038 59626 62102
rect 59690 62038 59734 62102
rect 59608 61993 59734 62038
rect 61855 62073 62385 62075
rect 61855 61993 62002 62073
rect 59608 61929 62002 61993
rect 54696 61922 54760 61923
rect 54695 61921 54761 61922
rect 56333 61921 56399 61922
rect 58566 61921 58632 61922
rect 54695 61857 54696 61921
rect 54760 61857 54761 61921
rect 56317 61857 56334 61921
rect 56398 61857 58567 61921
rect 58631 61857 58663 61921
rect 59608 61897 59708 61929
rect 54695 61856 54761 61857
rect 56333 61856 56399 61857
rect 58566 61856 58632 61857
rect 54279 61394 54343 61397
rect 54278 61393 54344 61394
rect 54278 61329 54279 61393
rect 54343 61329 54344 61393
rect 54278 61328 54344 61329
rect 52970 57872 53036 57873
rect 52970 57808 52971 57872
rect 53035 57808 53036 57872
rect 52970 57807 53036 57808
rect 41954 57201 42020 57202
rect 41954 57137 41955 57201
rect 42019 57137 42020 57201
rect 41954 57136 42020 57137
rect 29932 56822 30017 56886
rect 30081 56822 30172 56886
rect 29932 56806 30172 56822
rect 29932 56742 30017 56806
rect 30081 56789 30172 56806
rect 30081 56787 30390 56789
rect 29932 56726 30043 56742
rect 29932 56662 30017 56726
rect 29932 56646 30043 56662
rect 29932 56582 30017 56646
rect 29932 56566 30043 56582
rect 29932 56502 30017 56566
rect 30279 56551 30390 56787
rect 30081 56549 30390 56551
rect 30081 56502 30172 56549
rect 29932 56486 30172 56502
rect 29932 56422 30017 56486
rect 30081 56422 30172 56486
rect 29932 56351 30172 56422
rect 53175 53774 53241 53775
rect 53175 53710 53176 53774
rect 53240 53710 53241 53774
rect 53175 53709 53241 53710
rect 51815 53352 51879 53354
rect 51814 53351 51880 53352
rect 51814 53287 51815 53351
rect 51879 53287 51880 53351
rect 51814 53286 51880 53287
rect 41353 52730 41594 52731
rect 37856 52728 41594 52730
rect 37856 52492 38003 52728
rect 38239 52492 41594 52728
rect 37856 52490 41594 52492
rect 39394 51634 39634 52490
rect 41353 52085 41594 52490
rect 41353 52021 41399 52085
rect 41463 52021 41594 52085
rect 41353 52005 41594 52021
rect 41353 51941 41399 52005
rect 41463 51941 41594 52005
rect 41353 51925 41594 51941
rect 41353 51861 41399 51925
rect 41463 51861 41594 51925
rect 41353 51845 41594 51861
rect 41353 51781 41399 51845
rect 41463 51781 41594 51845
rect 41353 51765 41594 51781
rect 41353 51701 41399 51765
rect 41463 51701 41594 51765
rect 41353 51641 41594 51701
rect 44700 52087 44828 52111
rect 44700 52023 44709 52087
rect 44773 52025 44828 52087
rect 45857 52075 46387 52077
rect 45857 52025 46004 52075
rect 44773 52023 46004 52025
rect 44700 52007 46004 52023
rect 44700 51943 44709 52007
rect 44773 51943 46004 52007
rect 44700 51927 46004 51943
rect 44700 51863 44709 51927
rect 44773 51897 46004 51927
rect 44773 51863 44828 51897
rect 44700 51847 44828 51863
rect 44700 51783 44709 51847
rect 44773 51783 44828 51847
rect 44700 51767 44828 51783
rect 44700 51703 44709 51767
rect 44773 51703 44828 51767
rect 44700 51680 44828 51703
rect 39394 51570 39491 51634
rect 39555 51570 39634 51634
rect 39394 51483 39634 51570
rect 41860 51463 42390 51465
rect 41860 51227 42007 51463
rect 42243 51410 42390 51463
rect 44708 51450 44836 51483
rect 44699 51446 44836 51450
rect 44699 51410 44716 51446
rect 42243 51382 44716 51410
rect 44780 51410 44836 51446
rect 44780 51382 44847 51410
rect 42243 51366 44847 51382
rect 42243 51302 44716 51366
rect 44780 51302 44847 51366
rect 42243 51286 44847 51302
rect 42243 51282 44716 51286
rect 42243 51227 42390 51282
rect 41860 51225 42390 51227
rect 44699 51222 44716 51282
rect 44780 51282 44847 51286
rect 44780 51222 44836 51282
rect 44699 51219 44836 51222
rect 44708 51210 44836 51219
rect 21870 50928 22333 50930
rect 21870 50692 21983 50928
rect 22219 50692 22333 50928
rect 21870 50634 22333 50692
rect 18903 50616 22333 50634
rect 18903 50552 18939 50616
rect 19003 50552 19019 50616
rect 19083 50552 19099 50616
rect 19163 50552 19179 50616
rect 19243 50552 19259 50616
rect 19323 50552 19339 50616
rect 19403 50552 19419 50616
rect 19483 50552 19499 50616
rect 19563 50552 19579 50616
rect 19643 50552 19659 50616
rect 19723 50552 19739 50616
rect 19803 50552 19819 50616
rect 19883 50552 19899 50616
rect 19963 50552 19979 50616
rect 20043 50552 20059 50616
rect 20123 50552 20139 50616
rect 20203 50552 20219 50616
rect 20283 50552 20299 50616
rect 20363 50552 20379 50616
rect 20443 50552 20459 50616
rect 20523 50552 20539 50616
rect 20603 50552 20619 50616
rect 20683 50552 20699 50616
rect 20763 50552 20779 50616
rect 20843 50552 20859 50616
rect 20923 50552 20939 50616
rect 21003 50552 21019 50616
rect 21083 50552 21099 50616
rect 21163 50552 21179 50616
rect 21243 50552 21259 50616
rect 21323 50552 21339 50616
rect 21403 50552 21419 50616
rect 21483 50552 21499 50616
rect 21563 50552 21579 50616
rect 21643 50552 21659 50616
rect 21723 50552 21739 50616
rect 21803 50552 21819 50616
rect 21883 50552 21899 50616
rect 21963 50552 21979 50616
rect 22043 50552 22059 50616
rect 22123 50552 22139 50616
rect 22203 50552 22333 50616
rect 18903 50536 22333 50552
rect 18903 50535 22239 50536
rect 44672 50485 44800 50515
rect 39403 50405 39636 50483
rect 39403 50341 39491 50405
rect 39555 50341 39636 50405
rect 44672 50421 44713 50485
rect 44777 50421 44800 50485
rect 44672 50405 44800 50421
rect 39403 49832 39636 50341
rect 41352 50296 41585 50376
rect 41352 50232 41381 50296
rect 41445 50232 41585 50296
rect 41352 50216 41585 50232
rect 41352 50152 41381 50216
rect 41445 50152 41585 50216
rect 41352 50136 41585 50152
rect 41352 50072 41381 50136
rect 41445 50072 41585 50136
rect 44672 50341 44713 50405
rect 44777 50352 44800 50405
rect 45377 50352 45505 51897
rect 45857 51839 46004 51897
rect 46240 51839 46387 52075
rect 45857 51837 46387 51839
rect 51815 51555 51879 53286
rect 51814 51554 51880 51555
rect 51814 51490 51815 51554
rect 51879 51490 51880 51554
rect 51814 51489 51880 51490
rect 44777 50341 45505 50352
rect 44672 50325 45505 50341
rect 44672 50261 44713 50325
rect 44777 50261 45505 50325
rect 44672 50245 45505 50261
rect 44672 50181 44713 50245
rect 44777 50224 45505 50245
rect 44777 50181 44800 50224
rect 44672 50165 44800 50181
rect 44672 50101 44713 50165
rect 44777 50101 44800 50165
rect 44672 50075 44800 50101
rect 41352 49832 41585 50072
rect 41856 49838 42386 49840
rect 41856 49832 42003 49838
rect 37848 49830 38378 49832
rect 37848 49594 37995 49830
rect 38231 49821 38378 49830
rect 38234 49597 38378 49821
rect 38231 49594 38378 49597
rect 37848 49592 38378 49594
rect 39403 49602 42003 49832
rect 42239 49787 42386 49838
rect 44711 49787 44839 49878
rect 42239 49659 44839 49787
rect 42239 49602 42386 49659
rect 44711 49617 44839 49659
rect 39403 49600 42386 49602
rect 39403 49599 42247 49600
rect 29866 49534 30396 49536
rect 29866 49298 30013 49534
rect 30249 49455 30396 49534
rect 31644 49502 31726 49505
rect 31644 49455 31653 49502
rect 30249 49438 31653 49455
rect 31717 49455 31726 49502
rect 31717 49438 31778 49455
rect 30249 49422 31778 49438
rect 30249 49358 31653 49422
rect 31717 49358 31778 49422
rect 30249 49342 31778 49358
rect 30249 49327 31653 49342
rect 30249 49298 30396 49327
rect 29866 49296 30396 49298
rect 31644 49278 31653 49327
rect 31717 49327 31778 49342
rect 31717 49278 31726 49327
rect 31644 49262 31726 49278
rect 31644 49198 31653 49262
rect 31717 49198 31726 49262
rect 31644 49196 31726 49198
rect 39403 48992 39636 49599
rect 45377 49335 45505 50224
rect 45770 49687 45834 49688
rect 45769 49686 45835 49687
rect 45769 49622 45770 49686
rect 45834 49622 45835 49686
rect 45769 49621 45835 49622
rect 31641 48963 31730 48968
rect 31641 48899 31653 48963
rect 31717 48915 31730 48963
rect 33858 48937 34388 48939
rect 33858 48915 34005 48937
rect 31717 48899 34005 48915
rect 31641 48883 34005 48899
rect 31641 48819 31653 48883
rect 31717 48819 34005 48883
rect 31641 48803 34005 48819
rect 31641 48739 31653 48803
rect 31717 48787 34005 48803
rect 31717 48739 31730 48787
rect 31641 48735 31730 48739
rect 33858 48701 34005 48787
rect 34241 48701 34388 48937
rect 39403 48928 39491 48992
rect 39555 48928 39636 48992
rect 39403 48833 39636 48928
rect 44696 49207 45505 49335
rect 33858 48699 34388 48701
rect 44696 48719 44824 49207
rect 45116 48894 45182 48895
rect 45116 48830 45117 48894
rect 45181 48830 45182 48894
rect 45116 48829 45182 48830
rect 44696 48655 44701 48719
rect 44765 48655 44824 48719
rect 44696 48639 44824 48655
rect 44696 48575 44701 48639
rect 44765 48575 44824 48639
rect 44696 48559 44824 48575
rect 44696 48495 44701 48559
rect 44765 48495 44824 48559
rect 44696 48463 44824 48495
rect 44660 48255 44788 48286
rect 44660 48191 44705 48255
rect 44769 48191 44788 48255
rect 44660 48175 44788 48191
rect 44660 48111 44705 48175
rect 44769 48111 44788 48175
rect 44660 48095 44788 48111
rect 44660 48031 44705 48095
rect 44769 48031 44788 48095
rect 39402 47763 39642 47876
rect 39402 47753 39491 47763
rect 38283 47752 39491 47753
rect 37855 47750 39491 47752
rect 17889 47734 18352 47736
rect 17889 47498 18002 47734
rect 18238 47732 18352 47734
rect 18238 47608 22324 47732
rect 18238 47544 18945 47608
rect 19009 47544 19025 47608
rect 19089 47544 19105 47608
rect 19169 47544 19185 47608
rect 19249 47544 19265 47608
rect 19329 47544 19345 47608
rect 19409 47544 19425 47608
rect 19489 47544 19505 47608
rect 19569 47544 19585 47608
rect 19649 47544 19665 47608
rect 19729 47544 19745 47608
rect 19809 47544 19825 47608
rect 19889 47544 19905 47608
rect 19969 47544 19985 47608
rect 20049 47544 20065 47608
rect 20129 47544 20145 47608
rect 20209 47544 20225 47608
rect 20289 47544 20305 47608
rect 20369 47544 20385 47608
rect 20449 47544 20465 47608
rect 20529 47544 20545 47608
rect 20609 47544 20625 47608
rect 20689 47544 20705 47608
rect 20769 47544 20785 47608
rect 20849 47544 20865 47608
rect 20929 47544 20945 47608
rect 21009 47544 21025 47608
rect 21089 47544 21105 47608
rect 21169 47544 21185 47608
rect 21249 47544 21265 47608
rect 21329 47544 21345 47608
rect 21409 47544 21425 47608
rect 21489 47544 21505 47608
rect 21569 47544 21585 47608
rect 21649 47544 21665 47608
rect 21729 47544 21745 47608
rect 21809 47544 21825 47608
rect 21889 47544 21905 47608
rect 21969 47544 21985 47608
rect 22049 47544 22065 47608
rect 22129 47544 22145 47608
rect 22209 47544 22324 47608
rect 18238 47498 22324 47544
rect 37855 47514 38002 47750
rect 38238 47699 39491 47750
rect 39555 47699 39642 47763
rect 38238 47514 39642 47699
rect 37855 47513 39642 47514
rect 41368 47659 41601 47661
rect 41857 47659 42387 47661
rect 41368 47655 42004 47659
rect 41368 47591 41370 47655
rect 41434 47591 42004 47655
rect 41368 47575 42004 47591
rect 37855 47512 38385 47513
rect 17889 47496 22324 47498
rect 41368 47511 41370 47575
rect 41434 47511 42004 47575
rect 41368 47495 42004 47511
rect 41368 47431 41370 47495
rect 41434 47431 42004 47495
rect 41368 47426 42004 47431
rect 41857 47423 42004 47426
rect 42240 47614 42387 47659
rect 44660 47614 44788 48031
rect 42240 47486 44788 47614
rect 45117 47541 45181 48829
rect 45770 47910 45834 49621
rect 45769 47909 45835 47910
rect 45769 47845 45770 47909
rect 45834 47845 45835 47909
rect 45769 47844 45835 47845
rect 45116 47540 45182 47541
rect 42240 47423 42387 47486
rect 41857 47421 42387 47423
rect 40494 46746 40560 46747
rect 40494 46682 40495 46746
rect 40559 46682 40560 46746
rect 40494 46681 40560 46682
rect 40495 44674 40559 46681
rect 43209 46606 43337 47486
rect 45116 47476 45117 47540
rect 45181 47476 45182 47540
rect 45116 47475 45182 47476
rect 45117 47464 45181 47475
rect 44704 47299 44776 47300
rect 44704 47281 44836 47299
rect 44704 47217 44708 47281
rect 44772 47217 44836 47281
rect 44704 47201 44836 47217
rect 44704 47137 44708 47201
rect 44772 47137 44836 47201
rect 44704 47130 44836 47137
rect 45848 47174 46378 47176
rect 45848 47130 45995 47174
rect 44704 47121 45995 47130
rect 44704 47057 44708 47121
rect 44772 47057 45995 47121
rect 44704 47041 45995 47057
rect 44704 46977 44708 47041
rect 44772 47002 45995 47041
rect 44772 46977 44836 47002
rect 44704 46961 44836 46977
rect 44704 46897 44708 46961
rect 44772 46897 44836 46961
rect 45848 46938 45995 47002
rect 46231 46938 46378 47174
rect 45848 46936 46378 46938
rect 44704 46878 44836 46897
rect 44708 46859 44836 46878
rect 44694 46645 44822 46673
rect 44694 46606 44705 46645
rect 43209 46581 44705 46606
rect 44769 46581 44822 46645
rect 43209 46565 44822 46581
rect 43209 46501 44705 46565
rect 44769 46501 44822 46565
rect 43209 46485 44822 46501
rect 43209 46478 44705 46485
rect 44694 46421 44705 46478
rect 44769 46421 44822 46485
rect 44694 46372 44822 46421
rect 40494 44673 40560 44674
rect 40494 44609 40495 44673
rect 40559 44609 40560 44673
rect 40494 44608 40560 44609
rect 21876 43253 22339 43255
rect 21876 43088 21989 43253
rect 18925 43080 21989 43088
rect 18925 43016 18947 43080
rect 19011 43016 19027 43080
rect 19091 43016 19107 43080
rect 19171 43016 19187 43080
rect 19251 43016 19267 43080
rect 19331 43016 19347 43080
rect 19411 43016 19427 43080
rect 19491 43016 19507 43080
rect 19571 43016 19587 43080
rect 19651 43016 19667 43080
rect 19731 43016 19747 43080
rect 19811 43016 19827 43080
rect 19891 43016 19907 43080
rect 19971 43016 19987 43080
rect 20051 43016 20067 43080
rect 20131 43016 20147 43080
rect 20211 43016 20227 43080
rect 20291 43016 20307 43080
rect 20371 43016 20387 43080
rect 20451 43016 20467 43080
rect 20531 43016 20547 43080
rect 20611 43016 20627 43080
rect 20691 43016 20707 43080
rect 20771 43016 20787 43080
rect 20851 43016 20867 43080
rect 20931 43016 20947 43080
rect 21011 43016 21027 43080
rect 21091 43016 21107 43080
rect 21171 43016 21187 43080
rect 21251 43016 21267 43080
rect 21331 43016 21347 43080
rect 21411 43016 21427 43080
rect 21491 43016 21507 43080
rect 21571 43016 21587 43080
rect 21651 43016 21667 43080
rect 21731 43016 21747 43080
rect 21811 43016 21827 43080
rect 21891 43016 21907 43080
rect 21971 43016 21987 43080
rect 22225 43017 22339 43253
rect 51815 43066 51879 51489
rect 53176 50878 53240 53709
rect 53175 50877 53241 50878
rect 53175 50813 53176 50877
rect 53240 50813 53241 50877
rect 53175 50812 53241 50813
rect 53176 43066 53240 50812
rect 54279 43536 54343 61328
rect 54278 43535 54344 43536
rect 54278 43471 54279 43535
rect 54343 43471 54344 43535
rect 54278 43470 54344 43471
rect 54696 43235 54760 61856
rect 61855 61837 62002 61929
rect 62238 61837 62385 62073
rect 61855 61835 62385 61837
rect 56333 61392 56399 61393
rect 59089 61392 59155 61393
rect 56333 61328 56334 61392
rect 56398 61328 59090 61392
rect 59154 61328 59188 61392
rect 56333 61327 56399 61328
rect 59089 61327 59155 61328
rect 59261 61157 59327 61172
rect 57851 61115 58381 61117
rect 57851 60879 57998 61115
rect 58234 61018 58381 61115
rect 59261 61093 59262 61157
rect 59326 61093 59327 61157
rect 59261 61077 59327 61093
rect 59261 61018 59262 61077
rect 58234 61013 59262 61018
rect 59326 61013 59327 61077
rect 58234 60997 59327 61013
rect 58234 60954 59262 60997
rect 58234 60879 58381 60954
rect 59261 60933 59262 60954
rect 59326 60933 59327 60997
rect 59261 60919 59327 60933
rect 57851 60877 58381 60879
rect 59263 60691 59327 60702
rect 59262 60673 59328 60691
rect 59262 60609 59263 60673
rect 59327 60609 59328 60673
rect 59262 60593 59328 60609
rect 59262 60529 59263 60593
rect 59327 60589 59328 60593
rect 61862 60680 62392 60682
rect 61862 60589 62009 60680
rect 59327 60529 62009 60589
rect 59262 60525 62009 60529
rect 59262 60513 59328 60525
rect 59262 60449 59263 60513
rect 59327 60449 59328 60513
rect 59262 60433 59328 60449
rect 61862 60444 62009 60525
rect 62245 60444 62392 60680
rect 61862 60442 62392 60444
rect 59262 60369 59263 60433
rect 59327 60369 59328 60433
rect 59262 60353 59328 60369
rect 59262 60289 59263 60353
rect 59327 60289 59328 60353
rect 59262 60271 59328 60289
rect 60758 60117 60877 60137
rect 62273 60127 62337 60442
rect 60675 60116 60906 60117
rect 60675 60052 60678 60116
rect 60742 60052 60758 60116
rect 60822 60052 60838 60116
rect 60902 60052 60906 60116
rect 60675 60051 60906 60052
rect 62148 60115 62446 60127
rect 62723 60120 62842 60137
rect 62148 60051 62185 60115
rect 62249 60051 62265 60115
rect 62329 60051 62345 60115
rect 62409 60051 62446 60115
rect 57868 60036 58398 60038
rect 57868 59800 58015 60036
rect 58251 59979 58398 60036
rect 60758 59979 60877 60051
rect 62148 60039 62446 60051
rect 62667 60116 62896 60120
rect 62667 60052 62669 60116
rect 62733 60052 62749 60116
rect 62813 60052 62829 60116
rect 62893 60052 62896 60116
rect 64075 60112 64194 60147
rect 66739 60114 66858 60122
rect 62667 60048 62896 60052
rect 64029 60108 64252 60112
rect 62723 59979 62842 60048
rect 64029 60044 64068 60108
rect 64132 60044 64148 60108
rect 64212 60044 64252 60108
rect 66668 60111 66897 60114
rect 64029 60041 64252 60044
rect 65852 60048 66382 60050
rect 64075 59979 64194 60041
rect 65852 59979 65999 60048
rect 58251 59860 65999 59979
rect 58251 59800 58398 59860
rect 65852 59812 65999 59860
rect 66235 59979 66382 60048
rect 66668 60047 66670 60111
rect 66734 60047 66750 60111
rect 66814 60047 66830 60111
rect 66894 60047 66897 60111
rect 66668 60044 66897 60047
rect 66739 59979 66858 60044
rect 66235 59860 66858 59979
rect 66235 59812 66382 59860
rect 65852 59810 66382 59812
rect 57868 59798 58398 59800
rect 60214 59666 60335 59695
rect 60214 59602 60242 59666
rect 60306 59602 60335 59666
rect 60214 59574 60335 59602
rect 64596 59635 64717 59664
rect 60215 59440 60334 59574
rect 64596 59571 64624 59635
rect 64688 59571 64717 59635
rect 64596 59543 64717 59571
rect 66163 59644 66284 59673
rect 66163 59580 66191 59644
rect 66255 59580 66284 59644
rect 66163 59552 66284 59580
rect 61868 59502 62398 59504
rect 61868 59440 62015 59502
rect 60140 59321 62015 59440
rect 61868 59266 62015 59321
rect 62251 59440 62398 59502
rect 64597 59440 64716 59543
rect 66164 59440 66283 59552
rect 62251 59321 66283 59440
rect 62251 59266 62398 59321
rect 61868 59264 62398 59266
rect 61795 55472 61859 56194
rect 65059 55834 65123 56194
rect 65058 55833 65124 55834
rect 65058 55769 65059 55833
rect 65123 55769 65124 55833
rect 65058 55768 65124 55769
rect 61038 55408 61859 55472
rect 62035 55412 62833 55476
rect 64085 55412 64883 55476
rect 65059 55472 65123 55768
rect 61795 55394 61859 55408
rect 65059 55408 65880 55472
rect 68441 55414 68505 70591
rect 68440 55413 68506 55414
rect 65059 55394 65123 55408
rect 68440 55349 68441 55413
rect 68505 55349 68506 55413
rect 68440 55348 68506 55349
rect 60792 54411 60856 55209
rect 61447 54454 61513 54455
rect 61447 54390 61448 54454
rect 61512 54390 61799 54454
rect 63059 54416 63123 55214
rect 63795 54416 63859 55214
rect 65421 54459 65487 54460
rect 65122 54395 65422 54459
rect 65486 54395 65487 54459
rect 66062 54411 66126 55209
rect 65421 54394 65487 54395
rect 61447 54389 61513 54390
rect 60419 54327 60485 54328
rect 60419 54263 60420 54327
rect 60484 54263 60837 54327
rect 60419 54262 60485 54263
rect 60792 53411 60856 54209
rect 61795 53418 61859 54216
rect 63059 53416 63123 54214
rect 63795 53416 63859 54214
rect 65059 53418 65123 54216
rect 66062 53411 66126 54209
rect 60792 52411 60856 53189
rect 62061 52400 62125 53198
rect 63059 52416 63123 53214
rect 63795 52416 63859 53214
rect 64793 52400 64857 53198
rect 66062 52411 66126 53209
rect 67726 52826 67792 52827
rect 67726 52762 67727 52826
rect 67791 52762 67792 52826
rect 67726 52761 67792 52762
rect 60792 51411 60856 52209
rect 63059 51416 63123 52214
rect 63795 51416 63859 52214
rect 66062 51411 66126 52209
rect 61797 51210 61861 51222
rect 65057 51210 65121 51222
rect 61060 51146 61861 51210
rect 62060 51146 62858 51210
rect 64060 51146 64858 51210
rect 65057 51146 65858 51210
rect 61797 50424 61861 51146
rect 65057 50424 65121 51146
rect 64694 48870 64760 48871
rect 64694 48806 64695 48870
rect 64759 48806 64760 48870
rect 64694 48805 64760 48806
rect 62812 48617 62876 48739
rect 62808 48604 62878 48617
rect 62808 48540 62811 48604
rect 62875 48540 62878 48604
rect 64359 48615 64425 48616
rect 64359 48551 64360 48615
rect 64424 48551 64425 48615
rect 64359 48550 64425 48551
rect 62808 48524 62878 48540
rect 62808 48460 62811 48524
rect 62875 48460 62878 48524
rect 62808 48444 62878 48460
rect 62808 48380 62811 48444
rect 62875 48380 62878 48444
rect 62808 48364 62878 48380
rect 62808 48300 62811 48364
rect 62875 48300 62878 48364
rect 62808 48284 62878 48300
rect 62808 48220 62811 48284
rect 62875 48220 62878 48284
rect 62808 48207 62878 48220
rect 61873 47179 62338 47182
rect 61873 47173 61987 47179
rect 62223 47173 62338 47179
rect 61873 46949 61913 47173
rect 62297 46949 62338 47173
rect 62812 47086 62876 48207
rect 64360 47910 64424 48550
rect 64359 47909 64425 47910
rect 64359 47845 64360 47909
rect 64424 47845 64425 47909
rect 64359 47844 64425 47845
rect 62811 47085 62877 47086
rect 62811 47021 62812 47085
rect 62876 47021 62877 47085
rect 62811 47020 62877 47021
rect 61873 46943 61987 46949
rect 62223 46943 62338 46949
rect 61873 46940 62338 46943
rect 64695 46296 64759 48805
rect 65222 48552 65288 48553
rect 65222 48488 65223 48552
rect 65287 48488 65288 48552
rect 65222 48487 65288 48488
rect 65223 46747 65287 48487
rect 65868 47515 66331 47517
rect 65868 47355 65981 47515
rect 65868 47291 65887 47355
rect 65951 47291 65967 47355
rect 65868 47279 65981 47291
rect 66217 47279 66331 47515
rect 65868 47277 66331 47279
rect 65880 47267 66038 47277
rect 65222 46746 65288 46747
rect 65222 46682 65223 46746
rect 65287 46682 65288 46746
rect 65222 46681 65288 46682
rect 65223 46673 65287 46681
rect 64694 46295 64760 46296
rect 64694 46231 64695 46295
rect 64759 46231 64760 46295
rect 64694 46230 64760 46231
rect 67727 44972 67791 52761
rect 68441 50373 68505 55348
rect 69060 54795 69124 71214
rect 73809 70747 90321 70789
rect 73809 70683 75070 70747
rect 75134 70683 76158 70747
rect 76222 70683 77246 70747
rect 77310 70683 78334 70747
rect 78398 70683 79422 70747
rect 79486 70683 81598 70747
rect 81662 70683 82686 70747
rect 82750 70683 83774 70747
rect 83838 70683 84862 70747
rect 84926 70683 85950 70747
rect 86014 70683 87038 70747
rect 87102 70683 88126 70747
rect 88190 70739 90321 70747
rect 88190 70683 90384 70739
rect 73809 70667 90384 70683
rect 73809 70604 75070 70667
rect 73809 70368 74004 70604
rect 74240 70603 75070 70604
rect 75134 70603 76158 70667
rect 76222 70603 77246 70667
rect 77310 70603 78334 70667
rect 78398 70603 79422 70667
rect 79486 70603 81598 70667
rect 81662 70603 82686 70667
rect 82750 70603 83774 70667
rect 83838 70603 84862 70667
rect 84926 70603 85950 70667
rect 86014 70603 87038 70667
rect 87102 70603 88126 70667
rect 88190 70603 90384 70667
rect 74240 70597 90384 70603
rect 74240 70587 82000 70597
rect 74240 70523 75070 70587
rect 75134 70523 76158 70587
rect 76222 70523 77246 70587
rect 77310 70523 78334 70587
rect 78398 70523 79422 70587
rect 79486 70523 81598 70587
rect 81662 70523 82000 70587
rect 74240 70507 82000 70523
rect 74240 70443 75070 70507
rect 75134 70443 76158 70507
rect 76222 70443 77246 70507
rect 77310 70443 78334 70507
rect 78398 70443 79422 70507
rect 79486 70443 81598 70507
rect 81662 70443 82000 70507
rect 74240 70427 82000 70443
rect 74240 70368 75070 70427
rect 73809 70363 75070 70368
rect 75134 70363 76158 70427
rect 76222 70363 77246 70427
rect 77310 70363 78334 70427
rect 78398 70363 79422 70427
rect 79486 70363 81598 70427
rect 81662 70363 82000 70427
rect 73809 70361 82000 70363
rect 82236 70593 90384 70597
rect 82236 70587 90003 70593
rect 82236 70523 82686 70587
rect 82750 70523 83774 70587
rect 83838 70523 84862 70587
rect 84926 70523 85950 70587
rect 86014 70523 87038 70587
rect 87102 70523 88126 70587
rect 88190 70523 90003 70587
rect 82236 70507 90003 70523
rect 82236 70443 82686 70507
rect 82750 70443 83774 70507
rect 83838 70443 84862 70507
rect 84926 70443 85950 70507
rect 86014 70443 87038 70507
rect 87102 70443 88126 70507
rect 88190 70443 90003 70507
rect 82236 70427 90003 70443
rect 82236 70363 82686 70427
rect 82750 70363 83774 70427
rect 83838 70363 84862 70427
rect 84926 70363 85950 70427
rect 86014 70363 87038 70427
rect 87102 70363 88126 70427
rect 88190 70363 90003 70427
rect 82236 70361 90003 70363
rect 73809 70357 90003 70361
rect 90239 70357 90384 70593
rect 73809 70347 90384 70357
rect 73809 70283 75070 70347
rect 75134 70283 76158 70347
rect 76222 70283 77246 70347
rect 77310 70283 78334 70347
rect 78398 70283 79422 70347
rect 79486 70283 81598 70347
rect 81662 70283 82686 70347
rect 82750 70283 83774 70347
rect 83838 70283 84862 70347
rect 84926 70283 85950 70347
rect 86014 70283 87038 70347
rect 87102 70283 88126 70347
rect 88190 70283 90384 70347
rect 73809 70267 90384 70283
rect 73809 70203 75070 70267
rect 75134 70203 76158 70267
rect 76222 70203 77246 70267
rect 77310 70203 78334 70267
rect 78398 70203 79422 70267
rect 79486 70203 81598 70267
rect 81662 70203 82686 70267
rect 82750 70203 83774 70267
rect 83838 70203 84862 70267
rect 84926 70203 85950 70267
rect 86014 70203 87038 70267
rect 87102 70203 88126 70267
rect 88190 70211 90384 70267
rect 88190 70203 90321 70211
rect 73809 70169 90321 70203
rect 75338 69770 75404 69771
rect 75338 69706 75339 69770
rect 75403 69706 75404 69770
rect 75338 69705 75404 69706
rect 75884 69770 75950 69771
rect 75884 69706 75885 69770
rect 75949 69706 75950 69770
rect 83499 69764 83565 69765
rect 75884 69705 75950 69706
rect 76430 69761 76496 69762
rect 75339 68724 75403 69705
rect 75885 69095 75949 69705
rect 76430 69697 76431 69761
rect 76495 69697 76496 69761
rect 76430 69696 76496 69697
rect 76975 69760 77041 69761
rect 76975 69696 76976 69760
rect 77040 69696 77041 69760
rect 82956 69760 83022 69761
rect 80238 69749 80304 69750
rect 75884 69094 75950 69095
rect 75884 69030 75885 69094
rect 75949 69030 75950 69094
rect 75884 69029 75950 69030
rect 75338 68723 75404 68724
rect 75338 68659 75339 68723
rect 75403 68659 75404 68723
rect 75338 68658 75404 68659
rect 75339 62459 75403 68658
rect 70924 62458 70990 62459
rect 70924 62394 70925 62458
rect 70989 62394 70990 62458
rect 70924 62393 70990 62394
rect 75338 62458 75404 62459
rect 75338 62394 75339 62458
rect 75403 62394 75404 62458
rect 75338 62393 75404 62394
rect 70925 55414 70989 62393
rect 75885 61884 75949 69029
rect 76431 65034 76495 69696
rect 76975 69695 77041 69696
rect 78606 69748 78672 69749
rect 76976 65405 77040 69695
rect 78606 69684 78607 69748
rect 78671 69684 78672 69748
rect 78606 69683 78672 69684
rect 79149 69745 79215 69746
rect 76975 65404 77041 65405
rect 76975 65340 76976 65404
rect 77040 65340 77041 65404
rect 76975 65339 77041 65340
rect 76430 65033 76496 65034
rect 76430 64969 76431 65033
rect 76495 64969 76496 65033
rect 76430 64968 76496 64969
rect 71679 61883 71745 61884
rect 71679 61819 71680 61883
rect 71744 61819 71745 61883
rect 71679 61818 71745 61819
rect 75884 61883 75950 61884
rect 75884 61819 75885 61883
rect 75949 61819 75950 61883
rect 75884 61818 75950 61819
rect 70924 55413 70990 55414
rect 70924 55349 70925 55413
rect 70989 55349 70990 55413
rect 70924 55348 70990 55349
rect 71680 54795 71744 61818
rect 76431 61333 76495 64968
rect 72323 61332 72389 61333
rect 72323 61268 72324 61332
rect 72388 61268 72389 61332
rect 72323 61267 72389 61268
rect 76430 61332 76496 61333
rect 76430 61268 76431 61332
rect 76495 61268 76496 61332
rect 76430 61267 76496 61268
rect 69059 54794 69125 54795
rect 69059 54730 69060 54794
rect 69124 54730 69125 54794
rect 69059 54729 69125 54730
rect 71679 54794 71745 54795
rect 71679 54730 71680 54794
rect 71744 54730 71745 54794
rect 71679 54729 71745 54730
rect 69060 52827 69124 54729
rect 69059 52826 69125 52827
rect 69059 52762 69060 52826
rect 69124 52762 69125 52826
rect 69059 52761 69125 52762
rect 69060 52756 69124 52761
rect 68440 50372 68506 50373
rect 68440 50308 68441 50372
rect 68505 50308 68506 50372
rect 68440 50307 68506 50308
rect 68930 50372 68996 50373
rect 68930 50308 68931 50372
rect 68995 50308 68996 50372
rect 68930 50307 68996 50308
rect 68441 50302 68505 50307
rect 68174 48225 68238 48231
rect 68173 48224 68239 48225
rect 68173 48160 68174 48224
rect 68238 48160 68239 48224
rect 68173 48159 68239 48160
rect 67726 44908 67792 44972
rect 68174 44908 68238 48159
rect 68931 46939 68995 50307
rect 70943 50031 71009 50032
rect 70943 49967 70944 50031
rect 71008 49967 71009 50031
rect 70943 49966 71009 49967
rect 70359 49620 70425 49621
rect 70359 49556 70360 49620
rect 70424 49556 70425 49620
rect 70359 49555 70425 49556
rect 69682 47233 69746 47242
rect 69681 47232 69747 47233
rect 69681 47168 69682 47232
rect 69746 47168 69747 47232
rect 69681 47167 69747 47168
rect 68930 46938 68996 46939
rect 68569 46937 68635 46938
rect 68569 46873 68570 46937
rect 68634 46873 68635 46937
rect 68930 46874 68931 46938
rect 68995 46874 68996 46938
rect 68930 46873 68996 46874
rect 68569 46872 68635 46873
rect 67726 44842 68238 44908
rect 68174 44357 68238 44842
rect 68173 44356 68239 44357
rect 68173 44292 68174 44356
rect 68238 44292 68239 44356
rect 68173 44291 68239 44292
rect 68570 43826 68634 46872
rect 69166 45678 69230 45686
rect 69165 45677 69231 45678
rect 69165 45613 69166 45677
rect 69230 45613 69231 45677
rect 69165 45612 69231 45613
rect 68569 43825 68635 43826
rect 68569 43761 68570 43825
rect 68634 43761 68635 43825
rect 68569 43760 68635 43761
rect 61891 43253 62354 43255
rect 54695 43234 54761 43235
rect 54695 43170 54696 43234
rect 54760 43170 54761 43234
rect 54695 43169 54761 43170
rect 61891 43194 62004 43253
rect 62240 43194 62354 43253
rect 22051 43016 22067 43017
rect 22131 43016 22147 43017
rect 22211 43016 22339 43017
rect 18925 43015 22339 43016
rect 51814 43065 51880 43066
rect 18925 43008 22234 43015
rect 51814 43001 51815 43065
rect 51879 43001 51880 43065
rect 51814 43000 51880 43001
rect 53175 43065 53241 43066
rect 53175 43001 53176 43065
rect 53240 43001 53241 43065
rect 53175 43000 53241 43001
rect 29856 41983 30386 41985
rect 29856 41747 30003 41983
rect 30239 41935 30386 41983
rect 31641 41935 31708 41945
rect 30239 41908 31716 41935
rect 30239 41844 31642 41908
rect 31706 41844 31716 41908
rect 30239 41828 31716 41844
rect 30239 41807 31642 41828
rect 30239 41747 30386 41807
rect 29856 41745 30386 41747
rect 31641 41764 31642 41807
rect 31706 41807 31716 41828
rect 53882 41884 54347 41887
rect 53882 41878 53996 41884
rect 54232 41878 54347 41884
rect 31706 41764 31708 41807
rect 31641 41748 31708 41764
rect 31641 41684 31642 41748
rect 31706 41684 31708 41748
rect 31641 41648 31708 41684
rect 53882 41654 53922 41878
rect 54306 41654 54347 41878
rect 53882 41648 53996 41654
rect 54232 41648 54347 41654
rect 53882 41645 54347 41648
rect 31643 41420 31717 41427
rect 31643 41358 31648 41420
rect 31640 41356 31648 41358
rect 31712 41358 31717 41420
rect 31712 41356 32356 41358
rect 31640 41340 32356 41356
rect 31640 41276 31648 41340
rect 31712 41276 32356 41340
rect 31640 41260 32356 41276
rect 31640 41230 31648 41260
rect 31643 41196 31648 41230
rect 31712 41230 32356 41260
rect 31712 41196 31717 41230
rect 31643 41190 31717 41196
rect 17890 40220 18353 40222
rect 17890 39984 18003 40220
rect 18239 40100 18353 40220
rect 18239 40098 22237 40100
rect 18239 40085 22243 40098
rect 18239 40021 18949 40085
rect 19013 40021 19029 40085
rect 19093 40021 19109 40085
rect 19173 40021 19189 40085
rect 19253 40021 19269 40085
rect 19333 40021 19349 40085
rect 19413 40021 19429 40085
rect 19493 40021 19509 40085
rect 19573 40021 19589 40085
rect 19653 40021 19669 40085
rect 19733 40021 19749 40085
rect 19813 40021 19829 40085
rect 19893 40021 19909 40085
rect 19973 40021 19989 40085
rect 20053 40021 20069 40085
rect 20133 40021 20149 40085
rect 20213 40021 20229 40085
rect 20293 40021 20309 40085
rect 20373 40021 20389 40085
rect 20453 40021 20469 40085
rect 20533 40021 20549 40085
rect 20613 40021 20629 40085
rect 20693 40021 20709 40085
rect 20773 40021 20789 40085
rect 20853 40021 20869 40085
rect 20933 40021 20949 40085
rect 21013 40021 21029 40085
rect 21093 40021 21109 40085
rect 21173 40021 21189 40085
rect 21253 40021 21269 40085
rect 21333 40021 21349 40085
rect 21413 40021 21429 40085
rect 21493 40021 21509 40085
rect 21573 40021 21589 40085
rect 21653 40021 21669 40085
rect 21733 40021 21749 40085
rect 21813 40021 21829 40085
rect 21893 40021 21909 40085
rect 21973 40021 21989 40085
rect 22053 40021 22069 40085
rect 22133 40021 22149 40085
rect 22213 40021 22243 40085
rect 18239 40008 22243 40021
rect 18239 40006 22237 40008
rect 18239 39984 18353 40006
rect 17890 39982 18353 39984
rect 32228 39467 32356 41230
rect 38375 41167 39395 41231
rect 40975 41167 41995 41231
rect 43575 41167 44595 41231
rect 46677 41179 46743 41180
rect 46182 41115 46678 41179
rect 46742 41115 46743 41179
rect 46677 41114 46743 41115
rect 54696 41011 54760 43169
rect 61891 43050 61967 43194
rect 62271 43050 62354 43194
rect 61891 43017 62004 43050
rect 62240 43017 62354 43050
rect 61891 43015 62354 43017
rect 67325 43080 67391 43081
rect 67325 43016 67326 43080
rect 67390 43016 67391 43080
rect 67325 43015 67391 43016
rect 55589 42932 55655 42933
rect 55589 42868 55590 42932
rect 55654 42868 55655 42932
rect 55589 42867 55655 42868
rect 53166 40947 54760 41011
rect 33841 39510 34371 39512
rect 33841 39467 33988 39510
rect 32228 39339 33988 39467
rect 29863 38497 30393 38499
rect 29863 38261 30010 38497
rect 30246 38447 30393 38497
rect 31576 38447 31651 38469
rect 30246 38435 31680 38447
rect 30246 38371 31581 38435
rect 31645 38371 31680 38435
rect 30246 38355 31680 38371
rect 30246 38319 31581 38355
rect 30246 38261 30393 38319
rect 29863 38259 30393 38261
rect 31576 38291 31581 38319
rect 31645 38319 31680 38355
rect 31645 38291 31651 38319
rect 31576 38275 31651 38291
rect 31576 38211 31581 38275
rect 31645 38211 31651 38275
rect 31576 38178 31651 38211
rect 31575 37941 31649 37948
rect 31575 37896 31580 37941
rect 31574 37877 31580 37896
rect 31644 37896 31649 37941
rect 32228 37896 32356 39339
rect 33841 39274 33988 39339
rect 34224 39274 34371 39510
rect 33841 39272 34371 39274
rect 37081 38902 37145 39922
rect 42909 39392 43039 39425
rect 42909 39328 42942 39392
rect 43006 39328 43039 39392
rect 42909 39295 43039 39328
rect 42910 38914 43038 39295
rect 45839 38895 45903 39915
rect 49876 39832 50339 39834
rect 49876 39596 49989 39832
rect 50225 39730 50339 39832
rect 51307 39730 51373 39731
rect 50225 39666 51308 39730
rect 51372 39666 51373 39730
rect 50225 39596 50339 39666
rect 51307 39665 51373 39666
rect 49876 39594 50339 39596
rect 53166 39477 53230 40947
rect 53893 40470 54356 40472
rect 53893 40234 54006 40470
rect 54242 40234 54356 40470
rect 53893 40232 54356 40234
rect 53584 40227 53650 40228
rect 53584 40163 53585 40227
rect 53649 40163 53650 40227
rect 53584 40162 53650 40163
rect 53165 39476 53231 39477
rect 53165 39412 53166 39476
rect 53230 39412 53231 39476
rect 53165 39411 53231 39412
rect 49873 38472 50336 38474
rect 49873 38236 49986 38472
rect 50222 38367 50336 38472
rect 52191 38435 52263 38469
rect 52191 38371 52195 38435
rect 52259 38371 52263 38435
rect 52191 38367 52263 38371
rect 50222 38355 52266 38367
rect 50222 38303 52195 38355
rect 50222 38236 50336 38303
rect 52191 38291 52195 38303
rect 52259 38303 52266 38355
rect 52259 38291 52263 38303
rect 52191 38257 52263 38291
rect 49873 38234 50336 38236
rect 38870 38095 38936 38096
rect 38870 38031 38871 38095
rect 38935 38031 39362 38095
rect 38870 38030 38936 38031
rect 31644 37877 32356 37896
rect 31574 37861 32356 37877
rect 31574 37797 31580 37861
rect 31644 37797 32356 37861
rect 31574 37781 32356 37797
rect 31574 37768 31580 37781
rect 31575 37717 31580 37768
rect 31644 37768 32356 37781
rect 31644 37717 31649 37768
rect 31575 37711 31649 37717
rect 40970 37647 41990 37711
rect 37081 36302 37145 37322
rect 45839 36295 45903 37315
rect 38372 35017 39392 35081
rect 40972 35017 41992 35081
rect 43572 35017 44592 35081
rect 49873 34932 50336 34934
rect 49873 34696 49986 34932
rect 50222 34854 50336 34932
rect 50931 34854 51158 34856
rect 50222 34849 51165 34854
rect 50222 34790 50932 34849
rect 50222 34696 50336 34790
rect 50931 34785 50932 34790
rect 50996 34785 51012 34849
rect 51076 34785 51092 34849
rect 51156 34790 51165 34849
rect 51156 34785 51158 34790
rect 50931 34779 51158 34785
rect 49873 34694 50336 34696
rect 46123 34245 46189 34246
rect 46123 34181 46124 34245
rect 46188 34181 46189 34245
rect 46123 34180 46189 34181
rect 46124 33718 46188 34180
rect 49883 33682 50346 33684
rect 49883 33446 49996 33682
rect 50232 33594 50346 33682
rect 50926 33606 51166 33615
rect 50926 33594 50934 33606
rect 50232 33542 50934 33594
rect 50998 33542 51014 33606
rect 51078 33542 51094 33606
rect 51158 33594 51166 33606
rect 51158 33542 51185 33594
rect 50232 33530 51185 33542
rect 50232 33446 50346 33530
rect 49883 33444 50346 33446
rect 38375 33367 39395 33431
rect 40975 33367 41995 33431
rect 43575 33367 44595 33431
rect 37081 31102 37145 32122
rect 40312 31629 40442 31662
rect 40312 31565 40345 31629
rect 40409 31565 40442 31629
rect 40312 31532 40442 31565
rect 40313 31062 40441 31532
rect 45839 31095 45903 32115
rect 49879 31263 50344 31266
rect 49879 31257 49993 31263
rect 50229 31257 50344 31263
rect 49879 31033 49919 31257
rect 50303 31033 50344 31257
rect 49879 31027 49993 31033
rect 50229 31027 50344 31033
rect 49879 31024 50344 31027
rect 29855 30730 30385 30732
rect 29855 30494 30002 30730
rect 30238 30668 30385 30730
rect 31572 30672 31649 30692
rect 31572 30668 31578 30672
rect 30238 30608 31578 30668
rect 31642 30668 31649 30672
rect 31642 30608 31690 30668
rect 30238 30592 31690 30608
rect 30238 30540 31578 30592
rect 30238 30494 30385 30540
rect 29855 30492 30385 30494
rect 31572 30528 31578 30540
rect 31642 30540 31690 30592
rect 31642 30528 31649 30540
rect 31572 30512 31649 30528
rect 31572 30448 31578 30512
rect 31642 30448 31649 30512
rect 31572 30429 31649 30448
rect 38842 30325 38908 30326
rect 38842 30261 38843 30325
rect 38907 30261 39394 30325
rect 38842 30260 38908 30261
rect 31571 30185 31648 30197
rect 31571 30121 31577 30185
rect 31641 30163 31648 30185
rect 52183 30186 52247 30198
rect 31641 30121 31706 30163
rect 31571 30105 31706 30121
rect 31571 30041 31577 30105
rect 31641 30041 31706 30105
rect 31571 30025 31706 30041
rect 31571 29961 31577 30025
rect 31641 29961 31706 30025
rect 31571 29950 31706 29961
rect 31578 29006 31706 29950
rect 52183 30150 52254 30186
rect 52183 30086 52188 30150
rect 52252 30086 52254 30150
rect 52183 30070 52254 30086
rect 52183 30006 52188 30070
rect 52252 30006 52254 30070
rect 53166 30065 53230 39411
rect 53585 38667 53649 40162
rect 53960 39021 54024 39023
rect 53949 38992 54034 39021
rect 53949 38928 53959 38992
rect 54023 38928 54034 38992
rect 53949 38912 54034 38928
rect 53949 38848 53959 38912
rect 54023 38848 54034 38912
rect 53949 38832 54034 38848
rect 53949 38768 53959 38832
rect 54023 38768 54034 38832
rect 53949 38740 54034 38768
rect 53584 38666 53650 38667
rect 53584 38602 53585 38666
rect 53649 38602 53650 38666
rect 53584 38601 53650 38602
rect 52183 29971 52254 30006
rect 53165 30064 53231 30065
rect 53165 30000 53166 30064
rect 53230 30000 53231 30064
rect 53165 29999 53231 30000
rect 53166 29995 53230 29999
rect 40970 29847 41990 29911
rect 49883 29784 50346 29786
rect 49883 29548 49996 29784
rect 50232 29692 50346 29784
rect 52183 29692 52247 29971
rect 50232 29628 52247 29692
rect 50232 29548 50346 29628
rect 49883 29546 50346 29548
rect 33862 29064 34392 29066
rect 33862 29006 34009 29064
rect 31578 28878 34009 29006
rect 33862 28828 34009 28878
rect 34245 28828 34392 29064
rect 33862 28826 34392 28828
rect 37081 28502 37145 29522
rect 45839 28495 45903 29515
rect 53585 29256 53649 38601
rect 53960 38070 54024 38740
rect 53895 38068 54358 38070
rect 53895 37832 54008 38068
rect 54244 37964 54358 38068
rect 54244 37900 54789 37964
rect 54244 37832 54358 37900
rect 53895 37830 54358 37832
rect 54725 36977 54789 37900
rect 55285 37143 55370 37156
rect 55285 37079 55295 37143
rect 55359 37079 55370 37143
rect 55285 37063 55370 37079
rect 55285 36999 55295 37063
rect 55359 36999 55370 37063
rect 55285 36983 55370 36999
rect 55285 36977 55295 36983
rect 54725 36919 55295 36977
rect 55359 36919 55370 36983
rect 54725 36913 55370 36919
rect 54725 35412 54789 36913
rect 55285 36903 55370 36913
rect 55285 36839 55295 36903
rect 55359 36839 55370 36903
rect 55285 36823 55370 36839
rect 55285 36759 55295 36823
rect 55359 36759 55370 36823
rect 55285 36747 55370 36759
rect 55334 35548 55402 35552
rect 55334 35484 55336 35548
rect 55400 35484 55402 35548
rect 55334 35468 55402 35484
rect 55334 35412 55336 35468
rect 54725 35404 55336 35412
rect 55400 35404 55402 35468
rect 54725 35388 55402 35404
rect 54725 35348 55336 35388
rect 55334 35324 55336 35348
rect 55400 35324 55402 35388
rect 55334 35308 55402 35324
rect 55334 35244 55336 35308
rect 55400 35244 55402 35308
rect 55334 35228 55402 35244
rect 55334 35164 55336 35228
rect 55400 35164 55402 35228
rect 55334 35161 55402 35164
rect 55334 33945 55400 33953
rect 55334 33881 55335 33945
rect 55399 33881 55400 33945
rect 55334 33865 55400 33881
rect 55334 33801 55335 33865
rect 55399 33801 55400 33865
rect 55334 33797 55400 33801
rect 54704 33785 55400 33797
rect 54704 33733 55335 33785
rect 53893 32822 54356 32824
rect 53893 32729 54006 32822
rect 53893 32665 53909 32729
rect 53973 32665 54006 32729
rect 53893 32586 54006 32665
rect 54242 32732 54356 32822
rect 54704 32732 54768 33733
rect 55334 33721 55335 33733
rect 55399 33721 55400 33785
rect 55334 33705 55400 33721
rect 55334 33641 55335 33705
rect 55399 33641 55400 33705
rect 55334 33625 55400 33641
rect 55334 33561 55335 33625
rect 55399 33561 55400 33625
rect 55334 33553 55400 33561
rect 54242 32668 54768 32732
rect 54242 32586 54356 32668
rect 53893 32584 54356 32586
rect 54704 32201 54768 32668
rect 55335 32344 55405 32353
rect 55335 32280 55338 32344
rect 55402 32280 55405 32344
rect 55335 32264 55405 32280
rect 55335 32201 55338 32264
rect 54704 32200 55338 32201
rect 55402 32200 55405 32264
rect 54704 32184 55405 32200
rect 54704 32137 55338 32184
rect 55335 32120 55338 32137
rect 55402 32120 55405 32184
rect 55335 32104 55405 32120
rect 55335 32040 55338 32104
rect 55402 32040 55405 32104
rect 55335 32024 55405 32040
rect 55335 31960 55338 32024
rect 55402 31960 55405 32024
rect 55335 31951 55405 31960
rect 53895 30763 54358 30765
rect 53895 30671 54008 30763
rect 53895 30607 53910 30671
rect 53974 30607 54008 30671
rect 53895 30527 54008 30607
rect 54244 30673 54358 30763
rect 54244 30609 54759 30673
rect 54244 30527 54358 30609
rect 53895 30525 54358 30527
rect 53900 29570 53985 29600
rect 53900 29506 53910 29570
rect 53974 29506 53985 29570
rect 53900 29490 53985 29506
rect 53900 29433 53910 29490
rect 53893 29426 53910 29433
rect 53974 29433 53985 29490
rect 54695 29433 54759 30609
rect 53974 29426 54759 29433
rect 53893 29410 54759 29426
rect 53893 29369 53910 29410
rect 53900 29346 53910 29369
rect 53974 29369 54759 29410
rect 53974 29346 53985 29369
rect 53900 29317 53985 29346
rect 53584 29255 53650 29256
rect 53584 29191 53585 29255
rect 53649 29191 53650 29255
rect 53584 29190 53650 29191
rect 38372 27217 39392 27281
rect 40972 27217 41992 27281
rect 43572 27217 44592 27281
rect 55590 20962 55654 42867
rect 65373 42740 65439 42741
rect 65373 42676 65374 42740
rect 65438 42676 65439 42740
rect 65373 42675 65439 42676
rect 55960 42673 56026 42674
rect 55960 42609 55961 42673
rect 56025 42609 56026 42673
rect 55960 42608 56026 42609
rect 55961 21319 56025 42608
rect 56413 42334 56479 42335
rect 56413 42270 56414 42334
rect 56478 42270 56479 42334
rect 56413 42269 56479 42270
rect 56414 21734 56478 42269
rect 56809 42053 56875 42054
rect 56809 41989 56810 42053
rect 56874 41989 56875 42053
rect 56809 41988 56875 41989
rect 56810 22160 56874 41988
rect 57883 41638 58346 41640
rect 57883 41402 57996 41638
rect 58232 41402 58346 41638
rect 57883 41400 58346 41402
rect 61388 41311 61454 41312
rect 63320 41311 63386 41312
rect 65374 41311 65438 42675
rect 65883 41423 66346 41425
rect 65883 41311 65996 41423
rect 61388 41247 61389 41311
rect 61453 41247 63321 41311
rect 63385 41247 65996 41311
rect 61388 41246 61454 41247
rect 63320 41246 63386 41247
rect 65883 41187 65996 41247
rect 66232 41311 66346 41423
rect 67326 41311 67390 43015
rect 66232 41247 67390 41311
rect 66232 41187 66346 41247
rect 65883 41185 66346 41187
rect 61888 40615 62350 40768
rect 61888 40469 62001 40615
rect 57344 40436 62001 40469
rect 62237 40469 62350 40615
rect 62237 40436 68234 40469
rect 57344 40292 57357 40436
rect 68221 40292 68234 40436
rect 57344 40259 62001 40292
rect 61886 40212 62001 40259
rect 61888 40059 62001 40212
rect 62237 40259 68234 40292
rect 62237 40059 62350 40259
rect 61888 39906 62350 40059
rect 69166 36385 69230 45612
rect 69682 37193 69746 47167
rect 69955 45116 70197 45119
rect 69955 44880 69958 45116
rect 70194 44880 70197 45116
rect 69955 44877 70197 44880
rect 69943 42815 70185 42818
rect 69943 42579 69946 42815
rect 70182 42579 70185 42815
rect 69943 42576 70185 42579
rect 70360 41785 70424 49555
rect 70944 42593 71008 49966
rect 72324 48871 72388 61267
rect 76976 60751 77040 65339
rect 78607 64135 78671 69683
rect 79149 69681 79150 69745
rect 79214 69681 79215 69745
rect 79149 69680 79215 69681
rect 78606 64134 78672 64135
rect 78606 64070 78607 64134
rect 78671 64070 78672 64134
rect 78606 64069 78672 64070
rect 73083 60750 73149 60751
rect 73083 60686 73084 60750
rect 73148 60686 73149 60750
rect 73083 60685 73149 60686
rect 76975 60750 77041 60751
rect 76975 60686 76976 60750
rect 77040 60686 77041 60750
rect 76975 60685 77041 60686
rect 72323 48870 72389 48871
rect 72323 48806 72324 48870
rect 72388 48806 72389 48870
rect 72323 48805 72389 48806
rect 73084 48553 73148 60685
rect 73814 60072 73880 60073
rect 73814 60008 73815 60072
rect 73879 60008 73880 60072
rect 73814 60007 73880 60008
rect 73815 53775 73879 60007
rect 74505 59365 74571 59366
rect 74505 59301 74506 59365
rect 74570 59301 74571 59365
rect 74505 59300 74571 59301
rect 73814 53774 73880 53775
rect 73814 53710 73815 53774
rect 73879 53710 73880 53774
rect 73814 53709 73880 53710
rect 74506 53352 74570 59300
rect 75345 58605 75411 58606
rect 75345 58541 75346 58605
rect 75410 58541 75411 58605
rect 75345 58540 75411 58541
rect 74505 53351 74571 53352
rect 74505 53287 74506 53351
rect 74570 53287 74571 53351
rect 74505 53286 74571 53287
rect 74506 53283 74570 53286
rect 73083 48552 73149 48553
rect 73083 48488 73084 48552
rect 73148 48488 73149 48552
rect 73083 48487 73149 48488
rect 75346 47541 75410 58540
rect 78607 57769 78671 64069
rect 79151 63764 79215 69680
rect 79691 69744 79757 69745
rect 79691 69680 79692 69744
rect 79756 69680 79757 69744
rect 80238 69685 80239 69749
rect 80303 69685 80304 69749
rect 82956 69696 82957 69760
rect 83021 69696 83022 69760
rect 83499 69700 83500 69764
rect 83564 69700 83565 69764
rect 86222 69760 86288 69761
rect 83499 69699 83565 69700
rect 84041 69758 84107 69759
rect 82956 69695 83022 69696
rect 80238 69684 80304 69685
rect 79691 69679 79757 69680
rect 79692 67945 79756 69679
rect 79690 67944 79756 67945
rect 79690 67880 79691 67944
rect 79755 67880 79756 67944
rect 79690 67879 79756 67880
rect 79150 63763 79216 63764
rect 79150 63699 79151 63763
rect 79215 63699 79216 63763
rect 79150 63698 79216 63699
rect 79151 58606 79215 63698
rect 79692 59366 79756 67879
rect 80239 67574 80303 69684
rect 82957 68914 83021 69695
rect 82956 68913 83022 68914
rect 82956 68849 82957 68913
rect 83021 68849 83022 68913
rect 82956 68848 83022 68849
rect 80238 67573 80304 67574
rect 80238 67509 80239 67573
rect 80303 67509 80304 67573
rect 80238 67508 80304 67509
rect 80239 60073 80303 67508
rect 82957 62441 83021 68848
rect 83500 68549 83564 69699
rect 84041 69694 84042 69758
rect 84106 69694 84107 69758
rect 84041 69693 84107 69694
rect 84598 69749 84664 69750
rect 83499 68548 83565 68549
rect 83499 68484 83500 68548
rect 83564 68484 83565 68548
rect 83499 68483 83565 68484
rect 82956 62440 83022 62441
rect 82956 62376 82957 62440
rect 83021 62376 83022 62440
rect 82956 62375 83022 62376
rect 83500 61861 83564 68483
rect 84042 65224 84106 69693
rect 84598 69685 84599 69749
rect 84663 69685 84664 69749
rect 86222 69696 86223 69760
rect 86287 69696 86288 69760
rect 87316 69757 87382 69758
rect 86222 69695 86288 69696
rect 86766 69753 86832 69754
rect 84598 69684 84664 69685
rect 84041 65223 84107 65224
rect 84041 65159 84042 65223
rect 84106 65159 84107 65223
rect 84041 65158 84107 65159
rect 83499 61860 83565 61861
rect 83499 61796 83500 61860
rect 83564 61796 83565 61860
rect 83499 61795 83565 61796
rect 80238 60072 80304 60073
rect 80238 60008 80239 60072
rect 80303 60008 80304 60072
rect 80238 60007 80304 60008
rect 79691 59365 79757 59366
rect 79691 59301 79692 59365
rect 79756 59301 79757 59365
rect 79691 59300 79757 59301
rect 79692 59280 79756 59300
rect 79149 58605 79215 58606
rect 79149 58541 79150 58605
rect 79214 58541 79215 58605
rect 84042 58545 84106 65158
rect 84599 64859 84663 69684
rect 84598 64858 84664 64859
rect 84598 64794 84599 64858
rect 84663 64794 84664 64858
rect 84598 64793 84664 64794
rect 79149 58540 79215 58541
rect 84041 58544 84107 58545
rect 84041 58480 84042 58544
rect 84106 58480 84107 58544
rect 84041 58479 84107 58480
rect 84599 57836 84663 64793
rect 86223 63589 86287 69695
rect 86766 69689 86767 69753
rect 86831 69689 86832 69753
rect 86766 69688 86832 69689
rect 87316 69693 87317 69757
rect 87381 69693 87382 69757
rect 87316 69692 87382 69693
rect 87849 69757 87915 69758
rect 87849 69693 87850 69757
rect 87914 69693 87915 69757
rect 87849 69692 87915 69693
rect 86767 63954 86831 69688
rect 87316 67398 87380 69692
rect 87850 67764 87914 69692
rect 87849 67763 87915 67764
rect 87849 67699 87850 67763
rect 87914 67699 87915 67763
rect 87849 67698 87915 67699
rect 87315 67397 87381 67398
rect 87315 67333 87316 67397
rect 87380 67333 87381 67397
rect 87315 67332 87381 67333
rect 86766 63953 86832 63954
rect 86766 63889 86767 63953
rect 86831 63889 86832 63953
rect 86766 63888 86832 63889
rect 86222 63588 86288 63589
rect 86222 63524 86223 63588
rect 86287 63524 86288 63588
rect 86222 63523 86288 63524
rect 86223 59281 86287 63523
rect 86767 59993 86831 63888
rect 87316 60616 87380 67332
rect 87850 61252 87914 67698
rect 89507 62440 89573 62441
rect 89507 62376 89508 62440
rect 89572 62376 89573 62440
rect 89507 62375 89573 62376
rect 88917 61860 88983 61861
rect 88917 61796 88918 61860
rect 88982 61796 88983 61860
rect 88917 61795 88983 61796
rect 87849 61251 87915 61252
rect 87849 61187 87850 61251
rect 87914 61187 87915 61251
rect 87849 61186 87915 61187
rect 88324 61251 88390 61252
rect 88324 61187 88325 61251
rect 88389 61187 88390 61251
rect 88324 61186 88390 61187
rect 87315 60615 87381 60616
rect 87315 60551 87316 60615
rect 87380 60551 87381 60615
rect 87315 60550 87381 60551
rect 87677 60615 87743 60616
rect 87677 60551 87678 60615
rect 87742 60551 87743 60615
rect 87677 60550 87743 60551
rect 86766 59992 86832 59993
rect 86766 59928 86767 59992
rect 86831 59928 86832 59992
rect 86766 59927 86832 59928
rect 87083 59992 87149 59993
rect 87083 59928 87084 59992
rect 87148 59928 87149 59992
rect 87083 59927 87149 59928
rect 86222 59280 86288 59281
rect 86222 59216 86223 59280
rect 86287 59216 86288 59280
rect 86222 59215 86288 59216
rect 86500 59280 86566 59281
rect 86500 59216 86501 59280
rect 86565 59216 86566 59280
rect 86500 59215 86566 59216
rect 85921 58544 85987 58545
rect 85921 58480 85922 58544
rect 85986 58480 85987 58544
rect 85921 58479 85987 58480
rect 84598 57835 84664 57836
rect 84598 57771 84599 57835
rect 84663 57771 84664 57835
rect 84598 57770 84664 57771
rect 85408 57835 85474 57836
rect 85408 57771 85409 57835
rect 85473 57771 85474 57835
rect 85408 57770 85474 57771
rect 76348 57768 76414 57769
rect 76348 57704 76349 57768
rect 76413 57704 76414 57768
rect 76348 57703 76414 57704
rect 78606 57768 78673 57769
rect 78606 57704 78607 57768
rect 78671 57704 78673 57768
rect 78606 57703 78673 57704
rect 76349 47910 76413 57703
rect 82972 50031 83038 50032
rect 82972 49967 82973 50031
rect 83037 49967 83038 50031
rect 82972 49966 83038 49967
rect 76348 47909 76414 47910
rect 76348 47845 76349 47909
rect 76413 47845 76414 47909
rect 76348 47844 76414 47845
rect 75345 47540 75411 47541
rect 75345 47476 75346 47540
rect 75410 47476 75411 47540
rect 75345 47475 75411 47476
rect 80782 43404 80848 43405
rect 71780 43350 71844 43354
rect 71780 43349 71846 43350
rect 71780 43285 71781 43349
rect 71845 43285 71846 43349
rect 80782 43340 80783 43404
rect 80847 43340 80848 43404
rect 80782 43339 80848 43340
rect 71780 43284 71846 43285
rect 71780 43117 71844 43284
rect 73983 43207 74225 43210
rect 71780 43116 71847 43117
rect 73983 43116 73986 43207
rect 71780 43052 73986 43116
rect 71208 42593 71274 42594
rect 70944 42529 71209 42593
rect 71273 42529 71274 42593
rect 71208 42528 71274 42529
rect 71461 41785 71527 41786
rect 70360 41721 71462 41785
rect 71526 41721 71527 41785
rect 71461 41720 71527 41721
rect 71783 41565 71847 43052
rect 73983 42971 73986 43052
rect 74222 42971 74225 43207
rect 73983 42968 74225 42971
rect 77987 43180 78229 43183
rect 77987 42944 77990 43180
rect 78226 42944 78229 43180
rect 77987 42941 78229 42944
rect 80783 43105 80847 43339
rect 81997 43175 82239 43178
rect 81997 43105 82000 43175
rect 80783 43041 82000 43105
rect 80783 41575 80847 43041
rect 81997 42939 82000 43041
rect 82236 42939 82239 43175
rect 81997 42936 82239 42939
rect 82707 42593 82773 42594
rect 82973 42593 83037 49966
rect 83556 49620 83622 49621
rect 83556 49556 83557 49620
rect 83621 49556 83622 49620
rect 83556 49555 83622 49556
rect 82707 42529 82708 42593
rect 82772 42529 83037 42593
rect 82707 42528 82773 42529
rect 82454 41786 82520 41787
rect 83557 41786 83621 49555
rect 84205 47233 84269 47244
rect 84204 47232 84270 47233
rect 84204 47168 84205 47232
rect 84269 47168 84270 47232
rect 84204 47167 84270 47168
rect 82454 41722 82455 41786
rect 82519 41722 83621 41786
rect 82454 41721 82520 41722
rect 80782 41574 80848 41575
rect 71782 41564 71848 41565
rect 71782 41500 71783 41564
rect 71847 41500 71848 41564
rect 80782 41510 80783 41574
rect 80847 41510 80848 41574
rect 80782 41509 80848 41510
rect 71782 41499 71848 41500
rect 69937 41210 70179 41213
rect 69937 40974 69940 41210
rect 70176 40974 70179 41210
rect 69937 40971 70179 40974
rect 80779 39810 80845 39811
rect 71779 39756 71918 39791
rect 71758 39733 71918 39756
rect 80779 39746 80780 39810
rect 80844 39746 80845 39810
rect 80779 39745 80845 39746
rect 71758 39669 71780 39733
rect 71844 39669 71918 39733
rect 71758 39647 71918 39669
rect 71779 39546 71918 39647
rect 73891 39614 74133 39617
rect 73891 39546 73894 39614
rect 71779 39445 73894 39546
rect 69956 39339 70198 39342
rect 69956 39103 69959 39339
rect 70195 39103 70198 39339
rect 69956 39100 70198 39103
rect 71779 37988 71918 39445
rect 73891 39378 73894 39445
rect 74130 39378 74133 39614
rect 73891 39375 74133 39378
rect 77930 39609 78172 39612
rect 77930 39373 77933 39609
rect 78169 39373 78172 39609
rect 77930 39370 78172 39373
rect 80780 39495 80844 39745
rect 81999 39582 82241 39585
rect 81999 39495 82002 39582
rect 80780 39431 82002 39495
rect 80780 38020 80844 39431
rect 81999 39346 82002 39431
rect 82238 39346 82241 39582
rect 81999 39343 82241 39346
rect 71778 37987 71918 37988
rect 71778 37923 71779 37987
rect 71843 37923 71918 37987
rect 80779 38019 80845 38020
rect 80779 37955 80780 38019
rect 80844 37955 80845 38019
rect 80779 37954 80845 37955
rect 71778 37922 71918 37923
rect 69978 37638 70220 37641
rect 69978 37402 69981 37638
rect 70217 37402 70220 37638
rect 69978 37399 70220 37402
rect 71208 37193 71274 37194
rect 69682 37129 71209 37193
rect 71273 37129 71274 37193
rect 71208 37128 71274 37129
rect 71461 36385 71527 36386
rect 69166 36321 71462 36385
rect 71526 36321 71527 36385
rect 71461 36320 71527 36321
rect 71779 36202 71918 37922
rect 84205 37193 84269 47167
rect 84751 45678 84815 45687
rect 84750 45677 84816 45678
rect 84750 45613 84751 45677
rect 84815 45613 84816 45677
rect 84750 45612 84816 45613
rect 82772 37129 84269 37193
rect 84751 36386 84815 45612
rect 82519 36322 84815 36386
rect 71779 36138 71796 36202
rect 71860 36138 71918 36202
rect 80784 36212 80850 36213
rect 80784 36148 80785 36212
rect 80849 36148 80850 36212
rect 80784 36147 80850 36148
rect 69991 35783 70233 35786
rect 69991 35547 69994 35783
rect 70230 35547 70233 35783
rect 69991 35544 70233 35547
rect 69877 34673 70340 34675
rect 69877 34639 69990 34673
rect 67898 34560 69990 34639
rect 63576 34540 69990 34560
rect 63576 34396 63592 34540
rect 68296 34461 69990 34540
rect 68296 34396 68432 34461
rect 69877 34437 69990 34461
rect 70226 34639 70340 34673
rect 70226 34461 70383 34639
rect 70226 34437 70340 34461
rect 69877 34435 70340 34437
rect 63576 34377 68432 34396
rect 67898 34348 68432 34377
rect 71779 34405 71918 36138
rect 77984 36021 78226 36024
rect 77984 35785 77987 36021
rect 78223 35785 78226 36021
rect 77984 35782 78226 35785
rect 80785 35912 80849 36147
rect 81987 35991 82229 35994
rect 81987 35912 81990 35991
rect 80785 35848 81990 35912
rect 71779 34372 71785 34405
rect 71784 34341 71785 34372
rect 71849 34372 71918 34405
rect 80785 34403 80849 35848
rect 81987 35755 81990 35848
rect 82226 35755 82229 35991
rect 81987 35752 82229 35755
rect 80784 34402 80850 34403
rect 71849 34341 71850 34372
rect 71784 34340 71850 34341
rect 80784 34338 80785 34402
rect 80849 34338 80850 34402
rect 80784 34337 80850 34338
rect 65908 24357 66371 24359
rect 57888 24345 58351 24347
rect 57888 24255 58001 24345
rect 57415 24243 58001 24255
rect 58237 24255 58351 24345
rect 61697 24255 62011 24312
rect 65908 24255 66021 24357
rect 58237 24243 66021 24255
rect 66257 24255 66371 24357
rect 69263 24255 69514 24356
rect 73885 24345 74348 24347
rect 73885 24255 73998 24345
rect 66257 24243 73998 24255
rect 74234 24255 74348 24345
rect 74234 24243 78202 24255
rect 57415 24099 57416 24243
rect 78200 24099 78202 24243
rect 57415 24088 78202 24099
rect 85409 22160 85473 57770
rect 56810 22096 85473 22160
rect 85922 21734 85986 58479
rect 56414 21670 85986 21734
rect 86501 21319 86565 59215
rect 55961 21255 86565 21319
rect 87084 20962 87148 59927
rect 55590 20898 87148 20962
rect 78295 20513 78361 20514
rect 87678 20513 87742 60550
rect 78295 20449 78296 20513
rect 78360 20449 87742 20513
rect 78295 20448 78361 20449
rect 78295 20041 78361 20042
rect 88325 20041 88389 61186
rect 78295 19977 78296 20041
rect 78360 19977 88389 20041
rect 78295 19976 78361 19977
rect 78295 19506 78361 19507
rect 88918 19506 88982 61795
rect 78295 19442 78296 19506
rect 78360 19442 88982 19506
rect 78295 19441 78361 19442
rect 78295 19043 78361 19044
rect 89508 19043 89572 62375
rect 89885 48154 90348 48156
rect 89885 47918 89998 48154
rect 90234 48070 90348 48154
rect 90234 48006 92310 48070
rect 90234 47918 90348 48006
rect 89885 47916 90348 47918
rect 92246 47889 92310 48006
rect 92245 47888 92311 47889
rect 92245 47824 92246 47888
rect 92310 47824 92311 47888
rect 92245 47823 92311 47824
rect 89884 45694 90347 45696
rect 89884 45458 89997 45694
rect 90233 45607 90347 45694
rect 92245 45607 92311 45608
rect 90233 45543 92246 45607
rect 92310 45543 92311 45607
rect 90233 45458 90347 45543
rect 92245 45542 92311 45543
rect 89884 45456 90347 45458
rect 92571 45402 92635 92037
rect 93160 48041 93224 92660
rect 93159 48040 93225 48041
rect 93159 47976 93160 48040
rect 93224 47976 93225 48040
rect 93159 47975 93225 47976
rect 92570 45401 92636 45402
rect 92570 45337 92571 45401
rect 92635 45337 92636 45401
rect 92570 45336 92636 45337
rect 92571 32554 92635 45336
rect 93160 33177 93224 47975
rect 93159 33176 93225 33177
rect 93159 33112 93160 33176
rect 93224 33112 93225 33176
rect 93159 33111 93225 33112
rect 92571 32553 92648 32554
rect 92571 32489 92583 32553
rect 92647 32489 92648 32553
rect 92571 32488 92648 32489
rect 89887 31313 90350 31315
rect 89887 31077 90000 31313
rect 90236 31245 90350 31313
rect 92121 31245 92187 31246
rect 90236 31181 92122 31245
rect 92186 31181 92187 31245
rect 90236 31077 90350 31181
rect 92121 31180 92187 31181
rect 89887 31075 90350 31077
rect 89878 30013 90341 30015
rect 89878 29777 89991 30013
rect 90227 29907 90341 30013
rect 92120 29907 92186 29908
rect 90227 29843 92121 29907
rect 92185 29843 92186 29907
rect 90227 29777 90341 29843
rect 92120 29842 92186 29843
rect 89878 29775 90341 29777
rect 89884 28598 90347 28600
rect 89884 28362 89997 28598
rect 90233 28514 90347 28598
rect 92128 28514 92194 28515
rect 90233 28450 92129 28514
rect 92193 28450 92194 28514
rect 90233 28362 90347 28450
rect 92128 28449 92194 28450
rect 89884 28360 90347 28362
rect 89880 27225 90343 27227
rect 89880 26989 89993 27225
rect 90229 27144 90343 27225
rect 92124 27144 92190 27145
rect 90229 27080 92125 27144
rect 92189 27080 92190 27144
rect 90229 26989 90343 27080
rect 92124 27079 92190 27080
rect 89880 26987 90343 26989
rect 92571 25614 92635 32488
rect 93160 26237 93224 33111
rect 93725 32492 93789 93280
rect 101830 69194 102418 69201
rect 101830 69094 102002 69194
rect 102238 69094 102418 69194
rect 101830 69030 101852 69094
rect 101916 69030 101932 69094
rect 101996 69030 102002 69094
rect 102238 69030 102252 69094
rect 102316 69030 102332 69094
rect 102396 69030 102418 69094
rect 101830 68958 102002 69030
rect 102238 68958 102418 69030
rect 101830 68953 102418 68958
rect 98681 68550 98921 68573
rect 98609 68548 98969 68550
rect 98609 68484 98637 68548
rect 98701 68484 98717 68548
rect 98781 68484 98797 68548
rect 98861 68484 98877 68548
rect 98941 68484 98969 68548
rect 98609 68483 98969 68484
rect 98681 68326 98921 68483
rect 97894 68324 98921 68326
rect 97894 68088 98007 68324
rect 98243 68088 98921 68324
rect 97894 68086 98921 68088
rect 98681 67400 98921 68086
rect 101889 68033 102352 68035
rect 101889 67948 102002 68033
rect 101859 67943 102002 67948
rect 102238 67948 102352 68033
rect 102238 67943 102388 67948
rect 101859 67879 101891 67943
rect 101955 67879 101971 67943
rect 102275 67879 102291 67943
rect 102355 67879 102388 67943
rect 101859 67875 102002 67879
rect 101889 67797 102002 67875
rect 102238 67875 102388 67879
rect 102238 67797 102352 67875
rect 101889 67795 102352 67797
rect 98607 67398 98967 67400
rect 98607 67334 98635 67398
rect 98699 67334 98715 67398
rect 98779 67334 98795 67398
rect 98859 67334 98875 67398
rect 98939 67334 98967 67398
rect 98607 67333 98967 67334
rect 98681 67317 98921 67333
rect 101873 65524 102336 65526
rect 101873 65406 101986 65524
rect 101849 65401 101986 65406
rect 102222 65406 102336 65524
rect 102222 65401 102378 65406
rect 101849 65337 101881 65401
rect 101945 65337 101961 65401
rect 102265 65337 102281 65401
rect 102345 65337 102378 65401
rect 101849 65333 101986 65337
rect 101873 65288 101986 65333
rect 102222 65333 102378 65337
rect 102222 65288 102336 65333
rect 101873 65286 102336 65288
rect 98588 64859 98828 64877
rect 98525 64857 98885 64859
rect 98525 64793 98553 64857
rect 98617 64793 98633 64857
rect 98697 64793 98713 64857
rect 98777 64793 98793 64857
rect 98857 64793 98885 64857
rect 98525 64792 98885 64793
rect 98588 64581 98828 64792
rect 97902 64579 98828 64581
rect 97902 64343 98015 64579
rect 98251 64343 98828 64579
rect 97902 64341 98828 64343
rect 98588 63590 98828 64341
rect 101866 64213 102329 64215
rect 101866 64136 101979 64213
rect 101849 64131 101979 64136
rect 102215 64136 102329 64213
rect 102215 64131 102378 64136
rect 101849 64067 101881 64131
rect 101945 64067 101961 64131
rect 102265 64067 102281 64131
rect 102345 64067 102378 64131
rect 101849 64063 101979 64067
rect 101866 63977 101979 64063
rect 102215 64063 102378 64067
rect 102215 63977 102329 64063
rect 101866 63975 102329 63977
rect 98523 63588 98883 63590
rect 98523 63524 98551 63588
rect 98615 63524 98631 63588
rect 98695 63524 98711 63588
rect 98775 63524 98791 63588
rect 98855 63524 98883 63588
rect 98523 63523 98883 63524
rect 98588 63505 98828 63523
rect 99879 48272 103393 48274
rect 99879 48173 102008 48272
rect 102244 48173 103393 48272
rect 99879 48109 99985 48173
rect 100049 48109 100065 48173
rect 100129 48109 100145 48173
rect 100209 48109 100225 48173
rect 100289 48109 100305 48173
rect 100369 48109 100385 48173
rect 100449 48109 100465 48173
rect 100529 48109 100545 48173
rect 100609 48109 100625 48173
rect 100689 48109 100705 48173
rect 100769 48109 100785 48173
rect 100849 48109 100865 48173
rect 100929 48109 100945 48173
rect 101009 48109 101025 48173
rect 101089 48109 101105 48173
rect 101169 48109 101185 48173
rect 101249 48109 101265 48173
rect 101329 48109 101345 48173
rect 101409 48109 101425 48173
rect 101489 48109 101505 48173
rect 101569 48109 101585 48173
rect 101649 48109 101665 48173
rect 101729 48109 101745 48173
rect 101809 48109 101825 48173
rect 101889 48109 101905 48173
rect 101969 48109 101985 48173
rect 102289 48109 102305 48173
rect 102369 48109 102385 48173
rect 102449 48109 102465 48173
rect 102529 48109 102545 48173
rect 102609 48109 102625 48173
rect 102689 48109 102705 48173
rect 102769 48109 102785 48173
rect 102849 48109 102865 48173
rect 102929 48109 102945 48173
rect 103009 48109 103025 48173
rect 103089 48109 103105 48173
rect 103169 48109 103185 48173
rect 103249 48109 103393 48173
rect 99879 48036 102008 48109
rect 102244 48036 103393 48109
rect 99879 48034 103393 48036
rect 94755 47697 97269 47750
rect 94755 47633 96445 47697
rect 96509 47633 97269 47697
rect 94755 47617 97269 47633
rect 94755 47605 96445 47617
rect 94755 47541 94917 47605
rect 94981 47553 96445 47605
rect 96509 47553 97269 47617
rect 94981 47541 97269 47553
rect 94755 47510 97269 47541
rect 94912 47212 95000 47217
rect 96428 47212 96516 47223
rect 94368 47210 96591 47212
rect 94368 47204 96440 47210
rect 94368 47140 94924 47204
rect 94988 47146 96440 47204
rect 96504 47146 96591 47210
rect 94988 47140 96591 47146
rect 94368 47130 96591 47140
rect 94368 47124 96440 47130
rect 94368 47060 94924 47124
rect 94988 47066 96440 47124
rect 96504 47066 96591 47130
rect 94988 47060 96591 47066
rect 94368 47050 96591 47060
rect 94368 47044 96440 47050
rect 94368 46980 94924 47044
rect 94988 46986 96440 47044
rect 96504 46986 96591 47050
rect 94988 46980 96591 46986
rect 94368 46976 96591 46980
rect 94368 46838 94604 46976
rect 94912 46967 95000 46976
rect 96428 46973 96516 46976
rect 94007 46837 94604 46838
rect 94007 46601 94011 46837
rect 94247 46602 94604 46837
rect 94247 46601 94251 46602
rect 94007 46600 94251 46601
rect 94368 45849 94604 46602
rect 97029 46754 97269 47510
rect 97029 46752 98358 46754
rect 97029 46516 98008 46752
rect 98244 46516 98358 46752
rect 97029 46514 98358 46516
rect 97029 46424 97269 46514
rect 94826 46371 97269 46424
rect 94826 46307 96445 46371
rect 96509 46307 97269 46371
rect 94826 46291 97269 46307
rect 94826 46269 96445 46291
rect 94826 46205 94923 46269
rect 94987 46227 96445 46269
rect 96509 46227 97269 46291
rect 94987 46205 97269 46227
rect 94826 46184 97269 46205
rect 94919 46172 94991 46184
rect 96434 45849 96522 45857
rect 94368 45844 96591 45849
rect 94368 45816 96446 45844
rect 94368 45752 94918 45816
rect 94982 45780 96446 45816
rect 96510 45780 96591 45844
rect 94982 45764 96591 45780
rect 94982 45752 96446 45764
rect 94368 45736 96446 45752
rect 94368 45672 94918 45736
rect 94982 45700 96446 45736
rect 96510 45700 96591 45764
rect 94982 45684 96591 45700
rect 94982 45672 96446 45684
rect 94368 45620 96446 45672
rect 96510 45620 96591 45684
rect 94368 45613 96591 45620
rect 96434 45607 96522 45613
rect 105885 45266 106348 45267
rect 99823 45265 106348 45266
rect 99823 45177 105998 45265
rect 99823 45113 99983 45177
rect 100047 45113 100063 45177
rect 100127 45113 100143 45177
rect 100207 45113 100223 45177
rect 100287 45113 100303 45177
rect 100367 45113 100383 45177
rect 100447 45113 100463 45177
rect 100527 45113 100543 45177
rect 100607 45113 100623 45177
rect 100687 45113 100703 45177
rect 100767 45113 100783 45177
rect 100847 45113 100863 45177
rect 100927 45113 100943 45177
rect 101007 45113 101023 45177
rect 101087 45113 101103 45177
rect 101167 45113 101183 45177
rect 101247 45113 101263 45177
rect 101327 45113 101343 45177
rect 101407 45113 101423 45177
rect 101487 45113 101503 45177
rect 101567 45113 101583 45177
rect 101647 45113 101663 45177
rect 101727 45113 101743 45177
rect 101807 45113 101823 45177
rect 101887 45113 101903 45177
rect 101967 45113 101983 45177
rect 102047 45113 102063 45177
rect 102127 45113 102143 45177
rect 102207 45113 102223 45177
rect 102287 45113 102303 45177
rect 102367 45113 102383 45177
rect 102447 45113 102463 45177
rect 102527 45113 102543 45177
rect 102607 45113 102623 45177
rect 102687 45113 102703 45177
rect 102767 45113 102783 45177
rect 102847 45113 102863 45177
rect 102927 45113 102943 45177
rect 103007 45113 103023 45177
rect 103087 45113 103103 45177
rect 103167 45113 103183 45177
rect 103247 45113 105998 45177
rect 99823 45029 105998 45113
rect 106234 45029 106348 45265
rect 99823 45027 106348 45029
rect 99823 45026 106125 45027
rect 93975 32813 94249 32832
rect 93975 32577 93994 32813
rect 94230 32577 94249 32813
rect 93975 32559 94249 32577
rect 93724 32491 93790 32492
rect 93724 32427 93725 32491
rect 93789 32427 93790 32491
rect 93724 32426 93790 32427
rect 93159 26236 93225 26237
rect 93159 26172 93160 26236
rect 93224 26172 93225 26236
rect 93159 26171 93225 26172
rect 93160 26158 93224 26171
rect 92571 25613 92648 25614
rect 92571 25549 92583 25613
rect 92647 25549 92648 25613
rect 93725 25552 93789 32426
rect 94065 31372 94161 32559
rect 94989 31615 95225 32576
rect 94989 31563 95761 31615
rect 94989 31499 95670 31563
rect 95734 31499 95761 31563
rect 94989 31483 95761 31499
rect 94989 31419 95670 31483
rect 95734 31419 95761 31483
rect 94989 31379 95761 31419
rect 96496 31612 96732 32575
rect 96496 31576 97283 31612
rect 96496 31512 97189 31576
rect 97253 31512 97283 31576
rect 96496 31496 97283 31512
rect 96496 31432 97189 31496
rect 97253 31432 97283 31496
rect 94064 31355 94162 31372
rect 94064 31291 94081 31355
rect 94145 31291 94162 31355
rect 94064 31274 94162 31291
rect 94065 30547 94161 31274
rect 94989 31160 95225 31379
rect 94988 30924 95225 31160
rect 94989 30547 95225 30924
rect 96496 31376 97283 31432
rect 101890 31466 102353 31468
rect 96496 30547 96732 31376
rect 101890 31255 102003 31466
rect 99695 31241 102003 31255
rect 102239 31255 102353 31466
rect 102239 31241 103018 31255
rect 97894 31190 98359 31193
rect 97894 31184 98008 31190
rect 98244 31184 98359 31190
rect 97894 30960 97934 31184
rect 98318 30960 98359 31184
rect 99695 31177 99724 31241
rect 99788 31177 99804 31241
rect 99868 31177 99884 31241
rect 99948 31177 99964 31241
rect 100028 31177 100044 31241
rect 100108 31177 100124 31241
rect 100188 31177 100204 31241
rect 100268 31177 100284 31241
rect 100348 31177 100364 31241
rect 100428 31177 100444 31241
rect 100508 31177 100524 31241
rect 100588 31177 100604 31241
rect 100668 31177 100684 31241
rect 100748 31177 100764 31241
rect 100828 31177 100844 31241
rect 100908 31177 100924 31241
rect 100988 31177 101004 31241
rect 101068 31177 101084 31241
rect 101148 31177 101164 31241
rect 101228 31177 101244 31241
rect 101308 31177 101324 31241
rect 101388 31177 101404 31241
rect 101468 31177 101484 31241
rect 101548 31177 101564 31241
rect 101628 31177 101644 31241
rect 101708 31177 101724 31241
rect 101788 31177 101804 31241
rect 101868 31177 101884 31241
rect 101948 31177 101964 31241
rect 102028 31177 102044 31230
rect 102108 31177 102124 31230
rect 102188 31177 102204 31230
rect 102268 31177 102284 31241
rect 102348 31177 102364 31241
rect 102428 31177 102444 31241
rect 102508 31177 102524 31241
rect 102588 31177 102604 31241
rect 102668 31177 102684 31241
rect 102748 31177 102764 31241
rect 102828 31177 102844 31241
rect 102908 31177 102924 31241
rect 102988 31177 103018 31241
rect 99695 31164 103018 31177
rect 97894 30954 98008 30960
rect 98244 30954 98359 30960
rect 97894 30951 98359 30954
rect 94032 30311 94035 30547
rect 94271 30311 96732 30547
rect 94064 30271 94162 30311
rect 94064 30207 94081 30271
rect 94145 30207 94162 30271
rect 94064 30190 94162 30207
rect 94065 29200 94161 30190
rect 94064 29183 94162 29200
rect 94064 29131 94081 29183
rect 94145 29131 94162 29183
rect 94989 29131 95225 30311
rect 95656 30232 95740 30311
rect 95656 30168 95665 30232
rect 95729 30227 95740 30232
rect 96496 30297 96732 30311
rect 96496 30229 97269 30297
rect 95729 30168 95739 30227
rect 95656 30152 95739 30168
rect 95656 30088 95665 30152
rect 95729 30088 95739 30152
rect 95656 30065 95739 30088
rect 96496 30165 97194 30229
rect 97258 30165 97269 30229
rect 96496 30149 97269 30165
rect 96496 30085 97194 30149
rect 97258 30085 97269 30149
rect 96496 30061 97269 30085
rect 96496 29131 96732 30061
rect 93993 28895 93996 29131
rect 94232 28895 96732 29131
rect 94065 28112 94161 28895
rect 94065 28095 94163 28112
rect 94065 28031 94082 28095
rect 94146 28031 94163 28095
rect 94065 28014 94163 28031
rect 94065 26854 94161 28014
rect 94989 27522 95225 28895
rect 95655 28879 95738 28895
rect 95655 28815 95664 28879
rect 95728 28815 95738 28879
rect 95655 28799 95738 28815
rect 95655 28735 95664 28799
rect 95728 28735 95738 28799
rect 95655 28712 95738 28735
rect 96496 28857 97283 28895
rect 96496 28793 97194 28857
rect 97258 28793 97283 28857
rect 96496 28777 97283 28793
rect 96496 28713 97194 28777
rect 97258 28713 97283 28777
rect 96496 28659 97283 28713
rect 96496 27525 96732 28659
rect 97892 28289 98357 28290
rect 97892 28287 103096 28289
rect 97892 28281 98006 28287
rect 98242 28281 103096 28287
rect 97892 28057 97932 28281
rect 98316 28242 103096 28281
rect 98316 28178 99701 28242
rect 99765 28178 99781 28242
rect 99845 28178 99861 28242
rect 99925 28178 99941 28242
rect 100005 28178 100021 28242
rect 100085 28178 100101 28242
rect 100165 28178 100181 28242
rect 100245 28178 100261 28242
rect 100325 28178 100341 28242
rect 100405 28178 100421 28242
rect 100485 28178 100501 28242
rect 100565 28178 100581 28242
rect 100645 28178 100661 28242
rect 100725 28178 100741 28242
rect 100805 28178 100821 28242
rect 100885 28178 100901 28242
rect 100965 28178 100981 28242
rect 101045 28178 101061 28242
rect 101125 28178 101141 28242
rect 101205 28178 101221 28242
rect 101285 28178 101301 28242
rect 101365 28178 101381 28242
rect 101445 28178 101461 28242
rect 101525 28178 101541 28242
rect 101605 28178 101621 28242
rect 101685 28178 101701 28242
rect 101765 28178 101781 28242
rect 101845 28178 101861 28242
rect 101925 28178 101941 28242
rect 102005 28178 102021 28242
rect 102085 28178 102101 28242
rect 102165 28178 102181 28242
rect 102245 28178 102261 28242
rect 102325 28178 102341 28242
rect 102405 28178 102421 28242
rect 102485 28178 102501 28242
rect 102565 28178 102581 28242
rect 102645 28178 102661 28242
rect 102725 28178 102741 28242
rect 102805 28178 102821 28242
rect 102885 28178 102901 28242
rect 102965 28178 102981 28242
rect 103045 28178 103096 28242
rect 98316 28057 103096 28178
rect 97892 28051 98006 28057
rect 98242 28051 103096 28057
rect 97892 28049 103096 28051
rect 97892 28048 98357 28049
rect 94989 27502 95740 27522
rect 94989 27479 95741 27502
rect 94989 27415 95667 27479
rect 95731 27415 95741 27479
rect 94989 27399 95741 27415
rect 94989 27335 95667 27399
rect 95731 27335 95741 27399
rect 94989 27312 95741 27335
rect 96496 27473 97281 27525
rect 96496 27409 97191 27473
rect 97255 27409 97281 27473
rect 96496 27393 97281 27409
rect 96496 27329 97191 27393
rect 97255 27329 97281 27393
rect 94989 27286 95740 27312
rect 96496 27289 97281 27329
rect 93983 26835 94257 26854
rect 93983 26599 94002 26835
rect 94238 26599 94257 26835
rect 94989 26772 95225 27286
rect 96496 26842 96732 27289
rect 93983 26581 94257 26599
rect 93975 25873 94249 25892
rect 93975 25637 93994 25873
rect 94230 25637 94249 25873
rect 93975 25619 94249 25637
rect 92571 25548 92648 25549
rect 93724 25551 93790 25552
rect 92571 25515 92635 25548
rect 93724 25487 93725 25551
rect 93789 25487 93790 25551
rect 93724 25486 93790 25487
rect 93725 25458 93789 25486
rect 94065 24432 94161 25619
rect 94989 24675 95225 25636
rect 94989 24623 95761 24675
rect 94989 24559 95670 24623
rect 95734 24559 95761 24623
rect 94989 24543 95761 24559
rect 94989 24479 95670 24543
rect 95734 24479 95761 24543
rect 94989 24439 95761 24479
rect 96496 24672 96732 25635
rect 96496 24636 97283 24672
rect 96496 24572 97189 24636
rect 97253 24572 97283 24636
rect 96496 24556 97283 24572
rect 96496 24492 97189 24556
rect 97253 24492 97283 24556
rect 94064 24415 94162 24432
rect 89887 24373 90350 24375
rect 89887 24137 90000 24373
rect 90236 24305 90350 24373
rect 94064 24351 94081 24415
rect 94145 24351 94162 24415
rect 94064 24334 94162 24351
rect 92121 24305 92187 24306
rect 90236 24241 92122 24305
rect 92186 24241 92187 24305
rect 90236 24137 90350 24241
rect 92121 24240 92187 24241
rect 89887 24135 90350 24137
rect 94065 23607 94161 24334
rect 94989 24220 95225 24439
rect 94988 23984 95225 24220
rect 94989 23607 95225 23984
rect 96496 24436 97283 24492
rect 101893 24541 102356 24543
rect 96496 23607 96732 24436
rect 101893 24332 102006 24541
rect 99692 24308 102006 24332
rect 102242 24332 102356 24541
rect 102242 24308 103025 24332
rect 97894 24250 98359 24253
rect 97894 24244 98008 24250
rect 98244 24244 98359 24250
rect 97894 24020 97934 24244
rect 98318 24020 98359 24244
rect 99692 24244 99726 24308
rect 99790 24244 99806 24308
rect 99870 24244 99886 24308
rect 99950 24244 99966 24308
rect 100030 24244 100046 24308
rect 100110 24244 100126 24308
rect 100190 24244 100206 24308
rect 100270 24244 100286 24308
rect 100350 24244 100366 24308
rect 100430 24244 100446 24308
rect 100510 24244 100526 24308
rect 100590 24244 100606 24308
rect 100670 24244 100686 24308
rect 100750 24244 100766 24308
rect 100830 24244 100846 24308
rect 100910 24244 100926 24308
rect 100990 24244 101006 24308
rect 101070 24244 101086 24308
rect 101150 24244 101166 24308
rect 101230 24244 101246 24308
rect 101310 24244 101326 24308
rect 101390 24244 101406 24308
rect 101470 24244 101486 24308
rect 101550 24244 101566 24308
rect 101630 24244 101646 24308
rect 101710 24244 101726 24308
rect 101790 24244 101806 24308
rect 101870 24244 101886 24308
rect 101950 24244 101966 24308
rect 102030 24244 102046 24305
rect 102110 24244 102126 24305
rect 102190 24244 102206 24305
rect 102270 24244 102286 24308
rect 102350 24244 102366 24308
rect 102430 24244 102446 24308
rect 102510 24244 102526 24308
rect 102590 24244 102606 24308
rect 102670 24244 102686 24308
rect 102750 24244 102766 24308
rect 102830 24244 102846 24308
rect 102910 24244 102926 24308
rect 102990 24244 103025 24308
rect 99692 24220 103025 24244
rect 97894 24014 98008 24020
rect 98244 24014 98359 24020
rect 97894 24011 98359 24014
rect 94032 23371 94035 23607
rect 94271 23371 96732 23607
rect 94064 23331 94162 23371
rect 94064 23267 94081 23331
rect 94145 23267 94162 23331
rect 94064 23250 94162 23267
rect 89878 23073 90341 23075
rect 89878 22837 89991 23073
rect 90227 22967 90341 23073
rect 92120 22967 92186 22968
rect 90227 22903 92121 22967
rect 92185 22903 92186 22967
rect 90227 22837 90341 22903
rect 92120 22902 92186 22903
rect 89878 22835 90341 22837
rect 94065 22260 94161 23250
rect 94064 22243 94162 22260
rect 94064 22191 94081 22243
rect 94145 22191 94162 22243
rect 94989 22191 95225 23371
rect 95656 23292 95740 23371
rect 95656 23228 95665 23292
rect 95729 23287 95740 23292
rect 96496 23357 96732 23371
rect 96496 23289 97269 23357
rect 95729 23228 95739 23287
rect 95656 23212 95739 23228
rect 95656 23148 95665 23212
rect 95729 23148 95739 23212
rect 95656 23125 95739 23148
rect 96496 23225 97194 23289
rect 97258 23225 97269 23289
rect 96496 23209 97269 23225
rect 96496 23145 97194 23209
rect 97258 23145 97269 23209
rect 96496 23121 97269 23145
rect 96496 22191 96732 23121
rect 93993 21955 93996 22191
rect 94232 21955 96732 22191
rect 89884 21658 90347 21660
rect 89884 21422 89997 21658
rect 90233 21574 90347 21658
rect 92128 21574 92194 21575
rect 90233 21510 92129 21574
rect 92193 21510 92194 21574
rect 90233 21422 90347 21510
rect 92128 21509 92194 21510
rect 89884 21420 90347 21422
rect 94065 21172 94161 21955
rect 94065 21155 94163 21172
rect 94065 21091 94082 21155
rect 94146 21091 94163 21155
rect 94065 21074 94163 21091
rect 89880 20285 90343 20287
rect 89880 20049 89993 20285
rect 90229 20204 90343 20285
rect 92124 20204 92190 20205
rect 90229 20140 92125 20204
rect 92189 20140 92190 20204
rect 90229 20049 90343 20140
rect 92124 20139 92190 20140
rect 89880 20047 90343 20049
rect 94065 19914 94161 21074
rect 94989 20582 95225 21955
rect 95655 21939 95738 21955
rect 95655 21875 95664 21939
rect 95728 21875 95738 21939
rect 95655 21859 95738 21875
rect 95655 21795 95664 21859
rect 95728 21795 95738 21859
rect 95655 21772 95738 21795
rect 96496 21917 97283 21955
rect 96496 21853 97194 21917
rect 97258 21853 97283 21917
rect 96496 21837 97283 21853
rect 96496 21773 97194 21837
rect 97258 21773 97283 21837
rect 96496 21719 97283 21773
rect 96496 20585 96732 21719
rect 97892 21349 98357 21350
rect 97892 21343 98611 21349
rect 97892 21342 97999 21343
rect 97879 21341 97999 21342
rect 98235 21342 98611 21343
rect 98235 21341 103157 21342
rect 97879 21117 97932 21341
rect 98316 21302 103157 21341
rect 98316 21238 99682 21302
rect 99746 21238 99762 21302
rect 99826 21238 99842 21302
rect 99906 21238 99922 21302
rect 99986 21238 100002 21302
rect 100066 21238 100082 21302
rect 100146 21238 100162 21302
rect 100226 21238 100242 21302
rect 100306 21238 100322 21302
rect 100386 21238 100402 21302
rect 100466 21238 100482 21302
rect 100546 21238 100562 21302
rect 100626 21238 100642 21302
rect 100706 21238 100722 21302
rect 100786 21238 100802 21302
rect 100866 21238 100882 21302
rect 100946 21238 100962 21302
rect 101026 21238 101042 21302
rect 101106 21238 101122 21302
rect 101186 21238 101202 21302
rect 101266 21238 101282 21302
rect 101346 21238 101362 21302
rect 101426 21238 101442 21302
rect 101506 21238 101522 21302
rect 101586 21238 101602 21302
rect 101666 21238 101682 21302
rect 101746 21238 101762 21302
rect 101826 21238 101842 21302
rect 101906 21238 101922 21302
rect 101986 21238 102002 21302
rect 102066 21238 102082 21302
rect 102146 21238 102162 21302
rect 102226 21238 102242 21302
rect 102306 21238 102322 21302
rect 102386 21238 102402 21302
rect 102466 21238 102482 21302
rect 102546 21238 102562 21302
rect 102626 21238 102642 21302
rect 102706 21238 102722 21302
rect 102786 21238 102802 21302
rect 102866 21238 102882 21302
rect 102946 21238 102962 21302
rect 103026 21238 103157 21302
rect 98316 21117 103157 21238
rect 97879 21107 97999 21117
rect 98235 21107 103157 21117
rect 97879 21102 103157 21107
rect 94989 20562 95740 20582
rect 94989 20539 95741 20562
rect 94989 20475 95667 20539
rect 95731 20475 95741 20539
rect 94989 20459 95741 20475
rect 94989 20395 95667 20459
rect 95731 20395 95741 20459
rect 94989 20372 95741 20395
rect 96496 20533 97281 20585
rect 96496 20469 97191 20533
rect 97255 20469 97281 20533
rect 96496 20453 97281 20469
rect 96496 20389 97191 20453
rect 97255 20389 97281 20453
rect 94989 20346 95740 20372
rect 96496 20349 97281 20389
rect 93983 19895 94257 19914
rect 93983 19659 94002 19895
rect 94238 19659 94257 19895
rect 94989 19832 95225 20346
rect 96496 19902 96732 20349
rect 93983 19641 94257 19659
rect 78295 18979 78296 19043
rect 78360 18979 89572 19043
rect 78295 18978 78361 18979
rect 53896 17847 56607 17849
rect 53896 17611 54009 17847
rect 54245 17611 56607 17847
rect 53896 17609 56607 17611
rect 53498 17178 53592 17201
rect 56494 17198 56607 17609
rect 53498 17114 53513 17178
rect 53577 17114 53592 17178
rect 53498 17098 53592 17114
rect 53498 17034 53513 17098
rect 53577 17034 53592 17098
rect 53498 17018 53592 17034
rect 53498 16954 53513 17018
rect 53577 16954 53592 17018
rect 53498 16938 53592 16954
rect 53498 16874 53513 16938
rect 53577 16874 53592 16938
rect 53498 16858 53592 16874
rect 53498 16794 53513 16858
rect 53577 16794 53592 16858
rect 53498 16778 53592 16794
rect 53498 16714 53513 16778
rect 53577 16714 53592 16778
rect 53498 16698 53592 16714
rect 53498 16634 53513 16698
rect 53577 16634 53592 16698
rect 53498 16618 53592 16634
rect 53498 16554 53513 16618
rect 53577 16554 53592 16618
rect 53498 16538 53592 16554
rect 53498 16474 53513 16538
rect 53577 16474 53592 16538
rect 53498 16458 53592 16474
rect 53498 16394 53513 16458
rect 53577 16394 53592 16458
rect 53498 16378 53592 16394
rect 53498 16314 53513 16378
rect 53577 16314 53592 16378
rect 53498 16298 53592 16314
rect 53498 16234 53513 16298
rect 53577 16234 53592 16298
rect 53498 16218 53592 16234
rect 53498 16154 53513 16218
rect 53577 16154 53592 16218
rect 53498 16138 53592 16154
rect 53498 16074 53513 16138
rect 53577 16074 53592 16138
rect 53498 16058 53592 16074
rect 53498 15994 53513 16058
rect 53577 15994 53592 16058
rect 53498 15978 53592 15994
rect 53498 15914 53513 15978
rect 53577 15914 53592 15978
rect 53498 15898 53592 15914
rect 53498 15834 53513 15898
rect 53577 15834 53592 15898
rect 53498 15818 53592 15834
rect 53498 15754 53513 15818
rect 53577 15754 53592 15818
rect 53498 15746 53592 15754
rect 56493 17171 56609 17198
rect 56493 17107 56519 17171
rect 56583 17107 56609 17171
rect 56493 17091 56609 17107
rect 56493 17027 56519 17091
rect 56583 17027 56609 17091
rect 56493 17011 56609 17027
rect 56493 16947 56519 17011
rect 56583 16947 56609 17011
rect 56493 16931 56609 16947
rect 56493 16867 56519 16931
rect 56583 16867 56609 16931
rect 56493 16851 56609 16867
rect 56493 16787 56519 16851
rect 56583 16787 56609 16851
rect 56493 16771 56609 16787
rect 56493 16707 56519 16771
rect 56583 16707 56609 16771
rect 56493 16691 56609 16707
rect 56493 16627 56519 16691
rect 56583 16627 56609 16691
rect 56493 16611 56609 16627
rect 56493 16547 56519 16611
rect 56583 16547 56609 16611
rect 56493 16531 56609 16547
rect 56493 16467 56519 16531
rect 56583 16467 56609 16531
rect 56493 16451 56609 16467
rect 56493 16387 56519 16451
rect 56583 16387 56609 16451
rect 56493 16371 56609 16387
rect 56493 16307 56519 16371
rect 56583 16307 56609 16371
rect 56493 16291 56609 16307
rect 56493 16227 56519 16291
rect 56583 16227 56609 16291
rect 56493 16211 56609 16227
rect 56493 16147 56519 16211
rect 56583 16147 56609 16211
rect 56493 16131 56609 16147
rect 56493 16067 56519 16131
rect 56583 16067 56609 16131
rect 56493 16051 56609 16067
rect 56493 15987 56519 16051
rect 56583 15987 56609 16051
rect 56493 15971 56609 15987
rect 56493 15907 56519 15971
rect 56583 15907 56609 15971
rect 56493 15891 56609 15907
rect 56493 15827 56519 15891
rect 56583 15827 56609 15891
rect 56493 15811 56609 15827
rect 56493 15747 56519 15811
rect 56583 15747 56609 15811
rect 49890 15744 53600 15746
rect 49890 15508 50003 15744
rect 50239 15738 53600 15744
rect 50239 15674 53513 15738
rect 53577 15674 53600 15738
rect 50239 15658 53600 15674
rect 50239 15594 53513 15658
rect 53577 15594 53600 15658
rect 50239 15578 53600 15594
rect 50239 15514 53513 15578
rect 53577 15514 53600 15578
rect 50239 15508 53600 15514
rect 49890 15506 53600 15508
rect 56493 15731 56609 15747
rect 56493 15667 56519 15731
rect 56583 15667 56609 15731
rect 56493 15651 56609 15667
rect 56493 15587 56519 15651
rect 56583 15587 56609 15651
rect 56493 15571 56609 15587
rect 56493 15507 56519 15571
rect 56583 15507 56609 15571
rect 53498 15498 53592 15506
rect 53498 15434 53513 15498
rect 53577 15434 53592 15498
rect 53498 15418 53592 15434
rect 53498 15354 53513 15418
rect 53577 15354 53592 15418
rect 53498 15338 53592 15354
rect 53498 15274 53513 15338
rect 53577 15274 53592 15338
rect 53498 15258 53592 15274
rect 53498 15194 53513 15258
rect 53577 15194 53592 15258
rect 53498 15178 53592 15194
rect 53498 15114 53513 15178
rect 53577 15114 53592 15178
rect 53498 15098 53592 15114
rect 53498 15034 53513 15098
rect 53577 15034 53592 15098
rect 53498 15018 53592 15034
rect 53498 14954 53513 15018
rect 53577 14954 53592 15018
rect 53498 14938 53592 14954
rect 53498 14874 53513 14938
rect 53577 14874 53592 14938
rect 53498 14858 53592 14874
rect 53498 14794 53513 14858
rect 53577 14794 53592 14858
rect 53498 14778 53592 14794
rect 53498 14714 53513 14778
rect 53577 14714 53592 14778
rect 53498 14698 53592 14714
rect 53498 14634 53513 14698
rect 53577 14634 53592 14698
rect 53498 14618 53592 14634
rect 53498 14554 53513 14618
rect 53577 14554 53592 14618
rect 53498 14538 53592 14554
rect 53498 14474 53513 14538
rect 53577 14474 53592 14538
rect 53498 14458 53592 14474
rect 53498 14394 53513 14458
rect 53577 14394 53592 14458
rect 53498 14378 53592 14394
rect 53498 14314 53513 14378
rect 53577 14314 53592 14378
rect 53498 14298 53592 14314
rect 53498 14234 53513 14298
rect 53577 14234 53592 14298
rect 53498 14218 53592 14234
rect 53498 14154 53513 14218
rect 53577 14154 53592 14218
rect 53498 14138 53592 14154
rect 53498 14074 53513 14138
rect 53577 14074 53592 14138
rect 53498 14058 53592 14074
rect 53498 13994 53513 14058
rect 53577 13994 53592 14058
rect 53498 13978 53592 13994
rect 53498 13914 53513 13978
rect 53577 13914 53592 13978
rect 53498 13891 53592 13914
rect 56493 15491 56609 15507
rect 56493 15427 56519 15491
rect 56583 15427 56609 15491
rect 56493 15411 56609 15427
rect 56493 15347 56519 15411
rect 56583 15347 56609 15411
rect 56493 15331 56609 15347
rect 56493 15267 56519 15331
rect 56583 15267 56609 15331
rect 56493 15251 56609 15267
rect 56493 15187 56519 15251
rect 56583 15187 56609 15251
rect 56493 15171 56609 15187
rect 56493 15107 56519 15171
rect 56583 15107 56609 15171
rect 56493 15091 56609 15107
rect 56493 15027 56519 15091
rect 56583 15027 56609 15091
rect 56493 15011 56609 15027
rect 56493 14947 56519 15011
rect 56583 14947 56609 15011
rect 56493 14931 56609 14947
rect 56493 14867 56519 14931
rect 56583 14867 56609 14931
rect 56493 14851 56609 14867
rect 56493 14787 56519 14851
rect 56583 14787 56609 14851
rect 56493 14771 56609 14787
rect 56493 14707 56519 14771
rect 56583 14707 56609 14771
rect 56493 14691 56609 14707
rect 56493 14627 56519 14691
rect 56583 14627 56609 14691
rect 56493 14611 56609 14627
rect 56493 14547 56519 14611
rect 56583 14547 56609 14611
rect 56493 14531 56609 14547
rect 56493 14467 56519 14531
rect 56583 14467 56609 14531
rect 56493 14451 56609 14467
rect 56493 14387 56519 14451
rect 56583 14387 56609 14451
rect 56493 14371 56609 14387
rect 56493 14307 56519 14371
rect 56583 14307 56609 14371
rect 56493 14291 56609 14307
rect 56493 14227 56519 14291
rect 56583 14227 56609 14291
rect 56493 14211 56609 14227
rect 56493 14147 56519 14211
rect 56583 14147 56609 14211
rect 56493 14131 56609 14147
rect 56493 14067 56519 14131
rect 56583 14067 56609 14131
rect 56493 14051 56609 14067
rect 56493 13987 56519 14051
rect 56583 13987 56609 14051
rect 56493 13971 56609 13987
rect 56493 13907 56519 13971
rect 56583 13907 56609 13971
rect 56493 13881 56609 13907
rect 1 7919 120001 8001
rect 1 6083 2083 7919
rect 3919 6083 13841 7919
rect 14397 6083 21841 7919
rect 22397 6083 29841 7919
rect 30397 6083 37841 7919
rect 38397 6083 45841 7919
rect 46397 6083 53841 7919
rect 54397 6083 61841 7919
rect 62397 6083 69841 7919
rect 70397 6083 77841 7919
rect 78397 6083 85841 7919
rect 86397 6083 93841 7919
rect 94397 6083 101841 7919
rect 102397 6083 112083 7919
rect 113919 6083 120001 7919
rect 1 6001 120001 6083
rect 1 3919 120001 4001
rect 1 2083 6083 3919
rect 7919 2083 17841 3919
rect 18397 2083 25841 3919
rect 26397 2083 33841 3919
rect 34397 2083 41841 3919
rect 42397 2083 49841 3919
rect 50397 2083 57841 3919
rect 58397 2083 65841 3919
rect 66397 2083 73841 3919
rect 74397 2083 81841 3919
rect 82397 2083 89841 3919
rect 90397 2083 97841 3919
rect 98397 2083 105841 3919
rect 106397 2083 116083 3919
rect 117919 2083 120001 3919
rect 1 2001 120001 2083
<< via4 >>
rect 2083 110546 3919 112382
rect 13841 110546 14397 112382
rect 21841 110546 22397 112382
rect 29841 110546 30397 112382
rect 37841 110546 38397 112382
rect 45841 110546 46397 112382
rect 53841 110546 54397 112382
rect 61841 110546 62397 112382
rect 69841 110546 70397 112382
rect 77841 110546 78397 112382
rect 85841 110546 86397 112382
rect 93841 110546 94397 112382
rect 101841 110546 102397 112382
rect 112083 110546 113919 112382
rect 6083 106546 7919 108382
rect 17841 106546 18397 108382
rect 25841 106546 26397 108382
rect 33841 106546 34397 108382
rect 41841 106546 42397 108382
rect 49841 106546 50397 108382
rect 57841 106546 58397 108382
rect 65841 106546 66397 108382
rect 73841 106546 74397 108382
rect 81841 106546 82397 108382
rect 89841 106546 90397 108382
rect 97841 106546 98397 108382
rect 105841 106546 106397 108382
rect 116083 106546 117919 108382
rect 38000 98852 38236 99088
rect 41998 99037 42234 99273
rect 69999 98956 70235 99192
rect 73998 98948 74234 99184
rect 41999 94778 42235 95014
rect 38000 94021 38236 94257
rect 42002 92699 42238 92935
rect 37996 90906 38232 91142
rect 46072 87285 46308 87521
rect 78001 88359 78237 88595
rect 85995 88365 86231 88601
rect 50157 87220 50393 87226
rect 50157 86996 50163 87220
rect 50163 86996 50387 87220
rect 50387 86996 50393 87220
rect 50157 86990 50393 86996
rect 54000 87195 54236 87431
rect 57998 87246 58234 87252
rect 57998 87022 58234 87246
rect 57998 87016 58234 87022
rect 74004 86368 74240 86604
rect 82000 86361 82236 86597
rect 90003 86357 90239 86593
rect 38003 74618 38239 74710
rect 38003 74554 38089 74618
rect 38089 74554 38153 74618
rect 38153 74554 38239 74618
rect 38003 74474 38239 74554
rect 30005 73742 30241 73846
rect 30005 73678 30044 73742
rect 30044 73678 30108 73742
rect 30108 73678 30124 73742
rect 30124 73678 30188 73742
rect 30188 73678 30204 73742
rect 30204 73678 30241 73742
rect 30005 73610 30241 73678
rect 34007 73007 34243 73243
rect 30040 67156 30087 67176
rect 30087 67156 30276 67176
rect 30040 67140 30276 67156
rect 30040 67076 30087 67140
rect 30087 67076 30276 67140
rect 30040 67060 30276 67076
rect 30040 66996 30087 67060
rect 30087 66996 30276 67060
rect 30040 66980 30276 66996
rect 30040 66940 30087 66980
rect 30087 66940 30276 66980
rect 50134 79115 50370 79351
rect 50134 78795 50370 79031
rect 54004 78206 54240 78442
rect 57997 83908 58233 84144
rect 66002 83897 66238 84133
rect 57997 80533 58233 80769
rect 66001 80522 66237 80758
rect 57997 77158 58233 77394
rect 66001 77147 66237 77383
rect 50004 75485 50240 75721
rect 30045 63929 30092 63970
rect 30092 63929 30281 63970
rect 30045 63913 30281 63929
rect 30045 63849 30092 63913
rect 30092 63849 30281 63913
rect 30045 63833 30281 63849
rect 30045 63769 30092 63833
rect 30092 63769 30281 63833
rect 30045 63753 30281 63769
rect 30045 63734 30092 63753
rect 30092 63734 30281 63753
rect 21989 62282 22225 62518
rect 26001 62293 26237 62529
rect 25989 61195 26225 61431
rect 34015 61680 34251 61916
rect 42002 61953 42238 62189
rect 30045 59842 30089 59901
rect 30089 59842 30281 59901
rect 30045 59826 30281 59842
rect 30045 59762 30089 59826
rect 30089 59762 30281 59826
rect 30045 59746 30281 59762
rect 30045 59682 30089 59746
rect 30089 59682 30281 59746
rect 30045 59666 30281 59682
rect 30045 59665 30089 59666
rect 30089 59665 30281 59666
rect 54010 75079 54246 75121
rect 54010 74935 54246 75079
rect 54010 74885 54246 74935
rect 54004 72557 54240 72793
rect 57997 73783 58233 74019
rect 66001 73772 66237 74008
rect 78001 84359 78237 84595
rect 85995 84365 86231 84601
rect 74004 82368 74240 82604
rect 82000 82361 82236 82597
rect 90003 82357 90239 82593
rect 78001 80359 78237 80595
rect 85995 80365 86231 80601
rect 74004 78368 74240 78604
rect 82000 78361 82236 78597
rect 90003 78357 90239 78593
rect 78001 76359 78237 76595
rect 85995 76365 86231 76601
rect 74004 74368 74240 74604
rect 82000 74361 82236 74597
rect 90003 74357 90239 74593
rect 78001 72359 78237 72595
rect 85995 72365 86231 72601
rect 54000 68387 54236 68623
rect 57993 68298 58229 68534
rect 66001 67022 66237 67258
rect 54008 63850 54244 63906
rect 54008 63706 54244 63850
rect 58003 64653 58239 64889
rect 54008 63670 54244 63706
rect 57997 63224 58233 63460
rect 30043 56742 30081 56787
rect 30081 56742 30279 56787
rect 30043 56726 30279 56742
rect 30043 56662 30081 56726
rect 30081 56662 30279 56726
rect 30043 56646 30279 56662
rect 30043 56582 30081 56646
rect 30081 56582 30279 56646
rect 30043 56566 30279 56582
rect 30043 56551 30081 56566
rect 30081 56551 30279 56566
rect 38003 52492 38239 52728
rect 42007 51227 42243 51463
rect 21983 50692 22219 50928
rect 46004 51839 46240 52075
rect 37995 49821 38231 49830
rect 37995 49597 38010 49821
rect 38010 49597 38231 49821
rect 37995 49594 38231 49597
rect 42003 49602 42239 49838
rect 30013 49298 30249 49534
rect 34005 48701 34241 48937
rect 18002 47498 18238 47734
rect 38002 47514 38238 47750
rect 42004 47423 42240 47659
rect 45995 46938 46231 47174
rect 21989 43080 22225 43253
rect 21989 43017 22051 43080
rect 22051 43017 22067 43080
rect 22067 43017 22131 43080
rect 22131 43017 22147 43080
rect 22147 43017 22211 43080
rect 22211 43017 22225 43080
rect 62002 61837 62238 62073
rect 57998 60879 58234 61115
rect 62009 60444 62245 60680
rect 58015 59800 58251 60036
rect 65999 59812 66235 60048
rect 62015 59266 62251 59502
rect 61987 47173 62223 47179
rect 61987 46949 62223 47173
rect 61987 46943 62223 46949
rect 65981 47355 66217 47515
rect 65981 47291 66031 47355
rect 66031 47291 66217 47355
rect 65981 47279 66217 47291
rect 74004 70368 74240 70604
rect 82000 70361 82236 70597
rect 90003 70357 90239 70593
rect 62004 43194 62240 43253
rect 30003 41747 30239 41983
rect 53996 41878 54232 41884
rect 53996 41654 54232 41878
rect 53996 41648 54232 41654
rect 18003 39984 18239 40220
rect 62004 43050 62240 43194
rect 62004 43017 62240 43050
rect 30010 38261 30246 38497
rect 33988 39274 34224 39510
rect 49989 39596 50225 39832
rect 54006 40234 54242 40470
rect 49986 38236 50222 38472
rect 49986 34696 50222 34932
rect 49996 33446 50232 33682
rect 49993 31257 50229 31263
rect 49993 31033 50229 31257
rect 49993 31027 50229 31033
rect 30002 30494 30238 30730
rect 49996 29548 50232 29784
rect 34009 28828 34245 29064
rect 54008 37832 54244 38068
rect 54006 32586 54242 32822
rect 54008 30527 54244 30763
rect 57996 41547 58232 41638
rect 57996 41483 58075 41547
rect 58075 41483 58139 41547
rect 58139 41483 58232 41547
rect 57996 41402 58232 41483
rect 65996 41187 66232 41423
rect 62001 40436 62237 40615
rect 62001 40379 62237 40436
rect 62001 40292 62237 40295
rect 62001 40059 62237 40292
rect 69958 45049 70194 45116
rect 69958 44985 70030 45049
rect 70030 44985 70094 45049
rect 70094 44985 70194 45049
rect 69958 44880 70194 44985
rect 69946 42710 70182 42815
rect 69946 42646 70024 42710
rect 70024 42646 70088 42710
rect 70088 42646 70182 42710
rect 69946 42579 70182 42646
rect 73986 42971 74222 43207
rect 77990 43084 78226 43180
rect 77990 43020 78065 43084
rect 78065 43020 78129 43084
rect 78129 43020 78226 43084
rect 77990 42944 78226 43020
rect 82000 42939 82236 43175
rect 69940 41105 70176 41210
rect 69940 41041 70050 41105
rect 70050 41041 70114 41105
rect 70114 41041 70176 41105
rect 69940 40974 70176 41041
rect 69959 39250 70195 39339
rect 69959 39186 70067 39250
rect 70067 39186 70131 39250
rect 70131 39186 70195 39250
rect 69959 39103 70195 39186
rect 73894 39378 74130 39614
rect 77933 39518 78169 39609
rect 77933 39454 78022 39518
rect 78022 39454 78086 39518
rect 78086 39454 78169 39518
rect 77933 39373 78169 39454
rect 82002 39346 82238 39582
rect 69981 37550 70217 37638
rect 69981 37486 70097 37550
rect 70097 37486 70161 37550
rect 70161 37486 70217 37550
rect 69981 37402 70217 37486
rect 69994 35698 70230 35783
rect 69994 35634 70095 35698
rect 70095 35634 70159 35698
rect 70159 35634 70230 35698
rect 69994 35547 70230 35634
rect 69990 34437 70226 34673
rect 77987 35928 78223 36021
rect 77987 35864 78079 35928
rect 78079 35864 78143 35928
rect 78143 35864 78223 35928
rect 77987 35785 78223 35864
rect 81990 35755 82226 35991
rect 58001 24243 58237 24345
rect 66021 24243 66257 24357
rect 73998 24243 74234 24345
rect 58001 24109 58237 24243
rect 66021 24121 66257 24243
rect 73998 24109 74234 24243
rect 89998 47918 90234 48154
rect 89997 45458 90233 45694
rect 90000 31077 90236 31313
rect 89991 29777 90227 30013
rect 89997 28362 90233 28598
rect 89993 26989 90229 27225
rect 102002 69094 102238 69194
rect 102002 69030 102012 69094
rect 102012 69030 102076 69094
rect 102076 69030 102092 69094
rect 102092 69030 102156 69094
rect 102156 69030 102172 69094
rect 102172 69030 102236 69094
rect 102236 69030 102238 69094
rect 102002 68958 102238 69030
rect 98007 68088 98243 68324
rect 102002 67943 102238 68033
rect 102002 67879 102035 67943
rect 102035 67879 102051 67943
rect 102051 67879 102115 67943
rect 102115 67879 102131 67943
rect 102131 67879 102195 67943
rect 102195 67879 102211 67943
rect 102211 67879 102238 67943
rect 102002 67797 102238 67879
rect 101986 65401 102222 65524
rect 101986 65337 102025 65401
rect 102025 65337 102041 65401
rect 102041 65337 102105 65401
rect 102105 65337 102121 65401
rect 102121 65337 102185 65401
rect 102185 65337 102201 65401
rect 102201 65337 102222 65401
rect 101986 65288 102222 65337
rect 98015 64343 98251 64579
rect 101979 64131 102215 64213
rect 101979 64067 102025 64131
rect 102025 64067 102041 64131
rect 102041 64067 102105 64131
rect 102105 64067 102121 64131
rect 102121 64067 102185 64131
rect 102185 64067 102201 64131
rect 102201 64067 102215 64131
rect 101979 63977 102215 64067
rect 102008 48173 102244 48272
rect 102008 48109 102049 48173
rect 102049 48109 102065 48173
rect 102065 48109 102129 48173
rect 102129 48109 102145 48173
rect 102145 48109 102209 48173
rect 102209 48109 102225 48173
rect 102225 48109 102244 48173
rect 102008 48036 102244 48109
rect 94011 46831 94247 46837
rect 94011 46607 94017 46831
rect 94017 46607 94241 46831
rect 94241 46607 94247 46831
rect 94011 46601 94247 46607
rect 98008 46516 98244 46752
rect 105998 45029 106234 45265
rect 93994 32808 94230 32813
rect 93994 32584 94001 32808
rect 94001 32584 94225 32808
rect 94225 32584 94230 32808
rect 93994 32577 94230 32584
rect 102003 31241 102239 31466
rect 98008 31184 98244 31190
rect 98008 30960 98244 31184
rect 102003 31230 102028 31241
rect 102028 31230 102044 31241
rect 102044 31230 102108 31241
rect 102108 31230 102124 31241
rect 102124 31230 102188 31241
rect 102188 31230 102204 31241
rect 102204 31230 102239 31241
rect 98008 30954 98244 30960
rect 94035 30311 94271 30547
rect 93996 29119 94081 29131
rect 94081 29119 94145 29131
rect 94145 29119 94232 29131
rect 93996 28895 94232 29119
rect 98006 28281 98242 28287
rect 98006 28057 98242 28281
rect 98006 28051 98242 28057
rect 94002 26599 94238 26835
rect 93994 25868 94230 25873
rect 93994 25644 94001 25868
rect 94001 25644 94225 25868
rect 94225 25644 94230 25868
rect 93994 25637 94230 25644
rect 90000 24137 90236 24373
rect 102006 24308 102242 24541
rect 98008 24244 98244 24250
rect 98008 24020 98244 24244
rect 102006 24305 102030 24308
rect 102030 24305 102046 24308
rect 102046 24305 102110 24308
rect 102110 24305 102126 24308
rect 102126 24305 102190 24308
rect 102190 24305 102206 24308
rect 102206 24305 102242 24308
rect 98008 24014 98244 24020
rect 94035 23371 94271 23607
rect 89991 22837 90227 23073
rect 93996 22179 94081 22191
rect 94081 22179 94145 22191
rect 94145 22179 94232 22191
rect 93996 21955 94232 22179
rect 89997 21422 90233 21658
rect 89993 20049 90229 20285
rect 97999 21341 98235 21343
rect 97999 21117 98235 21341
rect 97999 21107 98235 21117
rect 94002 19659 94238 19895
rect 54009 17611 54245 17847
rect 50003 15508 50239 15744
rect 2083 6083 3919 7919
rect 13841 6083 14397 7919
rect 21841 6083 22397 7919
rect 29841 6083 30397 7919
rect 37841 6083 38397 7919
rect 45841 6083 46397 7919
rect 53841 6083 54397 7919
rect 61841 6083 62397 7919
rect 69841 6083 70397 7919
rect 77841 6083 78397 7919
rect 85841 6083 86397 7919
rect 93841 6083 94397 7919
rect 101841 6083 102397 7919
rect 112083 6083 113919 7919
rect 6083 2083 7919 3919
rect 17841 2083 18397 3919
rect 25841 2083 26397 3919
rect 33841 2083 34397 3919
rect 41841 2083 42397 3919
rect 49841 2083 50397 3919
rect 57841 2083 58397 3919
rect 65841 2083 66397 3919
rect 73841 2083 74397 3919
rect 81841 2083 82397 3919
rect 89841 2083 90397 3919
rect 97841 2083 98397 3919
rect 105841 2083 106397 3919
rect 116083 2083 117919 3919
<< metal5 >>
rect 2001 112488 4001 114464
rect 1977 112382 4025 112488
rect 1977 110546 2083 112382
rect 3919 110546 4025 112382
rect 1977 110440 4025 110546
rect 2001 8025 4001 110440
rect 6001 108488 8001 114463
rect 112001 112488 114001 114463
rect 13785 112382 14453 112488
rect 13785 110546 13841 112382
rect 14397 110546 14453 112382
rect 13785 110440 14453 110546
rect 5977 108382 8025 108488
rect 5977 106546 6083 108382
rect 7919 106546 8025 108382
rect 5977 106440 8025 106546
rect 1977 7919 4025 8025
rect 1977 6083 2083 7919
rect 3919 6083 4025 7919
rect 1977 5977 4025 6083
rect 2001 1 4001 5977
rect 6001 4025 8001 106440
rect 13809 8025 14429 110440
rect 17809 108488 18429 112488
rect 21785 112382 22453 112488
rect 21785 110546 21841 112382
rect 22397 110546 22453 112382
rect 21785 110440 22453 110546
rect 17785 108382 18453 108488
rect 17785 106546 17841 108382
rect 18397 106546 18453 108382
rect 17785 106440 18453 106546
rect 17809 47734 18429 106440
rect 17809 47498 18002 47734
rect 18238 47498 18429 47734
rect 17809 40220 18429 47498
rect 17809 39984 18003 40220
rect 18239 39984 18429 40220
rect 13785 7919 14453 8025
rect 13785 6083 13841 7919
rect 14397 6083 14453 7919
rect 13785 5977 14453 6083
rect 5977 3919 8025 4025
rect 5977 2083 6083 3919
rect 7919 2083 8025 3919
rect 5977 1977 8025 2083
rect 13809 1977 14429 5977
rect 17809 4025 18429 39984
rect 21809 62518 22429 110440
rect 25809 108488 26429 112488
rect 29785 112382 30453 112488
rect 29785 110546 29841 112382
rect 30397 110546 30453 112382
rect 29785 110440 30453 110546
rect 25785 108382 26453 108488
rect 25785 106546 25841 108382
rect 26397 106546 26453 108382
rect 25785 106440 26453 106546
rect 21809 62282 21989 62518
rect 22225 62282 22429 62518
rect 21809 50928 22429 62282
rect 21809 50692 21983 50928
rect 22219 50692 22429 50928
rect 21809 43253 22429 50692
rect 21809 43017 21989 43253
rect 22225 43017 22429 43253
rect 21809 8025 22429 43017
rect 25809 62529 26429 106440
rect 25809 62293 26001 62529
rect 26237 62293 26429 62529
rect 25809 61431 26429 62293
rect 25809 61195 25989 61431
rect 26225 61195 26429 61431
rect 21785 7919 22453 8025
rect 21785 6083 21841 7919
rect 22397 6083 22453 7919
rect 21785 5977 22453 6083
rect 17785 3919 18453 4025
rect 17785 2083 17841 3919
rect 18397 2083 18453 3919
rect 17785 1977 18453 2083
rect 21809 1977 22429 5977
rect 25809 4025 26429 61195
rect 29809 73846 30429 110440
rect 33809 108488 34429 112488
rect 37785 112382 38453 112488
rect 37785 110546 37841 112382
rect 38397 110546 38453 112382
rect 37785 110440 38453 110546
rect 33785 108382 34453 108488
rect 33785 106546 33841 108382
rect 34397 106546 34453 108382
rect 33785 106440 34453 106546
rect 29809 73610 30005 73846
rect 30241 73610 30429 73846
rect 29809 67176 30429 73610
rect 29809 66940 30040 67176
rect 30276 66940 30429 67176
rect 29809 63970 30429 66940
rect 29809 63734 30045 63970
rect 30281 63734 30429 63970
rect 29809 59901 30429 63734
rect 29809 59665 30045 59901
rect 30281 59665 30429 59901
rect 29809 56787 30429 59665
rect 29809 56551 30043 56787
rect 30279 56551 30429 56787
rect 29809 49534 30429 56551
rect 29809 49298 30013 49534
rect 30249 49298 30429 49534
rect 29809 41983 30429 49298
rect 29809 41747 30003 41983
rect 30239 41747 30429 41983
rect 29809 38497 30429 41747
rect 29809 38261 30010 38497
rect 30246 38261 30429 38497
rect 29809 30730 30429 38261
rect 29809 30494 30002 30730
rect 30238 30494 30429 30730
rect 29809 8025 30429 30494
rect 33809 73243 34429 106440
rect 33809 73007 34007 73243
rect 34243 73007 34429 73243
rect 33809 61916 34429 73007
rect 33809 61680 34015 61916
rect 34251 61680 34429 61916
rect 33809 48937 34429 61680
rect 33809 48701 34005 48937
rect 34241 48701 34429 48937
rect 33809 39510 34429 48701
rect 33809 39274 33988 39510
rect 34224 39274 34429 39510
rect 33809 29064 34429 39274
rect 33809 28828 34009 29064
rect 34245 28828 34429 29064
rect 29785 7919 30453 8025
rect 29785 6083 29841 7919
rect 30397 6083 30453 7919
rect 29785 5977 30453 6083
rect 25785 3919 26453 4025
rect 25785 2083 25841 3919
rect 26397 2083 26453 3919
rect 25785 1977 26453 2083
rect 29809 1977 30429 5977
rect 33809 4025 34429 28828
rect 37809 99088 38429 110440
rect 41809 108488 42429 112488
rect 45785 112382 46453 112488
rect 45785 110546 45841 112382
rect 46397 110546 46453 112382
rect 45785 110440 46453 110546
rect 41785 108382 42453 108488
rect 41785 106546 41841 108382
rect 42397 106546 42453 108382
rect 41785 106440 42453 106546
rect 37809 98852 38000 99088
rect 38236 98852 38429 99088
rect 37809 94257 38429 98852
rect 37809 94021 38000 94257
rect 38236 94021 38429 94257
rect 37809 91142 38429 94021
rect 37809 90906 37996 91142
rect 38232 90906 38429 91142
rect 37809 74710 38429 90906
rect 37809 74474 38003 74710
rect 38239 74474 38429 74710
rect 37809 52728 38429 74474
rect 37809 52492 38003 52728
rect 38239 52492 38429 52728
rect 37809 49830 38429 52492
rect 37809 49594 37995 49830
rect 38231 49594 38429 49830
rect 37809 47750 38429 49594
rect 37809 47514 38002 47750
rect 38238 47514 38429 47750
rect 37809 8025 38429 47514
rect 41809 99273 42429 106440
rect 41809 99037 41998 99273
rect 42234 99037 42429 99273
rect 41809 95014 42429 99037
rect 41809 94778 41999 95014
rect 42235 94778 42429 95014
rect 41809 92935 42429 94778
rect 41809 92699 42002 92935
rect 42238 92699 42429 92935
rect 41809 62189 42429 92699
rect 41809 61953 42002 62189
rect 42238 61953 42429 62189
rect 41809 51463 42429 61953
rect 41809 51227 42007 51463
rect 42243 51227 42429 51463
rect 41809 49838 42429 51227
rect 41809 49602 42003 49838
rect 42239 49602 42429 49838
rect 41809 47659 42429 49602
rect 41809 47423 42004 47659
rect 42240 47423 42429 47659
rect 37785 7919 38453 8025
rect 37785 6083 37841 7919
rect 38397 6083 38453 7919
rect 37785 5977 38453 6083
rect 33785 3919 34453 4025
rect 33785 2083 33841 3919
rect 34397 2083 34453 3919
rect 33785 1977 34453 2083
rect 37809 1977 38429 5977
rect 41809 4025 42429 47423
rect 45809 87521 46429 110440
rect 49809 108488 50429 112488
rect 53785 112382 54453 112488
rect 53785 110546 53841 112382
rect 54397 110546 54453 112382
rect 53785 110440 54453 110546
rect 49785 108382 50453 108488
rect 49785 106546 49841 108382
rect 50397 106546 50453 108382
rect 49785 106440 50453 106546
rect 45809 87285 46072 87521
rect 46308 87285 46429 87521
rect 45809 52075 46429 87285
rect 45809 51839 46004 52075
rect 46240 51839 46429 52075
rect 45809 47174 46429 51839
rect 45809 46938 45995 47174
rect 46231 46938 46429 47174
rect 45809 8025 46429 46938
rect 49809 87226 50429 106440
rect 49809 86990 50157 87226
rect 50393 86990 50429 87226
rect 49809 79351 50429 86990
rect 49809 79115 50134 79351
rect 50370 79115 50429 79351
rect 49809 79031 50429 79115
rect 49809 78795 50134 79031
rect 50370 78795 50429 79031
rect 49809 75721 50429 78795
rect 49809 75485 50004 75721
rect 50240 75485 50429 75721
rect 49809 39832 50429 75485
rect 49809 39596 49989 39832
rect 50225 39596 50429 39832
rect 49809 38472 50429 39596
rect 49809 38236 49986 38472
rect 50222 38236 50429 38472
rect 49809 34932 50429 38236
rect 49809 34696 49986 34932
rect 50222 34696 50429 34932
rect 49809 33682 50429 34696
rect 49809 33446 49996 33682
rect 50232 33446 50429 33682
rect 49809 31263 50429 33446
rect 49809 31027 49993 31263
rect 50229 31027 50429 31263
rect 49809 29784 50429 31027
rect 49809 29548 49996 29784
rect 50232 29548 50429 29784
rect 49809 15744 50429 29548
rect 49809 15508 50003 15744
rect 50239 15508 50429 15744
rect 45785 7919 46453 8025
rect 45785 6083 45841 7919
rect 46397 6083 46453 7919
rect 45785 5977 46453 6083
rect 41785 3919 42453 4025
rect 41785 2083 41841 3919
rect 42397 2083 42453 3919
rect 41785 1977 42453 2083
rect 45809 1977 46429 5977
rect 49809 4025 50429 15508
rect 53809 87431 54429 110440
rect 57809 108488 58429 112488
rect 61785 112382 62453 112488
rect 61785 110546 61841 112382
rect 62397 110546 62453 112382
rect 61785 110440 62453 110546
rect 57785 108382 58453 108488
rect 57785 106546 57841 108382
rect 58397 106546 58453 108382
rect 57785 106440 58453 106546
rect 53809 87195 54000 87431
rect 54236 87195 54429 87431
rect 53809 78442 54429 87195
rect 53809 78206 54004 78442
rect 54240 78206 54429 78442
rect 53809 75121 54429 78206
rect 53809 74885 54010 75121
rect 54246 74885 54429 75121
rect 53809 72793 54429 74885
rect 53809 72557 54004 72793
rect 54240 72557 54429 72793
rect 53809 68623 54429 72557
rect 53809 68387 54000 68623
rect 54236 68387 54429 68623
rect 53809 63906 54429 68387
rect 53809 63670 54008 63906
rect 54244 63670 54429 63906
rect 53809 41884 54429 63670
rect 53809 41648 53996 41884
rect 54232 41648 54429 41884
rect 53809 40470 54429 41648
rect 53809 40234 54006 40470
rect 54242 40234 54429 40470
rect 53809 38068 54429 40234
rect 53809 37832 54008 38068
rect 54244 37832 54429 38068
rect 53809 32822 54429 37832
rect 53809 32586 54006 32822
rect 54242 32586 54429 32822
rect 53809 30763 54429 32586
rect 53809 30527 54008 30763
rect 54244 30527 54429 30763
rect 53809 17847 54429 30527
rect 53809 17611 54009 17847
rect 54245 17611 54429 17847
rect 53809 8025 54429 17611
rect 57809 87252 58429 106440
rect 57809 87016 57998 87252
rect 58234 87016 58429 87252
rect 57809 84144 58429 87016
rect 57809 83908 57997 84144
rect 58233 83908 58429 84144
rect 57809 80769 58429 83908
rect 57809 80533 57997 80769
rect 58233 80533 58429 80769
rect 57809 77394 58429 80533
rect 57809 77158 57997 77394
rect 58233 77158 58429 77394
rect 57809 74019 58429 77158
rect 57809 73783 57997 74019
rect 58233 73783 58429 74019
rect 57809 68534 58429 73783
rect 57809 68298 57993 68534
rect 58229 68298 58429 68534
rect 57809 64889 58429 68298
rect 57809 64653 58003 64889
rect 58239 64653 58429 64889
rect 57809 63460 58429 64653
rect 57809 63224 57997 63460
rect 58233 63224 58429 63460
rect 57809 61115 58429 63224
rect 57809 60879 57998 61115
rect 58234 60879 58429 61115
rect 57809 60036 58429 60879
rect 57809 59800 58015 60036
rect 58251 59800 58429 60036
rect 57809 41638 58429 59800
rect 57809 41402 57996 41638
rect 58232 41402 58429 41638
rect 57809 24345 58429 41402
rect 57809 24109 58001 24345
rect 58237 24109 58429 24345
rect 53785 7919 54453 8025
rect 53785 6083 53841 7919
rect 54397 6083 54453 7919
rect 53785 5977 54453 6083
rect 49785 3919 50453 4025
rect 49785 2083 49841 3919
rect 50397 2083 50453 3919
rect 49785 1977 50453 2083
rect 53809 1977 54429 5977
rect 57809 4025 58429 24109
rect 61809 62073 62429 110440
rect 65809 108488 66429 112488
rect 69785 112382 70453 112488
rect 69785 110546 69841 112382
rect 70397 110546 70453 112382
rect 69785 110440 70453 110546
rect 65785 108382 66453 108488
rect 65785 106546 65841 108382
rect 66397 106546 66453 108382
rect 65785 106440 66453 106546
rect 61809 61837 62002 62073
rect 62238 61837 62429 62073
rect 61809 60680 62429 61837
rect 61809 60444 62009 60680
rect 62245 60444 62429 60680
rect 61809 59502 62429 60444
rect 61809 59266 62015 59502
rect 62251 59266 62429 59502
rect 61809 47179 62429 59266
rect 61809 46943 61987 47179
rect 62223 46943 62429 47179
rect 61809 43253 62429 46943
rect 61809 43017 62004 43253
rect 62240 43017 62429 43253
rect 61809 40615 62429 43017
rect 61809 40379 62001 40615
rect 62237 40379 62429 40615
rect 61809 40295 62429 40379
rect 61809 40059 62001 40295
rect 62237 40059 62429 40295
rect 61809 8025 62429 40059
rect 65809 84133 66429 106440
rect 65809 83897 66002 84133
rect 66238 83897 66429 84133
rect 65809 80758 66429 83897
rect 65809 80522 66001 80758
rect 66237 80522 66429 80758
rect 65809 77383 66429 80522
rect 65809 77147 66001 77383
rect 66237 77147 66429 77383
rect 65809 74008 66429 77147
rect 65809 73772 66001 74008
rect 66237 73772 66429 74008
rect 65809 67258 66429 73772
rect 65809 67022 66001 67258
rect 66237 67022 66429 67258
rect 65809 60048 66429 67022
rect 65809 59812 65999 60048
rect 66235 59812 66429 60048
rect 65809 47515 66429 59812
rect 65809 47279 65981 47515
rect 66217 47279 66429 47515
rect 65809 41423 66429 47279
rect 65809 41187 65996 41423
rect 66232 41187 66429 41423
rect 65809 24357 66429 41187
rect 65809 24121 66021 24357
rect 66257 24121 66429 24357
rect 61785 7919 62453 8025
rect 61785 6083 61841 7919
rect 62397 6083 62453 7919
rect 61785 5977 62453 6083
rect 57785 3919 58453 4025
rect 57785 2083 57841 3919
rect 58397 2083 58453 3919
rect 57785 1977 58453 2083
rect 61809 1977 62429 5977
rect 65809 4025 66429 24121
rect 69809 99192 70429 110440
rect 73809 108488 74429 112488
rect 77785 112382 78453 112488
rect 77785 110546 77841 112382
rect 78397 110546 78453 112382
rect 77785 110440 78453 110546
rect 73785 108382 74453 108488
rect 73785 106546 73841 108382
rect 74397 106546 74453 108382
rect 73785 106440 74453 106546
rect 69809 98956 69999 99192
rect 70235 98956 70429 99192
rect 69809 45116 70429 98956
rect 69809 44880 69958 45116
rect 70194 44880 70429 45116
rect 69809 42815 70429 44880
rect 69809 42579 69946 42815
rect 70182 42579 70429 42815
rect 69809 41210 70429 42579
rect 69809 40974 69940 41210
rect 70176 40974 70429 41210
rect 69809 39339 70429 40974
rect 69809 39103 69959 39339
rect 70195 39103 70429 39339
rect 69809 37638 70429 39103
rect 69809 37402 69981 37638
rect 70217 37402 70429 37638
rect 69809 35783 70429 37402
rect 69809 35547 69994 35783
rect 70230 35547 70429 35783
rect 69809 34673 70429 35547
rect 69809 34437 69990 34673
rect 70226 34437 70429 34673
rect 69809 8025 70429 34437
rect 73809 99184 74429 106440
rect 73809 98948 73998 99184
rect 74234 98948 74429 99184
rect 73809 86604 74429 98948
rect 73809 86368 74004 86604
rect 74240 86368 74429 86604
rect 73809 82604 74429 86368
rect 73809 82368 74004 82604
rect 74240 82368 74429 82604
rect 73809 78604 74429 82368
rect 73809 78368 74004 78604
rect 74240 78368 74429 78604
rect 73809 74604 74429 78368
rect 73809 74368 74004 74604
rect 74240 74368 74429 74604
rect 73809 70604 74429 74368
rect 73809 70368 74004 70604
rect 74240 70368 74429 70604
rect 73809 43207 74429 70368
rect 73809 42971 73986 43207
rect 74222 42971 74429 43207
rect 73809 39614 74429 42971
rect 73809 39378 73894 39614
rect 74130 39378 74429 39614
rect 73809 24345 74429 39378
rect 73809 24109 73998 24345
rect 74234 24109 74429 24345
rect 69785 7919 70453 8025
rect 69785 6083 69841 7919
rect 70397 6083 70453 7919
rect 69785 5977 70453 6083
rect 65785 3919 66453 4025
rect 65785 2083 65841 3919
rect 66397 2083 66453 3919
rect 65785 1977 66453 2083
rect 69809 1977 70429 5977
rect 73809 4025 74429 24109
rect 77809 88595 78429 110440
rect 81809 108488 82429 112488
rect 85785 112382 86453 112488
rect 85785 110546 85841 112382
rect 86397 110546 86453 112382
rect 85785 110440 86453 110546
rect 81785 108382 82453 108488
rect 81785 106546 81841 108382
rect 82397 106546 82453 108382
rect 81785 106440 82453 106546
rect 77809 88359 78001 88595
rect 78237 88359 78429 88595
rect 77809 84595 78429 88359
rect 77809 84359 78001 84595
rect 78237 84359 78429 84595
rect 77809 80595 78429 84359
rect 77809 80359 78001 80595
rect 78237 80359 78429 80595
rect 77809 76595 78429 80359
rect 77809 76359 78001 76595
rect 78237 76359 78429 76595
rect 77809 72595 78429 76359
rect 77809 72359 78001 72595
rect 78237 72359 78429 72595
rect 77809 43180 78429 72359
rect 77809 42944 77990 43180
rect 78226 42944 78429 43180
rect 77809 39609 78429 42944
rect 77809 39373 77933 39609
rect 78169 39373 78429 39609
rect 77809 36021 78429 39373
rect 77809 35785 77987 36021
rect 78223 35785 78429 36021
rect 77809 8025 78429 35785
rect 81809 86597 82429 106440
rect 81809 86361 82000 86597
rect 82236 86361 82429 86597
rect 81809 82597 82429 86361
rect 81809 82361 82000 82597
rect 82236 82361 82429 82597
rect 81809 78597 82429 82361
rect 81809 78361 82000 78597
rect 82236 78361 82429 78597
rect 81809 74597 82429 78361
rect 81809 74361 82000 74597
rect 82236 74361 82429 74597
rect 81809 70597 82429 74361
rect 81809 70361 82000 70597
rect 82236 70361 82429 70597
rect 81809 43175 82429 70361
rect 81809 42939 82000 43175
rect 82236 42939 82429 43175
rect 81809 39582 82429 42939
rect 81809 39346 82002 39582
rect 82238 39346 82429 39582
rect 81809 35991 82429 39346
rect 81809 35755 81990 35991
rect 82226 35755 82429 35991
rect 77785 7919 78453 8025
rect 77785 6083 77841 7919
rect 78397 6083 78453 7919
rect 77785 5977 78453 6083
rect 73785 3919 74453 4025
rect 73785 2083 73841 3919
rect 74397 2083 74453 3919
rect 73785 1977 74453 2083
rect 77809 1977 78429 5977
rect 81809 4025 82429 35755
rect 85809 88601 86429 110440
rect 89809 108488 90429 112488
rect 93785 112382 94453 112488
rect 93785 110546 93841 112382
rect 94397 110546 94453 112382
rect 93785 110440 94453 110546
rect 89785 108382 90453 108488
rect 89785 106546 89841 108382
rect 90397 106546 90453 108382
rect 89785 106440 90453 106546
rect 85809 88365 85995 88601
rect 86231 88365 86429 88601
rect 85809 84601 86429 88365
rect 85809 84365 85995 84601
rect 86231 84365 86429 84601
rect 85809 80601 86429 84365
rect 85809 80365 85995 80601
rect 86231 80365 86429 80601
rect 85809 76601 86429 80365
rect 85809 76365 85995 76601
rect 86231 76365 86429 76601
rect 85809 72601 86429 76365
rect 85809 72365 85995 72601
rect 86231 72365 86429 72601
rect 85809 8025 86429 72365
rect 89809 86593 90429 106440
rect 89809 86357 90003 86593
rect 90239 86357 90429 86593
rect 89809 82593 90429 86357
rect 89809 82357 90003 82593
rect 90239 82357 90429 82593
rect 89809 78593 90429 82357
rect 89809 78357 90003 78593
rect 90239 78357 90429 78593
rect 89809 74593 90429 78357
rect 89809 74357 90003 74593
rect 90239 74357 90429 74593
rect 89809 70593 90429 74357
rect 89809 70357 90003 70593
rect 90239 70357 90429 70593
rect 89809 48154 90429 70357
rect 89809 47918 89998 48154
rect 90234 47918 90429 48154
rect 89809 45694 90429 47918
rect 89809 45458 89997 45694
rect 90233 45458 90429 45694
rect 89809 31313 90429 45458
rect 89809 31077 90000 31313
rect 90236 31077 90429 31313
rect 89809 30013 90429 31077
rect 89809 29777 89991 30013
rect 90227 29777 90429 30013
rect 89809 28598 90429 29777
rect 89809 28362 89997 28598
rect 90233 28362 90429 28598
rect 89809 27225 90429 28362
rect 89809 26989 89993 27225
rect 90229 26989 90429 27225
rect 89809 24373 90429 26989
rect 89809 24137 90000 24373
rect 90236 24137 90429 24373
rect 89809 23073 90429 24137
rect 89809 22837 89991 23073
rect 90227 22837 90429 23073
rect 89809 21658 90429 22837
rect 89809 21422 89997 21658
rect 90233 21422 90429 21658
rect 89809 20285 90429 21422
rect 89809 20049 89993 20285
rect 90229 20049 90429 20285
rect 85785 7919 86453 8025
rect 85785 6083 85841 7919
rect 86397 6083 86453 7919
rect 85785 5977 86453 6083
rect 81785 3919 82453 4025
rect 81785 2083 81841 3919
rect 82397 2083 82453 3919
rect 81785 1977 82453 2083
rect 85809 1977 86429 5977
rect 89809 4025 90429 20049
rect 93809 46837 94429 110440
rect 97809 108488 98429 112488
rect 101785 112382 102453 112488
rect 101785 110546 101841 112382
rect 102397 110546 102453 112382
rect 101785 110440 102453 110546
rect 97785 108382 98453 108488
rect 97785 106546 97841 108382
rect 98397 106546 98453 108382
rect 97785 106440 98453 106546
rect 93809 46601 94011 46837
rect 94247 46601 94429 46837
rect 93809 32813 94429 46601
rect 93809 32577 93994 32813
rect 94230 32577 94429 32813
rect 93809 30547 94429 32577
rect 93809 30311 94035 30547
rect 94271 30311 94429 30547
rect 93809 29131 94429 30311
rect 93809 28895 93996 29131
rect 94232 28895 94429 29131
rect 93809 26835 94429 28895
rect 93809 26599 94002 26835
rect 94238 26599 94429 26835
rect 93809 25873 94429 26599
rect 93809 25637 93994 25873
rect 94230 25637 94429 25873
rect 93809 23607 94429 25637
rect 93809 23371 94035 23607
rect 94271 23371 94429 23607
rect 93809 22191 94429 23371
rect 93809 21955 93996 22191
rect 94232 21955 94429 22191
rect 93809 19895 94429 21955
rect 93809 19659 94002 19895
rect 94238 19659 94429 19895
rect 93809 8025 94429 19659
rect 97809 68324 98429 106440
rect 97809 68088 98007 68324
rect 98243 68088 98429 68324
rect 97809 64579 98429 68088
rect 97809 64343 98015 64579
rect 98251 64343 98429 64579
rect 97809 46752 98429 64343
rect 97809 46516 98008 46752
rect 98244 46516 98429 46752
rect 97809 31190 98429 46516
rect 97809 30954 98008 31190
rect 98244 30954 98429 31190
rect 97809 28287 98429 30954
rect 97809 28051 98006 28287
rect 98242 28051 98429 28287
rect 97809 24250 98429 28051
rect 97809 24014 98008 24250
rect 98244 24014 98429 24250
rect 97809 21343 98429 24014
rect 97809 21107 97999 21343
rect 98235 21107 98429 21343
rect 93785 7919 94453 8025
rect 93785 6083 93841 7919
rect 94397 6083 94453 7919
rect 93785 5977 94453 6083
rect 89785 3919 90453 4025
rect 89785 2083 89841 3919
rect 90397 2083 90453 3919
rect 89785 1977 90453 2083
rect 93809 1977 94429 5977
rect 97809 4025 98429 21107
rect 101809 69194 102429 110440
rect 105809 108488 106429 112488
rect 111977 112382 114025 112488
rect 111977 110546 112083 112382
rect 113919 110546 114025 112382
rect 111977 110440 114025 110546
rect 105785 108382 106453 108488
rect 105785 106546 105841 108382
rect 106397 106546 106453 108382
rect 105785 106440 106453 106546
rect 101809 68958 102002 69194
rect 102238 68958 102429 69194
rect 101809 68033 102429 68958
rect 101809 67797 102002 68033
rect 102238 67797 102429 68033
rect 101809 65524 102429 67797
rect 101809 65288 101986 65524
rect 102222 65288 102429 65524
rect 101809 64213 102429 65288
rect 101809 63977 101979 64213
rect 102215 63977 102429 64213
rect 101809 48272 102429 63977
rect 101809 48036 102008 48272
rect 102244 48036 102429 48272
rect 101809 31466 102429 48036
rect 101809 31230 102003 31466
rect 102239 31230 102429 31466
rect 101809 24541 102429 31230
rect 101809 24305 102006 24541
rect 102242 24305 102429 24541
rect 101809 8025 102429 24305
rect 105809 45265 106429 106440
rect 105809 45029 105998 45265
rect 106234 45029 106429 45265
rect 101785 7919 102453 8025
rect 101785 6083 101841 7919
rect 102397 6083 102453 7919
rect 101785 5977 102453 6083
rect 97785 3919 98453 4025
rect 97785 2083 97841 3919
rect 98397 2083 98453 3919
rect 97785 1977 98453 2083
rect 101809 1977 102429 5977
rect 105809 4025 106429 45029
rect 112001 8025 114001 110440
rect 116001 108488 118001 114463
rect 115977 108382 118025 108488
rect 115977 106546 116083 108382
rect 117919 106546 118025 108382
rect 115977 106440 118025 106546
rect 111977 7919 114025 8025
rect 111977 6083 112083 7919
rect 113919 6083 114025 7919
rect 111977 5977 114025 6083
rect 105785 3919 106453 4025
rect 105785 2083 105841 3919
rect 106397 2083 106453 3919
rect 105785 1977 106453 2083
rect 6001 1 8001 1977
rect 112001 1 114001 5977
rect 116001 4025 118001 106440
rect 115977 3919 118025 4025
rect 115977 2083 116083 3919
rect 117919 2083 118025 3919
rect 115977 1977 118025 2083
rect 116001 1 118001 1977
use a_mux2_en  a_mux2_en_0
timestamp 1654583406
transform 0 -1 40510 1 0 92748
box -2638 -2585 3429 115
use a_mux2_en  a_mux2_en_1
timestamp 1654583406
transform 1 0 93424 0 1 47919
box -2638 -2585 3429 115
use a_mux4_en  a_mux4_en_0
timestamp 1654583406
transform 1 0 94177 0 1 32348
box -3690 -5314 3456 148
use a_mux4_en  a_mux4_en_1
timestamp 1654583406
transform 1 0 94177 0 1 25408
box -3690 -5314 3456 148
use analog_top  analog_top_0
timestamp 1654583406
transform 1 0 57094 0 1 24022
box -57094 -24022 62907 90442
use clock_v2  clock_v2_0
timestamp 1654583406
transform 0 1 88714 -1 0 86659
box -3621 -14204 17033 36
use comparator_v2  comparator_v2_0
timestamp 1654583406
transform 0 -1 38113 -1 0 63586
box -3788 -193 7250 10729
use esd_cell  esd_cell_0
timestamp 1654583101
transform 0 -1 71300 1 0 97341
box -65 -55 3553 3095
use esd_cell  esd_cell_1
timestamp 1654583101
transform 0 -1 43296 1 0 97341
box -65 -55 3553 3095
use esd_cell  esd_cell_2
timestamp 1654583101
transform 1 0 99871 0 1 45144
box -65 -55 3553 3095
use esd_cell  esd_cell_3
timestamp 1654583101
transform 1 0 18834 0 1 40049
box -65 -55 3553 3095
use esd_cell  esd_cell_4
timestamp 1654583101
transform 1 0 18834 0 1 47579
box -65 -55 3553 3095
use esd_cell  esd_cell_5
timestamp 1654583101
transform 1 0 99616 0 1 28211
box -65 -55 3553 3095
use esd_cell  esd_cell_6
timestamp 1654583101
transform 1 0 99616 0 1 21271
box -65 -55 3553 3095
use esd_cell  esd_cell_7
timestamp 1654583101
transform 0 1 53546 -1 0 17286
box -65 -55 3553 3095
use onebit_dac  onebit_dac_0
timestamp 1654583101
transform 1 0 40003 0 1 48458
box -313 -1154 1895 1114
use onebit_dac  onebit_dac_1
timestamp 1654583101
transform 1 0 40008 0 1 51100
box -313 -1154 1895 1114
use ota  ota_0
timestamp 1654583101
transform 0 -1 49949 1 0 71337
box -7664 -17587 18520 2944
use ota_w_test  ota_w_test_0
timestamp 1654583101
transform 1 0 64758 0 1 41664
box -7664 -17587 18520 2944
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_0
timestamp 1654583101
transform 0 1 66959 -1 0 57260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_1
timestamp 1654583101
transform 0 1 66959 -1 0 56260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_2
timestamp 1654583101
transform 0 1 64959 -1 0 57260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_3
timestamp 1654583101
transform 0 1 64959 -1 0 56260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_4
timestamp 1654583101
transform 0 1 65959 -1 0 57260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_5
timestamp 1654583101
transform 0 1 65959 -1 0 56260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_6
timestamp 1654583101
transform 0 -1 61959 -1 0 57260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_7
timestamp 1654583101
transform 0 -1 62959 -1 0 57260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_8
timestamp 1654583101
transform 0 -1 61959 -1 0 56260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_9
timestamp 1654583101
transform 0 -1 62959 -1 0 56260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_10
timestamp 1654583101
transform 0 1 63959 -1 0 57260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_11
timestamp 1654583101
transform 0 1 63959 -1 0 56260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_12
timestamp 1654583101
transform 0 -1 59959 -1 0 57260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_13
timestamp 1654583101
transform 0 -1 60959 -1 0 57260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_14
timestamp 1654583101
transform 0 -1 59959 -1 0 56260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_15
timestamp 1654583101
transform 0 -1 60959 -1 0 56260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_16
timestamp 1654583101
transform 0 1 66959 -1 0 55260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_17
timestamp 1654583101
transform 0 1 66959 -1 0 53260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_18
timestamp 1654583101
transform 0 1 66959 -1 0 54260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_19
timestamp 1654583101
transform 0 1 64959 -1 0 55260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_20
timestamp 1654583101
transform 0 1 64959 -1 0 54260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_21
timestamp 1654583101
transform 0 1 64959 -1 0 53260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_22
timestamp 1654583101
transform 0 1 65959 -1 0 55260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_23
timestamp 1654583101
transform 0 1 65959 -1 0 54260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_24
timestamp 1654583101
transform 0 1 65959 -1 0 53260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_25
timestamp 1654583101
transform 0 -1 61959 -1 0 55260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_26
timestamp 1654583101
transform 0 -1 62959 -1 0 55260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_27
timestamp 1654583101
transform 0 -1 61959 -1 0 53260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_28
timestamp 1654583101
transform 0 -1 61959 -1 0 54260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_29
timestamp 1654583101
transform 0 -1 62959 -1 0 53260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_30
timestamp 1654583101
transform 0 -1 62959 -1 0 54260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_31
timestamp 1654583101
transform 0 1 63959 -1 0 55260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_32
timestamp 1654583101
transform 0 1 63959 -1 0 54260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_33
timestamp 1654583101
transform 0 1 63959 -1 0 53260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_34
timestamp 1654583101
transform 0 -1 59959 -1 0 55260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_35
timestamp 1654583101
transform 0 -1 60959 -1 0 55260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_36
timestamp 1654583101
transform 0 -1 59959 -1 0 54260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_37
timestamp 1654583101
transform 0 -1 59959 -1 0 53260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_38
timestamp 1654583101
transform 0 -1 60959 -1 0 53260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_39
timestamp 1654583101
transform 0 -1 60959 -1 0 54260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_40
timestamp 1654583101
transform 0 1 65959 -1 0 52260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_41
timestamp 1654583101
transform 0 1 66959 -1 0 52260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_42
timestamp 1654583101
transform 0 -1 62959 -1 0 52260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_43
timestamp 1654583101
transform 0 1 63959 -1 0 52260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_44
timestamp 1654583101
transform 0 1 64959 -1 0 52260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_45
timestamp 1654583101
transform 0 -1 61959 -1 0 52260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_46
timestamp 1654583101
transform 0 -1 59959 -1 0 52260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_47
timestamp 1654583101
transform 0 -1 60959 -1 0 52260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_48
timestamp 1654583101
transform 0 1 66959 -1 0 49260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_49
timestamp 1654583101
transform 0 1 65959 -1 0 51260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_50
timestamp 1654583101
transform 0 1 65959 -1 0 49260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_51
timestamp 1654583101
transform 0 1 65959 -1 0 50260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_52
timestamp 1654583101
transform 0 1 66959 -1 0 51260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_53
timestamp 1654583101
transform 0 1 66959 -1 0 50260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_54
timestamp 1654583101
transform 0 -1 62959 -1 0 51260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_55
timestamp 1654583101
transform 0 -1 62959 -1 0 49260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_56
timestamp 1654583101
transform 0 -1 62959 -1 0 50260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_57
timestamp 1654583101
transform 0 1 63959 -1 0 51260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_58
timestamp 1654583101
transform 0 1 63959 -1 0 49260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_59
timestamp 1654583101
transform 0 1 63959 -1 0 50260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_60
timestamp 1654583101
transform 0 1 64959 -1 0 51260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_61
timestamp 1654583101
transform 0 1 64959 -1 0 49260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_62
timestamp 1654583101
transform 0 1 64959 -1 0 50260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_63
timestamp 1654583101
transform 0 -1 61959 -1 0 51260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_64
timestamp 1654583101
transform 0 -1 61959 -1 0 49260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_65
timestamp 1654583101
transform 0 -1 61959 -1 0 50260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_66
timestamp 1654583101
transform 0 -1 59959 -1 0 51260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_67
timestamp 1654583101
transform 0 -1 60959 -1 0 51260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_68
timestamp 1654583101
transform 0 -1 59959 -1 0 49260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_69
timestamp 1654583101
transform 0 -1 59959 -1 0 50260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_70
timestamp 1654583101
transform 0 -1 60959 -1 0 49260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CEWQ64  sky130_fd_pr__cap_mim_m3_1_CEWQ64_71
timestamp 1654583101
transform 0 -1 60959 -1 0 50260
box -360 -310 260 310
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_0
timestamp 1654583101
transform 1 0 48026 0 1 43298
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_1
timestamp 1654583101
transform 1 0 45426 0 1 43298
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_2
timestamp 1654583101
transform 1 0 42826 0 1 43298
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_3
timestamp 1654583101
transform 1 0 40226 0 1 43298
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_4
timestamp 1654583101
transform 1 0 37626 0 1 43298
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_5
timestamp 1654583101
transform 1 0 35026 0 1 43298
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_6
timestamp 1654583101
transform 1 0 48026 0 1 38098
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_7
timestamp 1654583101
transform 1 0 48026 0 1 40698
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_8
timestamp 1654583101
transform 1 0 48026 0 1 32898
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_9
timestamp 1654583101
transform 1 0 48026 0 1 35498
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_10
timestamp 1654583101
transform 1 0 48026 0 1 30298
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_11
timestamp 1654583101
transform 1 0 48026 0 1 27698
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_12
timestamp 1654583101
transform 1 0 48026 0 1 25098
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_13
timestamp 1654583101
transform 1 0 45426 0 1 40698
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_14
timestamp 1654583101
transform 1 0 42826 0 1 40698
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_15
timestamp 1654583101
transform 1 0 40226 0 1 40698
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_16
timestamp 1654583101
transform 1 0 37626 0 1 40698
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_17
timestamp 1654583101
transform 1 0 35026 0 1 40698
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_18
timestamp 1654583101
transform 1 0 45426 0 1 38098
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_19
timestamp 1654583101
transform 1 0 42826 0 1 38098
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_20
timestamp 1654583101
transform 1 0 40226 0 1 38098
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_21
timestamp 1654583101
transform 1 0 37626 0 1 38098
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_22
timestamp 1654583101
transform 1 0 35026 0 1 38098
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_23
timestamp 1654583101
transform 1 0 45426 0 1 35498
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_24
timestamp 1654583101
transform 1 0 42826 0 1 35498
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_25
timestamp 1654583101
transform 1 0 45426 0 1 32898
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_26
timestamp 1654583101
transform 1 0 42826 0 1 32898
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_27
timestamp 1654583101
transform 1 0 40226 0 1 35498
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_28
timestamp 1654583101
transform 1 0 37626 0 1 35498
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_29
timestamp 1654583101
transform 1 0 40226 0 1 32898
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_30
timestamp 1654583101
transform 1 0 37626 0 1 32898
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_31
timestamp 1654583101
transform 1 0 35026 0 1 32898
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_32
timestamp 1654583101
transform 1 0 35026 0 1 35498
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_33
timestamp 1654583101
transform 1 0 45426 0 1 27698
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_34
timestamp 1654583101
transform 1 0 42826 0 1 27698
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_35
timestamp 1654583101
transform 1 0 45426 0 1 30298
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_36
timestamp 1654583101
transform 1 0 42826 0 1 30298
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_37
timestamp 1654583101
transform 1 0 37626 0 1 27698
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_38
timestamp 1654583101
transform 1 0 40226 0 1 27698
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_39
timestamp 1654583101
transform 1 0 40226 0 1 30298
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_40
timestamp 1654583101
transform 1 0 37626 0 1 30298
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_41
timestamp 1654583101
transform 1 0 35026 0 1 30298
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_42
timestamp 1654583101
transform 1 0 35026 0 1 27698
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_43
timestamp 1654583101
transform 1 0 42826 0 1 25098
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_44
timestamp 1654583101
transform 1 0 45426 0 1 25098
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_45
timestamp 1654583101
transform 1 0 37626 0 1 25098
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_46
timestamp 1654583101
transform 1 0 40226 0 1 25098
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_CGPBWM  sky130_fd_pr__cap_mim_m3_1_CGPBWM_47
timestamp 1654583101
transform 1 0 35026 0 1 25098
box -1031 -980 975 980
use sky130_fd_pr__cap_mim_m3_1_TABSMU  sky130_fd_pr__cap_mim_m3_1_TABSMU_0
timestamp 1654583101
transform 1 0 41148 0 -1 63799
box -1310 -1260 1210 1260
use sky130_fd_pr__cap_mim_m3_1_TABSMU  sky130_fd_pr__cap_mim_m3_1_TABSMU_1
timestamp 1654583101
transform 1 0 41148 0 -1 60389
box -1310 -1260 1210 1260
use sky130_fd_pr__nfet_01v8_CFEPS5  sky130_fd_pr__nfet_01v8_CFEPS5_0
timestamp 1654583101
transform 1 0 25574 0 -1 63011
box -301 -264 301 266
use sky130_fd_pr__pfet_01v8_hvt_XAYTAL  sky130_fd_pr__pfet_01v8_hvt_XAYTAL_0
timestamp 1654583101
transform 1 0 25574 0 1 62412
box -311 -319 311 319
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_0
timestamp 1654583406
transform 1 0 99516 0 1 68517
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_1
timestamp 1654583406
transform 1 0 99516 0 1 67367
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_2
timestamp 1654583406
transform 1 0 30466 0 1 73168
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_3
timestamp 1654583406
transform 1 0 99516 0 1 64827
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_4
timestamp 1654583406
transform 1 0 99516 0 1 63557
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_0
timestamp 1654583406
transform 1 0 100252 0 1 68517
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_1
timestamp 1654583406
transform 1 0 100252 0 1 67367
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_2
timestamp 1654583406
transform 1 0 100252 0 1 64827
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_3
timestamp 1654583406
transform 1 0 100252 0 1 63557
box -38 -48 2246 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_0
timestamp 1654583406
transform 1 0 102552 0 1 68517
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_1
timestamp 1654583406
transform 1 0 102552 0 1 67367
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_2
timestamp 1654583406
transform 1 0 99056 0 1 68517
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_3
timestamp 1654583406
transform 1 0 99056 0 1 67367
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_4
timestamp 1654583406
transform 1 0 31202 0 1 73168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_5
timestamp 1654583406
transform 1 0 30006 0 1 73168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_6
timestamp 1654583406
transform 1 0 102552 0 1 64827
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_7
timestamp 1654583406
transform 1 0 99056 0 1 64827
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_8
timestamp 1654583406
transform 1 0 102552 0 1 63557
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_9
timestamp 1654583406
transform 1 0 99056 0 1 63557
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  sky130_fd_sc_hd__mux4_1_0
timestamp 1654583101
transform 1 0 97032 0 1 68517
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  sky130_fd_sc_hd__mux4_1_1
timestamp 1654583101
transform 1 0 97032 0 1 67367
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  sky130_fd_sc_hd__mux4_1_2
timestamp 1654583101
transform 1 0 97032 0 1 64827
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  sky130_fd_sc_hd__mux4_1_3
timestamp 1654583101
transform 1 0 97032 0 1 63557
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1654583406
transform 1 0 102460 0 1 68517
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1654583406
transform 1 0 102460 0 1 67367
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1654583406
transform 1 0 99424 0 1 68517
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1654583406
transform 1 0 100160 0 1 68517
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1654583406
transform 1 0 99424 0 1 67367
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1654583406
transform 1 0 100160 0 1 67367
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1654583406
transform 1 0 98964 0 1 68517
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1654583406
transform 1 0 98964 0 1 67367
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_8
timestamp 1654583406
transform 1 0 96940 0 1 68517
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_9
timestamp 1654583406
transform 1 0 96940 0 1 67367
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_10
timestamp 1654583406
transform 1 0 30374 0 1 73168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_11
timestamp 1654583406
transform 1 0 31110 0 1 73168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_12
timestamp 1654583406
transform 1 0 102460 0 1 64827
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_13
timestamp 1654583406
transform 1 0 99424 0 1 64827
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_14
timestamp 1654583406
transform 1 0 100160 0 1 64827
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_15
timestamp 1654583406
transform 1 0 98964 0 1 64827
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_16
timestamp 1654583406
transform 1 0 102460 0 1 63557
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_17
timestamp 1654583406
transform 1 0 99424 0 1 63557
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_18
timestamp 1654583406
transform 1 0 100160 0 1 63557
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_19
timestamp 1654583406
transform 1 0 98964 0 1 63557
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_20
timestamp 1654583406
transform 1 0 96940 0 1 64827
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_21
timestamp 1654583406
transform 1 0 96940 0 1 63557
box -38 -48 130 592
use transmission_gate  transmission_gate_0
timestamp 1654583101
transform -1 0 49476 0 -1 75337
box -216 -51 1283 1063
use transmission_gate  transmission_gate_1
timestamp 1654583101
transform 1 0 58453 0 -1 62969
box -216 -51 1283 1063
use transmission_gate  transmission_gate_2
timestamp 1654583101
transform 0 -1 66967 1 0 58890
box -216 -51 1283 1063
use transmission_gate  transmission_gate_3
timestamp 1654583101
transform 0 1 63955 1 0 58890
box -216 -51 1283 1063
use transmission_gate  transmission_gate_4
timestamp 1654583101
transform 0 -1 62967 1 0 58890
box -216 -51 1283 1063
use transmission_gate  transmission_gate_5
timestamp 1654583101
transform 0 -1 60967 1 0 58890
box -216 -51 1283 1063
use transmission_gate  transmission_gate_6
timestamp 1654583101
transform 1 0 58101 0 -1 61219
box -216 -51 1283 1063
use transmission_gate  transmission_gate_7
timestamp 1654583101
transform 0 1 66116 1 0 46196
box -216 -51 1283 1063
use transmission_gate  transmission_gate_8
timestamp 1654583101
transform -1 0 64042 0 1 47676
box -216 -51 1283 1063
use transmission_gate  transmission_gate_9
timestamp 1654583101
transform 0 -1 60939 1 0 46196
box -216 -51 1283 1063
use transmission_gate  transmission_gate_10
timestamp 1654583101
transform 0 -1 66933 1 0 41855
box -216 -51 1283 1063
use transmission_gate  transmission_gate_11
timestamp 1654583101
transform 0 -1 64933 1 0 41855
box -216 -51 1283 1063
use transmission_gate  transmission_gate_12
timestamp 1654583101
transform 0 -1 62933 1 0 41855
box -216 -51 1283 1063
use transmission_gate  transmission_gate_13
timestamp 1654583101
transform 0 -1 60933 1 0 41855
box -216 -51 1283 1063
use transmission_gate  transmission_gate_14
timestamp 1654583101
transform 0 1 56268 -1 0 42944
box -216 -51 1283 1063
use transmission_gate  transmission_gate_15
timestamp 1654583101
transform 1 0 43546 0 1 51153
box -216 -51 1283 1063
use transmission_gate  transmission_gate_16
timestamp 1654583101
transform 1 0 43546 0 1 49553
box -216 -51 1283 1063
use transmission_gate  transmission_gate_17
timestamp 1654583101
transform 1 0 43546 0 1 47953
box -216 -51 1283 1063
use transmission_gate  transmission_gate_18
timestamp 1654583101
transform 1 0 43546 0 1 46353
box -216 -51 1283 1063
use transmission_gate  transmission_gate_19
timestamp 1654583101
transform 1 0 30487 0 1 48666
box -216 -51 1283 1063
use transmission_gate  transmission_gate_20
timestamp 1654583101
transform 1 0 30487 0 1 41123
box -216 -51 1283 1063
use transmission_gate  transmission_gate_21
timestamp 1654583101
transform -1 0 55193 0 -1 39544
box -216 -51 1283 1063
use transmission_gate  transmission_gate_22
timestamp 1654583101
transform 1 0 51023 0 -1 38548
box -216 -51 1283 1063
use transmission_gate  transmission_gate_23
timestamp 1654583101
transform 0 1 50863 1 0 32376
box -216 -51 1283 1063
use transmission_gate  transmission_gate_24
timestamp 1654583101
transform 0 1 50863 -1 0 36013
box -216 -51 1283 1063
use transmission_gate  transmission_gate_25
timestamp 1654583101
transform 1 0 54127 0 1 33017
box -216 -51 1283 1063
use transmission_gate  transmission_gate_26
timestamp 1654583101
transform 1 0 54127 0 1 34617
box -216 -51 1283 1063
use transmission_gate  transmission_gate_27
timestamp 1654583101
transform 1 0 54127 0 1 36217
box -216 -51 1283 1063
use transmission_gate  transmission_gate_28
timestamp 1654583101
transform -1 0 55191 0 -1 30132
box -216 -51 1283 1063
use transmission_gate  transmission_gate_29
timestamp 1654583101
transform 1 0 51023 0 1 29891
box -216 -51 1283 1063
use transmission_gate  transmission_gate_30
timestamp 1654583101
transform 1 0 54127 0 1 31417
box -216 -51 1283 1063
use transmission_gate  transmission_gate_31
timestamp 1654583101
transform 1 0 30419 0 1 37649
box -216 -51 1283 1063
use transmission_gate  transmission_gate_32
timestamp 1654583101
transform 1 0 30419 0 1 29881
box -216 -51 1283 1063
<< labels >>
flabel metal3 s 119 49049 119 49049 1 FreeSans 20000 0 0 0 ip
port 1 nsew
flabel metal3 s 88 41514 88 41514 1 FreeSans 20000 0 0 0 in
port 2 nsew
flabel metal3 s 228 61469 228 61469 1 FreeSans 20000 0 0 0 op
port 3 nsew
flabel metal3 s 137 74067 137 74067 1 FreeSans 20000 0 0 0 rst_n
port 4 nsew
flabel metal3 s 40231 114276 40231 114276 1 FreeSans 20000 0 0 0 a_probe_1
port 5 nsew
flabel metal3 s 68195 114299 68195 114299 1 FreeSans 20000 0 0 0 i_bias_2
port 6 nsew
flabel metal3 s 80129 114286 80129 114286 1 FreeSans 20000 0 0 0 clk
port 7 nsew
flabel metal3 s 119812 100090 119812 100090 1 FreeSans 20000 0 0 0 a_mod_grp_ctrl_1
port 8 nsew
flabel metal3 s 119870 92728 119870 92728 1 FreeSans 20000 0 0 0 a_mod_grp_ctrl_0
port 9 nsew
flabel metal3 s 119870 85288 119870 85288 1 FreeSans 20000 0 0 0 debug
port 10 nsew
flabel metal3 s 119887 79244 119887 79244 1 FreeSans 20000 0 0 0 d_clk_grp_1_ctrl_0
port 11 nsew
flabel metal3 s 119877 75014 119877 75014 1 FreeSans 20000 0 0 0 d_clk_grp_1_ctrl_1
port 12 nsew
flabel metal3 s 119832 71272 119832 71272 1 FreeSans 20000 0 0 0 d_probe_0
port 13 nsew
flabel metal3 s 119824 67682 119824 67682 1 FreeSans 20000 0 0 0 d_probe_1
port 14 nsew
flabel metal3 s 119849 57563 119849 57563 1 FreeSans 20000 0 0 0 d_probe_2
port 15 nsew
flabel metal3 s 119915 54345 119915 54345 1 FreeSans 20000 0 0 0 d_probe_3
port 16 nsew
flabel metal3 s 119780 64273 119780 64273 1 FreeSans 20000 0 0 0 d_clk_grp_2_ctrl_0
port 17 nsew
flabel metal3 s 119905 61017 119905 61017 1 FreeSans 20000 0 0 0 d_clk_grp_2_ctrl_1
port 18 nsew
flabel metal3 s 119863 46658 119863 46658 1 FreeSans 20000 0 0 0 a_probe_0
port 19 nsew
flabel metal3 s 119904 29715 119904 29715 1 FreeSans 20000 0 0 0 a_probe_2
port 20 nsew
flabel metal3 s 119819 22781 119819 22781 1 FreeSans 20000 0 0 0 a_probe_3
port 21 nsew
flabel metal3 s 56096 120 56096 120 1 FreeSans 20000 0 0 0 i_bias_1
port 22 nsew
flabel metal5 s 3002 114114 3002 114114 1 FreeSans 20000 0 0 0 VDD
port 23 nsew
flabel metal5 s 7042 114074 7042 114074 1 FreeSans 20000 0 0 0 VSS
port 24 nsew
flabel metal5 s 112994 114160 112994 114160 1 FreeSans 20000 0 0 0 VDD
port 23 nsew
flabel metal5 s 117008 114116 117008 114116 1 FreeSans 20000 0 0 0 VSS
port 24 nsew
flabel metal5 s 2992 384 2992 384 1 FreeSans 20000 0 0 0 VDD
port 23 nsew
flabel metal5 s 6986 384 6986 384 1 FreeSans 20000 0 0 0 VSS
port 24 nsew
flabel metal5 s 113022 388 113022 388 1 FreeSans 20000 0 0 0 VDD
port 23 nsew
flabel metal5 s 117006 514 117006 514 1 FreeSans 20000 0 0 0 VSS
port 24 nsew
<< end >>
