* NGSPICE file created from transmission_gate.ext - technology: sky130A

.subckt pmos_tgate a_n416_n136# a_352_n136# a_n128_n136# a_n224_n136# a_64_n136# a_160_n136#
+ a_n320_n136# w_n646_n356# a_n32_n136# a_n508_n136# a_448_n136# a_n512_n234# a_256_n136#
+ VSUBS
X0 a_n224_n136# a_n512_n234# a_n320_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X1 a_352_n136# a_n512_n234# a_256_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X2 a_n128_n136# a_n512_n234# a_n224_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X3 a_256_n136# a_n512_n234# a_160_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X4 a_n416_n136# a_n512_n234# a_n508_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.216e+11p ps=3.34e+06u w=1.36e+06u l=150000u
X5 a_n320_n136# a_n512_n234# a_n416_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X6 a_n32_n136# a_n512_n234# a_n128_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X7 a_448_n136# a_n512_n234# a_352_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.216e+11p pd=3.34e+06u as=0p ps=0u w=1.36e+06u l=150000u
X8 a_64_n136# a_n512_n234# a_n32_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X9 a_160_n136# a_n512_n234# a_64_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
C0 a_n320_n136# a_n512_n234# 0.03fF
C1 a_448_n136# a_n224_n136# 0.03fF
C2 a_160_n136# a_n128_n136# 0.07fF
C3 a_256_n136# a_64_n136# 0.12fF
C4 a_160_n136# a_n224_n136# 0.05fF
C5 a_352_n136# a_n320_n136# 0.03fF
C6 a_256_n136# a_n32_n136# 0.07fF
C7 a_64_n136# w_n646_n356# 0.05fF
C8 a_n32_n136# w_n646_n356# 0.05fF
C9 a_256_n136# w_n646_n356# 0.06fF
C10 a_64_n136# a_n512_n234# 0.03fF
C11 a_n32_n136# a_n512_n234# 0.03fF
C12 a_352_n136# a_64_n136# 0.07fF
C13 a_352_n136# a_n32_n136# 0.05fF
C14 a_256_n136# a_n512_n234# 0.03fF
C15 a_256_n136# a_352_n136# 0.33fF
C16 a_n512_n234# w_n646_n356# 1.47fF
C17 a_160_n136# a_448_n136# 0.07fF
C18 a_n320_n136# a_n508_n136# 0.12fF
C19 a_n320_n136# a_n416_n136# 0.33fF
C20 a_352_n136# w_n646_n356# 0.08fF
C21 a_352_n136# a_n512_n234# 0.03fF
C22 a_n128_n136# a_n320_n136# 0.12fF
C23 a_64_n136# a_n508_n136# 0.03fF
C24 a_64_n136# a_n416_n136# 0.04fF
C25 a_n508_n136# a_n32_n136# 0.04fF
C26 a_n320_n136# a_n224_n136# 0.33fF
C27 a_n416_n136# a_n32_n136# 0.05fF
C28 a_256_n136# a_n508_n136# 0.02fF
C29 a_256_n136# a_n416_n136# 0.03fF
C30 a_n508_n136# w_n646_n356# 0.13fF
C31 a_n416_n136# w_n646_n356# 0.08fF
C32 a_64_n136# a_n128_n136# 0.12fF
C33 a_64_n136# a_n224_n136# 0.07fF
C34 a_n128_n136# a_n32_n136# 0.33fF
C35 a_n32_n136# a_n224_n136# 0.12fF
C36 a_n508_n136# a_n512_n234# 0.03fF
C37 a_n416_n136# a_n512_n234# 0.03fF
C38 a_256_n136# a_n128_n136# 0.05fF
C39 a_352_n136# a_n508_n136# 0.02fF
C40 a_352_n136# a_n416_n136# 0.02fF
C41 a_256_n136# a_n224_n136# 0.04fF
C42 a_448_n136# a_n320_n136# 0.02fF
C43 a_n128_n136# w_n646_n356# 0.05fF
C44 a_160_n136# a_n320_n136# 0.04fF
C45 a_n224_n136# w_n646_n356# 0.06fF
C46 a_n128_n136# a_n512_n234# 0.03fF
C47 a_n224_n136# a_n512_n234# 0.03fF
C48 a_352_n136# a_n128_n136# 0.04fF
C49 a_352_n136# a_n224_n136# 0.03fF
C50 a_448_n136# a_64_n136# 0.05fF
C51 a_448_n136# a_n32_n136# 0.04fF
C52 a_160_n136# a_64_n136# 0.33fF
C53 a_160_n136# a_n32_n136# 0.12fF
C54 a_256_n136# a_448_n136# 0.12fF
C55 a_n508_n136# a_n416_n136# 0.33fF
C56 a_256_n136# a_160_n136# 0.33fF
C57 a_448_n136# w_n646_n356# 0.13fF
C58 a_160_n136# w_n646_n356# 0.06fF
C59 a_448_n136# a_n512_n234# 0.03fF
C60 a_160_n136# a_n512_n234# 0.03fF
C61 a_n128_n136# a_n508_n136# 0.05fF
C62 a_n128_n136# a_n416_n136# 0.07fF
C63 a_448_n136# a_352_n136# 0.33fF
C64 a_n508_n136# a_n224_n136# 0.07fF
C65 a_n416_n136# a_n224_n136# 0.12fF
C66 a_160_n136# a_352_n136# 0.12fF
C67 a_n128_n136# a_n224_n136# 0.33fF
C68 a_64_n136# a_n320_n136# 0.05fF
C69 a_n320_n136# a_n32_n136# 0.07fF
C70 a_448_n136# a_n508_n136# 0.02fF
C71 a_448_n136# a_n416_n136# 0.02fF
C72 a_160_n136# a_n508_n136# 0.03fF
C73 a_160_n136# a_n416_n136# 0.03fF
C74 a_256_n136# a_n320_n136# 0.03fF
C75 a_n320_n136# w_n646_n356# 0.06fF
C76 a_64_n136# a_n32_n136# 0.33fF
C77 a_448_n136# a_n128_n136# 0.03fF
C78 w_n646_n356# VSUBS 2.52fF
.ends

.subckt nmos_tgate a_256_n52# a_n32_n52# a_n224_n52# a_448_n52# a_n416_n52# a_160_n52#
+ a_n610_n226# a_n128_n52# a_352_n52# a_n320_n52# a_n508_n52# a_n512_n149# a_64_n52#
X0 a_n32_n52# a_n512_n149# a_n128_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X1 a_n416_n52# a_n512_n149# a_n508_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.612e+11p ps=1.66e+06u w=520000u l=150000u
X2 a_n224_n52# a_n512_n149# a_n320_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X3 a_n128_n52# a_n512_n149# a_n224_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4 a_n320_n52# a_n512_n149# a_n416_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X5 a_160_n52# a_n512_n149# a_64_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X6 a_352_n52# a_n512_n149# a_256_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X7 a_256_n52# a_n512_n149# a_160_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X8 a_448_n52# a_n512_n149# a_352_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.612e+11p pd=1.66e+06u as=0p ps=0u w=520000u l=150000u
X9 a_64_n52# a_n512_n149# a_n32_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
C0 a_256_n52# a_n320_n52# 0.01fF
C1 a_n32_n52# a_64_n52# 0.13fF
C2 a_n320_n52# a_448_n52# 0.01fF
C3 a_160_n52# a_n224_n52# 0.02fF
C4 a_n512_n149# a_64_n52# 0.03fF
C5 a_n224_n52# a_352_n52# 0.01fF
C6 a_256_n52# a_n224_n52# 0.02fF
C7 a_n224_n52# a_448_n52# 0.01fF
C8 a_n508_n52# a_n416_n52# 0.13fF
C9 a_160_n52# a_64_n52# 0.13fF
C10 a_n320_n52# a_n224_n52# 0.13fF
C11 a_64_n52# a_352_n52# 0.03fF
C12 a_256_n52# a_64_n52# 0.05fF
C13 a_n416_n52# a_n128_n52# 0.03fF
C14 a_64_n52# a_448_n52# 0.02fF
C15 a_n32_n52# a_n416_n52# 0.02fF
C16 a_n508_n52# a_n128_n52# 0.02fF
C17 a_n320_n52# a_64_n52# 0.02fF
C18 a_n32_n52# a_n508_n52# 0.02fF
C19 a_n512_n149# a_n416_n52# 0.03fF
C20 a_n512_n149# a_n508_n52# 0.03fF
C21 a_n32_n52# a_n128_n52# 0.13fF
C22 a_n224_n52# a_64_n52# 0.03fF
C23 a_160_n52# a_n416_n52# 0.01fF
C24 a_n416_n52# a_352_n52# 0.01fF
C25 a_n512_n149# a_n128_n52# 0.03fF
C26 a_160_n52# a_n508_n52# 0.01fF
C27 a_256_n52# a_n416_n52# 0.01fF
C28 a_n32_n52# a_n512_n149# 0.03fF
C29 a_n508_n52# a_352_n52# 0.01fF
C30 a_256_n52# a_n508_n52# 0.01fF
C31 a_n416_n52# a_448_n52# 0.01fF
C32 a_160_n52# a_n128_n52# 0.03fF
C33 a_n508_n52# a_448_n52# 0.01fF
C34 a_n320_n52# a_n416_n52# 0.13fF
C35 a_160_n52# a_n32_n52# 0.05fF
C36 a_n128_n52# a_352_n52# 0.02fF
C37 a_256_n52# a_n128_n52# 0.02fF
C38 a_n320_n52# a_n508_n52# 0.05fF
C39 a_n32_n52# a_352_n52# 0.02fF
C40 a_256_n52# a_n32_n52# 0.03fF
C41 a_n128_n52# a_448_n52# 0.01fF
C42 a_160_n52# a_n512_n149# 0.03fF
C43 a_n224_n52# a_n416_n52# 0.05fF
C44 a_n32_n52# a_448_n52# 0.02fF
C45 a_n512_n149# a_352_n52# 0.03fF
C46 a_n320_n52# a_n128_n52# 0.05fF
C47 a_256_n52# a_n512_n149# 0.03fF
C48 a_n224_n52# a_n508_n52# 0.03fF
C49 a_n320_n52# a_n32_n52# 0.03fF
C50 a_n512_n149# a_448_n52# 0.03fF
C51 a_160_n52# a_352_n52# 0.05fF
C52 a_n416_n52# a_64_n52# 0.02fF
C53 a_160_n52# a_256_n52# 0.13fF
C54 a_n224_n52# a_n128_n52# 0.13fF
C55 a_n320_n52# a_n512_n149# 0.03fF
C56 a_n508_n52# a_64_n52# 0.01fF
C57 a_256_n52# a_352_n52# 0.13fF
C58 a_n32_n52# a_n224_n52# 0.05fF
C59 a_160_n52# a_448_n52# 0.03fF
C60 a_352_n52# a_448_n52# 0.13fF
C61 a_256_n52# a_448_n52# 0.05fF
C62 a_160_n52# a_n320_n52# 0.02fF
C63 a_n224_n52# a_n512_n149# 0.03fF
C64 a_64_n52# a_n128_n52# 0.05fF
C65 a_n320_n52# a_352_n52# 0.01fF
C66 a_448_n52# a_n610_n226# 0.07fF
C67 a_352_n52# a_n610_n226# 0.05fF
C68 a_256_n52# a_n610_n226# 0.04fF
C69 a_160_n52# a_n610_n226# 0.04fF
C70 a_64_n52# a_n610_n226# 0.04fF
C71 a_n32_n52# a_n610_n226# 0.04fF
C72 a_n128_n52# a_n610_n226# 0.04fF
C73 a_n224_n52# a_n610_n226# 0.04fF
C74 a_n320_n52# a_n610_n226# 0.04fF
C75 a_n416_n52# a_n610_n226# 0.05fF
C76 a_n508_n52# a_n610_n226# 0.07fF
C77 a_n512_n149# a_n610_n226# 1.83fF
.ends

.subckt transmission_gate in out en en_b VDD VSS
Xpmos_tgate_0 in in out in out in out VDD in out out en_b out VSS pmos_tgate
Xnmos_tgate_0 out in in out in in VSS out in out out en out nmos_tgate
C0 out en 0.01fF
C1 out VDD 0.29fF
C2 out en_b 0.01fF
C3 out in 0.77fF
C4 en VDD 0.12fF
C5 en_b en 0.07fF
C6 en in 0.13fF
C7 en_b VDD -0.11fF
C8 in VDD 0.70fF
C9 en_b in 0.15fF
C10 en VSS 1.70fF
C11 out VSS 0.57fF
C12 in VSS 1.13fF
C13 en_b VSS 0.09fF
C14 VDD VSS 3.16fF
.ends

