magic
tech sky130A
magscale 1 2
timestamp 1654599767
<< error_p >>
rect -559 192 -501 198
rect -135 192 -77 198
rect 289 192 347 198
rect 713 192 771 198
rect -559 158 -547 192
rect -135 158 -123 192
rect 289 158 301 192
rect 713 158 725 192
rect -559 152 -501 158
rect -135 152 -77 158
rect 289 152 347 158
rect 713 152 771 158
rect -771 -158 -713 -152
rect -347 -158 -289 -152
rect 77 -158 135 -152
rect 501 -158 559 -152
rect -771 -192 -759 -158
rect -347 -192 -335 -158
rect 77 -192 89 -158
rect 501 -192 513 -158
rect -771 -198 -713 -192
rect -347 -198 -289 -192
rect 77 -198 135 -192
rect 501 -198 559 -192
<< nmoslvt >>
rect -762 -120 -722 120
rect -550 -120 -510 120
rect -338 -120 -298 120
rect -126 -120 -86 120
rect 86 -120 126 120
rect 298 -120 338 120
rect 510 -120 550 120
rect 722 -120 762 120
<< ndiff >>
rect -820 108 -762 120
rect -820 -108 -808 108
rect -774 -108 -762 108
rect -820 -120 -762 -108
rect -722 108 -664 120
rect -722 -108 -710 108
rect -676 -108 -664 108
rect -722 -120 -664 -108
rect -608 108 -550 120
rect -608 -108 -596 108
rect -562 -108 -550 108
rect -608 -120 -550 -108
rect -510 108 -452 120
rect -510 -108 -498 108
rect -464 -108 -452 108
rect -510 -120 -452 -108
rect -396 108 -338 120
rect -396 -108 -384 108
rect -350 -108 -338 108
rect -396 -120 -338 -108
rect -298 108 -240 120
rect -298 -108 -286 108
rect -252 -108 -240 108
rect -298 -120 -240 -108
rect -184 108 -126 120
rect -184 -108 -172 108
rect -138 -108 -126 108
rect -184 -120 -126 -108
rect -86 108 -28 120
rect -86 -108 -74 108
rect -40 -108 -28 108
rect -86 -120 -28 -108
rect 28 108 86 120
rect 28 -108 40 108
rect 74 -108 86 108
rect 28 -120 86 -108
rect 126 108 184 120
rect 126 -108 138 108
rect 172 -108 184 108
rect 126 -120 184 -108
rect 240 108 298 120
rect 240 -108 252 108
rect 286 -108 298 108
rect 240 -120 298 -108
rect 338 108 396 120
rect 338 -108 350 108
rect 384 -108 396 108
rect 338 -120 396 -108
rect 452 108 510 120
rect 452 -108 464 108
rect 498 -108 510 108
rect 452 -120 510 -108
rect 550 108 608 120
rect 550 -108 562 108
rect 596 -108 608 108
rect 550 -120 608 -108
rect 664 108 722 120
rect 664 -108 676 108
rect 710 -108 722 108
rect 664 -120 722 -108
rect 762 108 820 120
rect 762 -108 774 108
rect 808 -108 820 108
rect 762 -120 820 -108
<< ndiffc >>
rect -808 -108 -774 108
rect -710 -108 -676 108
rect -596 -108 -562 108
rect -498 -108 -464 108
rect -384 -108 -350 108
rect -286 -108 -252 108
rect -172 -108 -138 108
rect -74 -108 -40 108
rect 40 -108 74 108
rect 138 -108 172 108
rect 252 -108 286 108
rect 350 -108 384 108
rect 464 -108 498 108
rect 562 -108 596 108
rect 676 -108 710 108
rect 774 -108 808 108
<< poly >>
rect -563 192 -497 208
rect -563 158 -547 192
rect -513 158 -497 192
rect -762 120 -722 146
rect -563 142 -497 158
rect -139 192 -73 208
rect -139 158 -123 192
rect -89 158 -73 192
rect -550 120 -510 142
rect -338 120 -298 146
rect -139 142 -73 158
rect 285 192 351 208
rect 285 158 301 192
rect 335 158 351 192
rect -126 120 -86 142
rect 86 120 126 146
rect 285 142 351 158
rect 709 192 775 208
rect 709 158 725 192
rect 759 158 775 192
rect 298 120 338 142
rect 510 120 550 146
rect 709 142 775 158
rect 722 120 762 142
rect -762 -142 -722 -120
rect -775 -158 -709 -142
rect -550 -146 -510 -120
rect -338 -142 -298 -120
rect -775 -192 -759 -158
rect -725 -192 -709 -158
rect -775 -208 -709 -192
rect -351 -158 -285 -142
rect -126 -146 -86 -120
rect 86 -142 126 -120
rect -351 -192 -335 -158
rect -301 -192 -285 -158
rect -351 -208 -285 -192
rect 73 -158 139 -142
rect 298 -146 338 -120
rect 510 -142 550 -120
rect 73 -192 89 -158
rect 123 -192 139 -158
rect 73 -208 139 -192
rect 497 -158 563 -142
rect 722 -146 762 -120
rect 497 -192 513 -158
rect 547 -192 563 -158
rect 497 -208 563 -192
<< polycont >>
rect -547 158 -513 192
rect -123 158 -89 192
rect 301 158 335 192
rect 725 158 759 192
rect -759 -192 -725 -158
rect -335 -192 -301 -158
rect 89 -192 123 -158
rect 513 -192 547 -158
<< locali >>
rect -563 158 -547 192
rect -513 158 -497 192
rect -139 158 -123 192
rect -89 158 -73 192
rect 285 158 301 192
rect 335 158 351 192
rect 709 158 725 192
rect 759 158 775 192
rect -808 108 -774 124
rect -808 -124 -774 -108
rect -710 108 -676 124
rect -710 -124 -676 -108
rect -596 108 -562 124
rect -596 -124 -562 -108
rect -498 108 -464 124
rect -498 -124 -464 -108
rect -384 108 -350 124
rect -384 -124 -350 -108
rect -286 108 -252 124
rect -286 -124 -252 -108
rect -172 108 -138 124
rect -172 -124 -138 -108
rect -74 108 -40 124
rect -74 -124 -40 -108
rect 40 108 74 124
rect 40 -124 74 -108
rect 138 108 172 124
rect 138 -124 172 -108
rect 252 108 286 124
rect 252 -124 286 -108
rect 350 108 384 124
rect 350 -124 384 -108
rect 464 108 498 124
rect 464 -124 498 -108
rect 562 108 596 124
rect 562 -124 596 -108
rect 676 108 710 124
rect 676 -124 710 -108
rect 774 108 808 124
rect 774 -124 808 -108
rect -775 -192 -759 -158
rect -725 -192 -709 -158
rect -351 -192 -335 -158
rect -301 -192 -285 -158
rect 73 -192 89 -158
rect 123 -192 139 -158
rect 497 -192 513 -158
rect 547 -192 563 -158
<< viali >>
rect -547 158 -513 192
rect -123 158 -89 192
rect 301 158 335 192
rect 725 158 759 192
rect -759 -192 -725 -158
rect -335 -192 -301 -158
rect 89 -192 123 -158
rect 513 -192 547 -158
<< metal1 >>
rect -559 192 -501 198
rect -559 158 -547 192
rect -513 158 -501 192
rect -559 152 -501 158
rect -135 192 -77 198
rect -135 158 -123 192
rect -89 158 -77 192
rect -135 152 -77 158
rect 289 192 347 198
rect 289 158 301 192
rect 335 158 347 192
rect 289 152 347 158
rect 713 192 771 198
rect 713 158 725 192
rect 759 158 771 192
rect 713 152 771 158
rect -771 -158 -713 -152
rect -771 -192 -759 -158
rect -725 -192 -713 -158
rect -771 -198 -713 -192
rect -347 -158 -289 -152
rect -347 -192 -335 -158
rect -301 -192 -289 -158
rect -347 -198 -289 -192
rect 77 -158 135 -152
rect 77 -192 89 -158
rect 123 -192 135 -158
rect 77 -198 135 -192
rect 501 -158 559 -152
rect 501 -192 513 -158
rect 547 -192 559 -158
rect 501 -198 559 -192
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1.2 l 0.2 m 1 nf 8 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 0 viadrn 0 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
