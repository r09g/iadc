magic
tech sky130A
magscale 1 2
timestamp 1653911004
<< error_p >>
rect -1530 581 -1472 587
rect -1372 581 -1314 587
rect -1214 581 -1156 587
rect -1056 581 -998 587
rect -898 581 -840 587
rect -740 581 -682 587
rect -582 581 -524 587
rect -424 581 -366 587
rect -266 581 -208 587
rect -108 581 -50 587
rect 50 581 108 587
rect 208 581 266 587
rect 366 581 424 587
rect 524 581 582 587
rect 682 581 740 587
rect 840 581 898 587
rect 998 581 1056 587
rect 1156 581 1214 587
rect 1314 581 1372 587
rect 1472 581 1530 587
rect -1530 547 -1518 581
rect -1372 547 -1360 581
rect -1214 547 -1202 581
rect -1056 547 -1044 581
rect -898 547 -886 581
rect -740 547 -728 581
rect -582 547 -570 581
rect -424 547 -412 581
rect -266 547 -254 581
rect -108 547 -96 581
rect 50 547 62 581
rect 208 547 220 581
rect 366 547 378 581
rect 524 547 536 581
rect 682 547 694 581
rect 840 547 852 581
rect 998 547 1010 581
rect 1156 547 1168 581
rect 1314 547 1326 581
rect 1472 547 1484 581
rect -1530 541 -1472 547
rect -1372 541 -1314 547
rect -1214 541 -1156 547
rect -1056 541 -998 547
rect -898 541 -840 547
rect -740 541 -682 547
rect -582 541 -524 547
rect -424 541 -366 547
rect -266 541 -208 547
rect -108 541 -50 547
rect 50 541 108 547
rect 208 541 266 547
rect 366 541 424 547
rect 524 541 582 547
rect 682 541 740 547
rect 840 541 898 547
rect 998 541 1056 547
rect 1156 541 1214 547
rect 1314 541 1372 547
rect 1472 541 1530 547
rect -1530 -547 -1472 -541
rect -1372 -547 -1314 -541
rect -1214 -547 -1156 -541
rect -1056 -547 -998 -541
rect -898 -547 -840 -541
rect -740 -547 -682 -541
rect -582 -547 -524 -541
rect -424 -547 -366 -541
rect -266 -547 -208 -541
rect -108 -547 -50 -541
rect 50 -547 108 -541
rect 208 -547 266 -541
rect 366 -547 424 -541
rect 524 -547 582 -541
rect 682 -547 740 -541
rect 840 -547 898 -541
rect 998 -547 1056 -541
rect 1156 -547 1214 -541
rect 1314 -547 1372 -541
rect 1472 -547 1530 -541
rect -1530 -581 -1518 -547
rect -1372 -581 -1360 -547
rect -1214 -581 -1202 -547
rect -1056 -581 -1044 -547
rect -898 -581 -886 -547
rect -740 -581 -728 -547
rect -582 -581 -570 -547
rect -424 -581 -412 -547
rect -266 -581 -254 -547
rect -108 -581 -96 -547
rect 50 -581 62 -547
rect 208 -581 220 -547
rect 366 -581 378 -547
rect 524 -581 536 -547
rect 682 -581 694 -547
rect 840 -581 852 -547
rect 998 -581 1010 -547
rect 1156 -581 1168 -547
rect 1314 -581 1326 -547
rect 1472 -581 1484 -547
rect -1530 -587 -1472 -581
rect -1372 -587 -1314 -581
rect -1214 -587 -1156 -581
rect -1056 -587 -998 -581
rect -898 -587 -840 -581
rect -740 -587 -682 -581
rect -582 -587 -524 -581
rect -424 -587 -366 -581
rect -266 -587 -208 -581
rect -108 -587 -50 -581
rect 50 -587 108 -581
rect 208 -587 266 -581
rect 366 -587 424 -581
rect 524 -587 582 -581
rect 682 -587 740 -581
rect 840 -587 898 -581
rect 998 -587 1056 -581
rect 1156 -587 1214 -581
rect 1314 -587 1372 -581
rect 1472 -587 1530 -581
<< nwell >>
rect -1809 -797 1809 797
<< mvpmos >>
rect -1551 -500 -1451 500
rect -1393 -500 -1293 500
rect -1235 -500 -1135 500
rect -1077 -500 -977 500
rect -919 -500 -819 500
rect -761 -500 -661 500
rect -603 -500 -503 500
rect -445 -500 -345 500
rect -287 -500 -187 500
rect -129 -500 -29 500
rect 29 -500 129 500
rect 187 -500 287 500
rect 345 -500 445 500
rect 503 -500 603 500
rect 661 -500 761 500
rect 819 -500 919 500
rect 977 -500 1077 500
rect 1135 -500 1235 500
rect 1293 -500 1393 500
rect 1451 -500 1551 500
<< mvpdiff >>
rect -1609 488 -1551 500
rect -1609 -488 -1597 488
rect -1563 -488 -1551 488
rect -1609 -500 -1551 -488
rect -1451 488 -1393 500
rect -1451 -488 -1439 488
rect -1405 -488 -1393 488
rect -1451 -500 -1393 -488
rect -1293 488 -1235 500
rect -1293 -488 -1281 488
rect -1247 -488 -1235 488
rect -1293 -500 -1235 -488
rect -1135 488 -1077 500
rect -1135 -488 -1123 488
rect -1089 -488 -1077 488
rect -1135 -500 -1077 -488
rect -977 488 -919 500
rect -977 -488 -965 488
rect -931 -488 -919 488
rect -977 -500 -919 -488
rect -819 488 -761 500
rect -819 -488 -807 488
rect -773 -488 -761 488
rect -819 -500 -761 -488
rect -661 488 -603 500
rect -661 -488 -649 488
rect -615 -488 -603 488
rect -661 -500 -603 -488
rect -503 488 -445 500
rect -503 -488 -491 488
rect -457 -488 -445 488
rect -503 -500 -445 -488
rect -345 488 -287 500
rect -345 -488 -333 488
rect -299 -488 -287 488
rect -345 -500 -287 -488
rect -187 488 -129 500
rect -187 -488 -175 488
rect -141 -488 -129 488
rect -187 -500 -129 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 129 488 187 500
rect 129 -488 141 488
rect 175 -488 187 488
rect 129 -500 187 -488
rect 287 488 345 500
rect 287 -488 299 488
rect 333 -488 345 488
rect 287 -500 345 -488
rect 445 488 503 500
rect 445 -488 457 488
rect 491 -488 503 488
rect 445 -500 503 -488
rect 603 488 661 500
rect 603 -488 615 488
rect 649 -488 661 488
rect 603 -500 661 -488
rect 761 488 819 500
rect 761 -488 773 488
rect 807 -488 819 488
rect 761 -500 819 -488
rect 919 488 977 500
rect 919 -488 931 488
rect 965 -488 977 488
rect 919 -500 977 -488
rect 1077 488 1135 500
rect 1077 -488 1089 488
rect 1123 -488 1135 488
rect 1077 -500 1135 -488
rect 1235 488 1293 500
rect 1235 -488 1247 488
rect 1281 -488 1293 488
rect 1235 -500 1293 -488
rect 1393 488 1451 500
rect 1393 -488 1405 488
rect 1439 -488 1451 488
rect 1393 -500 1451 -488
rect 1551 488 1609 500
rect 1551 -488 1563 488
rect 1597 -488 1609 488
rect 1551 -500 1609 -488
<< mvpdiffc >>
rect -1597 -488 -1563 488
rect -1439 -488 -1405 488
rect -1281 -488 -1247 488
rect -1123 -488 -1089 488
rect -965 -488 -931 488
rect -807 -488 -773 488
rect -649 -488 -615 488
rect -491 -488 -457 488
rect -333 -488 -299 488
rect -175 -488 -141 488
rect -17 -488 17 488
rect 141 -488 175 488
rect 299 -488 333 488
rect 457 -488 491 488
rect 615 -488 649 488
rect 773 -488 807 488
rect 931 -488 965 488
rect 1089 -488 1123 488
rect 1247 -488 1281 488
rect 1405 -488 1439 488
rect 1563 -488 1597 488
<< mvnsubdiff >>
rect -1743 719 1743 731
rect -1743 685 -1635 719
rect 1635 685 1743 719
rect -1743 673 1743 685
rect -1743 623 -1685 673
rect -1743 -623 -1731 623
rect -1697 -623 -1685 623
rect 1685 623 1743 673
rect -1743 -673 -1685 -623
rect 1685 -623 1697 623
rect 1731 -623 1743 623
rect 1685 -673 1743 -623
rect -1743 -685 1743 -673
rect -1743 -719 -1635 -685
rect 1635 -719 1743 -685
rect -1743 -731 1743 -719
<< mvnsubdiffcont >>
rect -1635 685 1635 719
rect -1731 -623 -1697 623
rect 1697 -623 1731 623
rect -1635 -719 1635 -685
<< poly >>
rect -1551 581 -1451 597
rect -1551 547 -1535 581
rect -1467 547 -1451 581
rect -1551 500 -1451 547
rect -1393 581 -1293 597
rect -1393 547 -1377 581
rect -1309 547 -1293 581
rect -1393 500 -1293 547
rect -1235 581 -1135 597
rect -1235 547 -1219 581
rect -1151 547 -1135 581
rect -1235 500 -1135 547
rect -1077 581 -977 597
rect -1077 547 -1061 581
rect -993 547 -977 581
rect -1077 500 -977 547
rect -919 581 -819 597
rect -919 547 -903 581
rect -835 547 -819 581
rect -919 500 -819 547
rect -761 581 -661 597
rect -761 547 -745 581
rect -677 547 -661 581
rect -761 500 -661 547
rect -603 581 -503 597
rect -603 547 -587 581
rect -519 547 -503 581
rect -603 500 -503 547
rect -445 581 -345 597
rect -445 547 -429 581
rect -361 547 -345 581
rect -445 500 -345 547
rect -287 581 -187 597
rect -287 547 -271 581
rect -203 547 -187 581
rect -287 500 -187 547
rect -129 581 -29 597
rect -129 547 -113 581
rect -45 547 -29 581
rect -129 500 -29 547
rect 29 581 129 597
rect 29 547 45 581
rect 113 547 129 581
rect 29 500 129 547
rect 187 581 287 597
rect 187 547 203 581
rect 271 547 287 581
rect 187 500 287 547
rect 345 581 445 597
rect 345 547 361 581
rect 429 547 445 581
rect 345 500 445 547
rect 503 581 603 597
rect 503 547 519 581
rect 587 547 603 581
rect 503 500 603 547
rect 661 581 761 597
rect 661 547 677 581
rect 745 547 761 581
rect 661 500 761 547
rect 819 581 919 597
rect 819 547 835 581
rect 903 547 919 581
rect 819 500 919 547
rect 977 581 1077 597
rect 977 547 993 581
rect 1061 547 1077 581
rect 977 500 1077 547
rect 1135 581 1235 597
rect 1135 547 1151 581
rect 1219 547 1235 581
rect 1135 500 1235 547
rect 1293 581 1393 597
rect 1293 547 1309 581
rect 1377 547 1393 581
rect 1293 500 1393 547
rect 1451 581 1551 597
rect 1451 547 1467 581
rect 1535 547 1551 581
rect 1451 500 1551 547
rect -1551 -547 -1451 -500
rect -1551 -581 -1535 -547
rect -1467 -581 -1451 -547
rect -1551 -597 -1451 -581
rect -1393 -547 -1293 -500
rect -1393 -581 -1377 -547
rect -1309 -581 -1293 -547
rect -1393 -597 -1293 -581
rect -1235 -547 -1135 -500
rect -1235 -581 -1219 -547
rect -1151 -581 -1135 -547
rect -1235 -597 -1135 -581
rect -1077 -547 -977 -500
rect -1077 -581 -1061 -547
rect -993 -581 -977 -547
rect -1077 -597 -977 -581
rect -919 -547 -819 -500
rect -919 -581 -903 -547
rect -835 -581 -819 -547
rect -919 -597 -819 -581
rect -761 -547 -661 -500
rect -761 -581 -745 -547
rect -677 -581 -661 -547
rect -761 -597 -661 -581
rect -603 -547 -503 -500
rect -603 -581 -587 -547
rect -519 -581 -503 -547
rect -603 -597 -503 -581
rect -445 -547 -345 -500
rect -445 -581 -429 -547
rect -361 -581 -345 -547
rect -445 -597 -345 -581
rect -287 -547 -187 -500
rect -287 -581 -271 -547
rect -203 -581 -187 -547
rect -287 -597 -187 -581
rect -129 -547 -29 -500
rect -129 -581 -113 -547
rect -45 -581 -29 -547
rect -129 -597 -29 -581
rect 29 -547 129 -500
rect 29 -581 45 -547
rect 113 -581 129 -547
rect 29 -597 129 -581
rect 187 -547 287 -500
rect 187 -581 203 -547
rect 271 -581 287 -547
rect 187 -597 287 -581
rect 345 -547 445 -500
rect 345 -581 361 -547
rect 429 -581 445 -547
rect 345 -597 445 -581
rect 503 -547 603 -500
rect 503 -581 519 -547
rect 587 -581 603 -547
rect 503 -597 603 -581
rect 661 -547 761 -500
rect 661 -581 677 -547
rect 745 -581 761 -547
rect 661 -597 761 -581
rect 819 -547 919 -500
rect 819 -581 835 -547
rect 903 -581 919 -547
rect 819 -597 919 -581
rect 977 -547 1077 -500
rect 977 -581 993 -547
rect 1061 -581 1077 -547
rect 977 -597 1077 -581
rect 1135 -547 1235 -500
rect 1135 -581 1151 -547
rect 1219 -581 1235 -547
rect 1135 -597 1235 -581
rect 1293 -547 1393 -500
rect 1293 -581 1309 -547
rect 1377 -581 1393 -547
rect 1293 -597 1393 -581
rect 1451 -547 1551 -500
rect 1451 -581 1467 -547
rect 1535 -581 1551 -547
rect 1451 -597 1551 -581
<< polycont >>
rect -1535 547 -1467 581
rect -1377 547 -1309 581
rect -1219 547 -1151 581
rect -1061 547 -993 581
rect -903 547 -835 581
rect -745 547 -677 581
rect -587 547 -519 581
rect -429 547 -361 581
rect -271 547 -203 581
rect -113 547 -45 581
rect 45 547 113 581
rect 203 547 271 581
rect 361 547 429 581
rect 519 547 587 581
rect 677 547 745 581
rect 835 547 903 581
rect 993 547 1061 581
rect 1151 547 1219 581
rect 1309 547 1377 581
rect 1467 547 1535 581
rect -1535 -581 -1467 -547
rect -1377 -581 -1309 -547
rect -1219 -581 -1151 -547
rect -1061 -581 -993 -547
rect -903 -581 -835 -547
rect -745 -581 -677 -547
rect -587 -581 -519 -547
rect -429 -581 -361 -547
rect -271 -581 -203 -547
rect -113 -581 -45 -547
rect 45 -581 113 -547
rect 203 -581 271 -547
rect 361 -581 429 -547
rect 519 -581 587 -547
rect 677 -581 745 -547
rect 835 -581 903 -547
rect 993 -581 1061 -547
rect 1151 -581 1219 -547
rect 1309 -581 1377 -547
rect 1467 -581 1535 -547
<< locali >>
rect -1731 685 -1635 719
rect 1635 685 1731 719
rect -1731 623 -1697 685
rect 1697 623 1731 685
rect -1551 547 -1535 581
rect -1467 547 -1451 581
rect -1393 547 -1377 581
rect -1309 547 -1293 581
rect -1235 547 -1219 581
rect -1151 547 -1135 581
rect -1077 547 -1061 581
rect -993 547 -977 581
rect -919 547 -903 581
rect -835 547 -819 581
rect -761 547 -745 581
rect -677 547 -661 581
rect -603 547 -587 581
rect -519 547 -503 581
rect -445 547 -429 581
rect -361 547 -345 581
rect -287 547 -271 581
rect -203 547 -187 581
rect -129 547 -113 581
rect -45 547 -29 581
rect 29 547 45 581
rect 113 547 129 581
rect 187 547 203 581
rect 271 547 287 581
rect 345 547 361 581
rect 429 547 445 581
rect 503 547 519 581
rect 587 547 603 581
rect 661 547 677 581
rect 745 547 761 581
rect 819 547 835 581
rect 903 547 919 581
rect 977 547 993 581
rect 1061 547 1077 581
rect 1135 547 1151 581
rect 1219 547 1235 581
rect 1293 547 1309 581
rect 1377 547 1393 581
rect 1451 547 1467 581
rect 1535 547 1551 581
rect -1597 488 -1563 504
rect -1597 -504 -1563 -488
rect -1439 488 -1405 504
rect -1439 -504 -1405 -488
rect -1281 488 -1247 504
rect -1281 -504 -1247 -488
rect -1123 488 -1089 504
rect -1123 -504 -1089 -488
rect -965 488 -931 504
rect -965 -504 -931 -488
rect -807 488 -773 504
rect -807 -504 -773 -488
rect -649 488 -615 504
rect -649 -504 -615 -488
rect -491 488 -457 504
rect -491 -504 -457 -488
rect -333 488 -299 504
rect -333 -504 -299 -488
rect -175 488 -141 504
rect -175 -504 -141 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 141 488 175 504
rect 141 -504 175 -488
rect 299 488 333 504
rect 299 -504 333 -488
rect 457 488 491 504
rect 457 -504 491 -488
rect 615 488 649 504
rect 615 -504 649 -488
rect 773 488 807 504
rect 773 -504 807 -488
rect 931 488 965 504
rect 931 -504 965 -488
rect 1089 488 1123 504
rect 1089 -504 1123 -488
rect 1247 488 1281 504
rect 1247 -504 1281 -488
rect 1405 488 1439 504
rect 1405 -504 1439 -488
rect 1563 488 1597 504
rect 1563 -504 1597 -488
rect -1551 -581 -1535 -547
rect -1467 -581 -1451 -547
rect -1393 -581 -1377 -547
rect -1309 -581 -1293 -547
rect -1235 -581 -1219 -547
rect -1151 -581 -1135 -547
rect -1077 -581 -1061 -547
rect -993 -581 -977 -547
rect -919 -581 -903 -547
rect -835 -581 -819 -547
rect -761 -581 -745 -547
rect -677 -581 -661 -547
rect -603 -581 -587 -547
rect -519 -581 -503 -547
rect -445 -581 -429 -547
rect -361 -581 -345 -547
rect -287 -581 -271 -547
rect -203 -581 -187 -547
rect -129 -581 -113 -547
rect -45 -581 -29 -547
rect 29 -581 45 -547
rect 113 -581 129 -547
rect 187 -581 203 -547
rect 271 -581 287 -547
rect 345 -581 361 -547
rect 429 -581 445 -547
rect 503 -581 519 -547
rect 587 -581 603 -547
rect 661 -581 677 -547
rect 745 -581 761 -547
rect 819 -581 835 -547
rect 903 -581 919 -547
rect 977 -581 993 -547
rect 1061 -581 1077 -547
rect 1135 -581 1151 -547
rect 1219 -581 1235 -547
rect 1293 -581 1309 -547
rect 1377 -581 1393 -547
rect 1451 -581 1467 -547
rect 1535 -581 1551 -547
rect -1731 -685 -1697 -623
rect 1697 -685 1731 -623
rect -1731 -719 -1635 -685
rect 1635 -719 1731 -685
<< viali >>
rect -1518 547 -1484 581
rect -1360 547 -1326 581
rect -1202 547 -1168 581
rect -1044 547 -1010 581
rect -886 547 -852 581
rect -728 547 -694 581
rect -570 547 -536 581
rect -412 547 -378 581
rect -254 547 -220 581
rect -96 547 -62 581
rect 62 547 96 581
rect 220 547 254 581
rect 378 547 412 581
rect 536 547 570 581
rect 694 547 728 581
rect 852 547 886 581
rect 1010 547 1044 581
rect 1168 547 1202 581
rect 1326 547 1360 581
rect 1484 547 1518 581
rect -1597 -488 -1563 488
rect -1439 -488 -1405 488
rect -1281 -488 -1247 488
rect -1123 -488 -1089 488
rect -965 -488 -931 488
rect -807 -488 -773 488
rect -649 -488 -615 488
rect -491 -488 -457 488
rect -333 -488 -299 488
rect -175 -488 -141 488
rect -17 -488 17 488
rect 141 -488 175 488
rect 299 -488 333 488
rect 457 -488 491 488
rect 615 -488 649 488
rect 773 -488 807 488
rect 931 -488 965 488
rect 1089 -488 1123 488
rect 1247 -488 1281 488
rect 1405 -488 1439 488
rect 1563 -488 1597 488
rect -1518 -581 -1484 -547
rect -1360 -581 -1326 -547
rect -1202 -581 -1168 -547
rect -1044 -581 -1010 -547
rect -886 -581 -852 -547
rect -728 -581 -694 -547
rect -570 -581 -536 -547
rect -412 -581 -378 -547
rect -254 -581 -220 -547
rect -96 -581 -62 -547
rect 62 -581 96 -547
rect 220 -581 254 -547
rect 378 -581 412 -547
rect 536 -581 570 -547
rect 694 -581 728 -547
rect 852 -581 886 -547
rect 1010 -581 1044 -547
rect 1168 -581 1202 -547
rect 1326 -581 1360 -547
rect 1484 -581 1518 -547
<< metal1 >>
rect -1530 581 -1472 587
rect -1530 547 -1518 581
rect -1484 547 -1472 581
rect -1530 541 -1472 547
rect -1372 581 -1314 587
rect -1372 547 -1360 581
rect -1326 547 -1314 581
rect -1372 541 -1314 547
rect -1214 581 -1156 587
rect -1214 547 -1202 581
rect -1168 547 -1156 581
rect -1214 541 -1156 547
rect -1056 581 -998 587
rect -1056 547 -1044 581
rect -1010 547 -998 581
rect -1056 541 -998 547
rect -898 581 -840 587
rect -898 547 -886 581
rect -852 547 -840 581
rect -898 541 -840 547
rect -740 581 -682 587
rect -740 547 -728 581
rect -694 547 -682 581
rect -740 541 -682 547
rect -582 581 -524 587
rect -582 547 -570 581
rect -536 547 -524 581
rect -582 541 -524 547
rect -424 581 -366 587
rect -424 547 -412 581
rect -378 547 -366 581
rect -424 541 -366 547
rect -266 581 -208 587
rect -266 547 -254 581
rect -220 547 -208 581
rect -266 541 -208 547
rect -108 581 -50 587
rect -108 547 -96 581
rect -62 547 -50 581
rect -108 541 -50 547
rect 50 581 108 587
rect 50 547 62 581
rect 96 547 108 581
rect 50 541 108 547
rect 208 581 266 587
rect 208 547 220 581
rect 254 547 266 581
rect 208 541 266 547
rect 366 581 424 587
rect 366 547 378 581
rect 412 547 424 581
rect 366 541 424 547
rect 524 581 582 587
rect 524 547 536 581
rect 570 547 582 581
rect 524 541 582 547
rect 682 581 740 587
rect 682 547 694 581
rect 728 547 740 581
rect 682 541 740 547
rect 840 581 898 587
rect 840 547 852 581
rect 886 547 898 581
rect 840 541 898 547
rect 998 581 1056 587
rect 998 547 1010 581
rect 1044 547 1056 581
rect 998 541 1056 547
rect 1156 581 1214 587
rect 1156 547 1168 581
rect 1202 547 1214 581
rect 1156 541 1214 547
rect 1314 581 1372 587
rect 1314 547 1326 581
rect 1360 547 1372 581
rect 1314 541 1372 547
rect 1472 581 1530 587
rect 1472 547 1484 581
rect 1518 547 1530 581
rect 1472 541 1530 547
rect -1603 488 -1557 500
rect -1603 -488 -1597 488
rect -1563 -488 -1557 488
rect -1603 -500 -1557 -488
rect -1445 488 -1399 500
rect -1445 -488 -1439 488
rect -1405 -488 -1399 488
rect -1445 -500 -1399 -488
rect -1287 488 -1241 500
rect -1287 -488 -1281 488
rect -1247 -488 -1241 488
rect -1287 -500 -1241 -488
rect -1129 488 -1083 500
rect -1129 -488 -1123 488
rect -1089 -488 -1083 488
rect -1129 -500 -1083 -488
rect -971 488 -925 500
rect -971 -488 -965 488
rect -931 -488 -925 488
rect -971 -500 -925 -488
rect -813 488 -767 500
rect -813 -488 -807 488
rect -773 -488 -767 488
rect -813 -500 -767 -488
rect -655 488 -609 500
rect -655 -488 -649 488
rect -615 -488 -609 488
rect -655 -500 -609 -488
rect -497 488 -451 500
rect -497 -488 -491 488
rect -457 -488 -451 488
rect -497 -500 -451 -488
rect -339 488 -293 500
rect -339 -488 -333 488
rect -299 -488 -293 488
rect -339 -500 -293 -488
rect -181 488 -135 500
rect -181 -488 -175 488
rect -141 -488 -135 488
rect -181 -500 -135 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 135 488 181 500
rect 135 -488 141 488
rect 175 -488 181 488
rect 135 -500 181 -488
rect 293 488 339 500
rect 293 -488 299 488
rect 333 -488 339 488
rect 293 -500 339 -488
rect 451 488 497 500
rect 451 -488 457 488
rect 491 -488 497 488
rect 451 -500 497 -488
rect 609 488 655 500
rect 609 -488 615 488
rect 649 -488 655 488
rect 609 -500 655 -488
rect 767 488 813 500
rect 767 -488 773 488
rect 807 -488 813 488
rect 767 -500 813 -488
rect 925 488 971 500
rect 925 -488 931 488
rect 965 -488 971 488
rect 925 -500 971 -488
rect 1083 488 1129 500
rect 1083 -488 1089 488
rect 1123 -488 1129 488
rect 1083 -500 1129 -488
rect 1241 488 1287 500
rect 1241 -488 1247 488
rect 1281 -488 1287 488
rect 1241 -500 1287 -488
rect 1399 488 1445 500
rect 1399 -488 1405 488
rect 1439 -488 1445 488
rect 1399 -500 1445 -488
rect 1557 488 1603 500
rect 1557 -488 1563 488
rect 1597 -488 1603 488
rect 1557 -500 1603 -488
rect -1530 -547 -1472 -541
rect -1530 -581 -1518 -547
rect -1484 -581 -1472 -547
rect -1530 -587 -1472 -581
rect -1372 -547 -1314 -541
rect -1372 -581 -1360 -547
rect -1326 -581 -1314 -547
rect -1372 -587 -1314 -581
rect -1214 -547 -1156 -541
rect -1214 -581 -1202 -547
rect -1168 -581 -1156 -547
rect -1214 -587 -1156 -581
rect -1056 -547 -998 -541
rect -1056 -581 -1044 -547
rect -1010 -581 -998 -547
rect -1056 -587 -998 -581
rect -898 -547 -840 -541
rect -898 -581 -886 -547
rect -852 -581 -840 -547
rect -898 -587 -840 -581
rect -740 -547 -682 -541
rect -740 -581 -728 -547
rect -694 -581 -682 -547
rect -740 -587 -682 -581
rect -582 -547 -524 -541
rect -582 -581 -570 -547
rect -536 -581 -524 -547
rect -582 -587 -524 -581
rect -424 -547 -366 -541
rect -424 -581 -412 -547
rect -378 -581 -366 -547
rect -424 -587 -366 -581
rect -266 -547 -208 -541
rect -266 -581 -254 -547
rect -220 -581 -208 -547
rect -266 -587 -208 -581
rect -108 -547 -50 -541
rect -108 -581 -96 -547
rect -62 -581 -50 -547
rect -108 -587 -50 -581
rect 50 -547 108 -541
rect 50 -581 62 -547
rect 96 -581 108 -547
rect 50 -587 108 -581
rect 208 -547 266 -541
rect 208 -581 220 -547
rect 254 -581 266 -547
rect 208 -587 266 -581
rect 366 -547 424 -541
rect 366 -581 378 -547
rect 412 -581 424 -547
rect 366 -587 424 -581
rect 524 -547 582 -541
rect 524 -581 536 -547
rect 570 -581 582 -547
rect 524 -587 582 -581
rect 682 -547 740 -541
rect 682 -581 694 -547
rect 728 -581 740 -547
rect 682 -587 740 -581
rect 840 -547 898 -541
rect 840 -581 852 -547
rect 886 -581 898 -547
rect 840 -587 898 -581
rect 998 -547 1056 -541
rect 998 -581 1010 -547
rect 1044 -581 1056 -547
rect 998 -587 1056 -581
rect 1156 -547 1214 -541
rect 1156 -581 1168 -547
rect 1202 -581 1214 -547
rect 1156 -587 1214 -581
rect 1314 -547 1372 -541
rect 1314 -581 1326 -547
rect 1360 -581 1372 -547
rect 1314 -587 1372 -581
rect 1472 -547 1530 -541
rect 1472 -581 1484 -547
rect 1518 -581 1530 -547
rect 1472 -587 1530 -581
<< properties >>
string FIXED_BBOX -1714 -702 1714 702
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 5 l 0.5 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
