magic
tech sky130A
timestamp 1654408082
<< nmoslvt >>
rect -386 -70 -326 70
rect -297 -70 -237 70
rect -208 -70 -148 70
rect -119 -70 -59 70
rect -30 -70 30 70
rect 59 -70 119 70
rect 148 -70 208 70
rect 237 -70 297 70
rect 326 -70 386 70
<< ndiff >>
rect -415 64 -386 70
rect -415 -64 -409 64
rect -392 -64 -386 64
rect -415 -70 -386 -64
rect -326 64 -297 70
rect -326 -64 -320 64
rect -303 -64 -297 64
rect -326 -70 -297 -64
rect -237 64 -208 70
rect -237 -64 -231 64
rect -214 -64 -208 64
rect -237 -70 -208 -64
rect -148 64 -119 70
rect -148 -64 -142 64
rect -125 -64 -119 64
rect -148 -70 -119 -64
rect -59 64 -30 70
rect -59 -64 -53 64
rect -36 -64 -30 64
rect -59 -70 -30 -64
rect 30 64 59 70
rect 30 -64 36 64
rect 53 -64 59 64
rect 30 -70 59 -64
rect 119 64 148 70
rect 119 -64 125 64
rect 142 -64 148 64
rect 119 -70 148 -64
rect 208 64 237 70
rect 208 -64 214 64
rect 231 -64 237 64
rect 208 -70 237 -64
rect 297 64 326 70
rect 297 -64 303 64
rect 320 -64 326 64
rect 297 -70 326 -64
rect 386 64 415 70
rect 386 -64 392 64
rect 409 -64 415 64
rect 386 -70 415 -64
<< ndiffc >>
rect -409 -64 -392 64
rect -320 -64 -303 64
rect -231 -64 -214 64
rect -142 -64 -125 64
rect -53 -64 -36 64
rect 36 -64 53 64
rect 125 -64 142 64
rect 214 -64 231 64
rect 303 -64 320 64
rect 392 -64 409 64
<< poly >>
rect -375 106 -337 114
rect -375 97 -367 106
rect -386 89 -367 97
rect -345 97 -337 106
rect -286 106 -248 114
rect -286 97 -278 106
rect -345 89 -326 97
rect -386 70 -326 89
rect -297 89 -278 97
rect -256 97 -248 106
rect -197 106 -159 114
rect -197 97 -189 106
rect -256 89 -237 97
rect -297 70 -237 89
rect -208 89 -189 97
rect -167 97 -159 106
rect -108 106 -70 114
rect -108 97 -100 106
rect -167 89 -148 97
rect -208 70 -148 89
rect -119 89 -100 97
rect -78 97 -70 106
rect -19 106 19 114
rect -19 97 -11 106
rect -78 89 -59 97
rect -119 70 -59 89
rect -30 89 -11 97
rect 11 97 19 106
rect 70 106 108 114
rect 70 97 78 106
rect 11 89 30 97
rect -30 70 30 89
rect 59 89 78 97
rect 100 97 108 106
rect 159 106 197 114
rect 159 97 167 106
rect 100 89 119 97
rect 59 70 119 89
rect 148 89 167 97
rect 189 97 197 106
rect 248 106 286 114
rect 248 97 256 106
rect 189 89 208 97
rect 148 70 208 89
rect 237 89 256 97
rect 278 97 286 106
rect 337 106 375 114
rect 337 97 345 106
rect 278 89 297 97
rect 237 70 297 89
rect 326 89 345 97
rect 367 97 375 106
rect 367 89 386 97
rect 326 70 386 89
rect -386 -89 -326 -70
rect -386 -97 -367 -89
rect -375 -106 -367 -97
rect -345 -97 -326 -89
rect -297 -89 -237 -70
rect -297 -97 -278 -89
rect -345 -106 -337 -97
rect -375 -114 -337 -106
rect -286 -106 -278 -97
rect -256 -97 -237 -89
rect -208 -89 -148 -70
rect -208 -97 -189 -89
rect -256 -106 -248 -97
rect -286 -114 -248 -106
rect -197 -106 -189 -97
rect -167 -97 -148 -89
rect -119 -89 -59 -70
rect -119 -97 -100 -89
rect -167 -106 -159 -97
rect -197 -114 -159 -106
rect -108 -106 -100 -97
rect -78 -97 -59 -89
rect -30 -89 30 -70
rect -30 -97 -11 -89
rect -78 -106 -70 -97
rect -108 -114 -70 -106
rect -19 -106 -11 -97
rect 11 -97 30 -89
rect 59 -89 119 -70
rect 59 -97 78 -89
rect 11 -106 19 -97
rect -19 -114 19 -106
rect 70 -106 78 -97
rect 100 -97 119 -89
rect 148 -89 208 -70
rect 148 -97 167 -89
rect 100 -106 108 -97
rect 70 -114 108 -106
rect 159 -106 167 -97
rect 189 -97 208 -89
rect 237 -89 297 -70
rect 237 -97 256 -89
rect 189 -106 197 -97
rect 159 -114 197 -106
rect 248 -106 256 -97
rect 278 -97 297 -89
rect 326 -89 386 -70
rect 326 -97 345 -89
rect 278 -106 286 -97
rect 248 -114 286 -106
rect 337 -106 345 -97
rect 367 -97 386 -89
rect 367 -106 375 -97
rect 337 -114 375 -106
<< polycont >>
rect -367 89 -345 106
rect -278 89 -256 106
rect -189 89 -167 106
rect -100 89 -78 106
rect -11 89 11 106
rect 78 89 100 106
rect 167 89 189 106
rect 256 89 278 106
rect 345 89 367 106
rect -367 -106 -345 -89
rect -278 -106 -256 -89
rect -189 -106 -167 -89
rect -100 -106 -78 -89
rect -11 -106 11 -89
rect 78 -106 100 -89
rect 167 -106 189 -89
rect 256 -106 278 -89
rect 345 -106 367 -89
<< locali >>
rect -375 89 -367 106
rect -345 89 -337 106
rect -286 89 -278 106
rect -256 89 -248 106
rect -197 89 -189 106
rect -167 89 -159 106
rect -108 89 -100 106
rect -78 89 -70 106
rect -19 89 -11 106
rect 11 89 19 106
rect 70 89 78 106
rect 100 89 108 106
rect 159 89 167 106
rect 189 89 197 106
rect 248 89 256 106
rect 278 89 286 106
rect 337 89 345 106
rect 367 89 375 106
rect -409 64 -392 72
rect -409 -72 -392 -64
rect -320 64 -303 72
rect -320 -72 -303 -64
rect -231 64 -214 72
rect -231 -72 -214 -64
rect -142 64 -125 72
rect -142 -72 -125 -64
rect -53 64 -36 72
rect -53 -72 -36 -64
rect 36 64 53 72
rect 36 -72 53 -64
rect 125 64 142 72
rect 125 -72 142 -64
rect 214 64 231 72
rect 214 -72 231 -64
rect 303 64 320 72
rect 303 -72 320 -64
rect 392 64 409 72
rect 392 -72 409 -64
rect -375 -106 -367 -89
rect -345 -106 -337 -89
rect -286 -106 -278 -89
rect -256 -106 -248 -89
rect -197 -106 -189 -89
rect -167 -106 -159 -89
rect -108 -106 -100 -89
rect -78 -106 -70 -89
rect -19 -106 -11 -89
rect 11 -106 19 -89
rect 70 -106 78 -89
rect 100 -106 108 -89
rect 159 -106 167 -89
rect 189 -106 197 -89
rect 248 -106 256 -89
rect 278 -106 286 -89
rect 337 -106 345 -89
rect 367 -106 375 -89
<< viali >>
rect -367 89 -345 106
rect -278 89 -256 106
rect -189 89 -167 106
rect -100 89 -78 106
rect -11 89 11 106
rect 78 89 100 106
rect 167 89 189 106
rect 256 89 278 106
rect 345 89 367 106
rect -409 -64 -392 64
rect -320 -64 -303 64
rect -231 -64 -214 64
rect -142 -64 -125 64
rect -53 -64 -36 64
rect 36 -64 53 64
rect 125 -64 142 64
rect 214 -64 231 64
rect 303 -64 320 64
rect 392 -64 409 64
rect -367 -106 -345 -89
rect -278 -106 -256 -89
rect -189 -106 -167 -89
rect -100 -106 -78 -89
rect -11 -106 11 -89
rect 78 -106 100 -89
rect 167 -106 189 -89
rect 256 -106 278 -89
rect 345 -106 367 -89
<< metal1 >>
rect -375 106 -337 114
rect -375 89 -367 106
rect -345 89 -337 106
rect -375 86 -337 89
rect -286 106 -248 114
rect -286 89 -278 106
rect -256 89 -248 106
rect -286 86 -248 89
rect -197 106 -159 114
rect -197 89 -189 106
rect -167 89 -159 106
rect -197 86 -159 89
rect -108 106 -70 114
rect -108 89 -100 106
rect -78 89 -70 106
rect -108 86 -70 89
rect -19 106 19 114
rect -19 89 -11 106
rect 11 89 19 106
rect -19 86 19 89
rect 70 106 108 114
rect 70 89 78 106
rect 100 89 108 106
rect 70 86 108 89
rect 159 106 197 114
rect 159 89 167 106
rect 189 89 197 106
rect 159 86 197 89
rect 248 106 286 114
rect 248 89 256 106
rect 278 89 286 106
rect 248 86 286 89
rect 337 106 375 114
rect 337 89 345 106
rect 367 89 375 106
rect 337 86 375 89
rect -412 64 -389 70
rect -412 -64 -409 64
rect -392 -64 -389 64
rect -412 -70 -389 -64
rect -323 64 -300 70
rect -323 -64 -320 64
rect -303 -64 -300 64
rect -323 -70 -300 -64
rect -234 64 -211 70
rect -234 -64 -231 64
rect -214 -64 -211 64
rect -234 -70 -211 -64
rect -145 64 -122 70
rect -145 -64 -142 64
rect -125 -64 -122 64
rect -145 -70 -122 -64
rect -56 64 -33 70
rect -56 -64 -53 64
rect -36 -64 -33 64
rect -56 -70 -33 -64
rect 33 64 56 70
rect 33 -64 36 64
rect 53 -64 56 64
rect 33 -70 56 -64
rect 122 64 145 70
rect 122 -64 125 64
rect 142 -64 145 64
rect 122 -70 145 -64
rect 211 64 234 70
rect 211 -64 214 64
rect 231 -64 234 64
rect 211 -70 234 -64
rect 300 64 323 70
rect 300 -64 303 64
rect 320 -64 323 64
rect 300 -70 323 -64
rect 389 64 412 70
rect 389 -64 392 64
rect 409 -64 412 64
rect 389 -70 412 -64
rect -375 -89 -337 -86
rect -375 -106 -367 -89
rect -345 -106 -337 -89
rect -375 -114 -337 -106
rect -286 -89 -248 -86
rect -286 -106 -278 -89
rect -256 -106 -248 -89
rect -286 -114 -248 -106
rect -197 -89 -159 -86
rect -197 -106 -189 -89
rect -167 -106 -159 -89
rect -197 -114 -159 -106
rect -108 -89 -70 -86
rect -108 -106 -100 -89
rect -78 -106 -70 -89
rect -108 -114 -70 -106
rect -19 -89 19 -86
rect -19 -106 -11 -89
rect 11 -106 19 -89
rect -19 -114 19 -106
rect 70 -89 108 -86
rect 70 -106 78 -89
rect 100 -106 108 -89
rect 70 -114 108 -106
rect 159 -89 197 -86
rect 159 -106 167 -89
rect 189 -106 197 -89
rect 159 -114 197 -106
rect 248 -89 286 -86
rect 248 -106 256 -89
rect 278 -106 286 -89
rect 248 -114 286 -106
rect 337 -89 375 -86
rect 337 -106 345 -89
rect 367 -106 375 -89
rect 337 -114 375 -106
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1.4 l 0.6 m 1 nf 9 diffcov 100 polycov 50 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
