* NGSPICE file created from transmission_gate_flat.ext - technology: sky130A

.subckt transmission_gate_flat in out en en_b VDD VSS
X0 in en out VSS sky130_fd_pr__nfet_01v8 ad=1.537e+12p pd=1.118e+07u as=1.537e+12p ps=1.118e+07u w=5.3e+06u l=150000u
X1 out en_b in VDD sky130_fd_pr__pfet_01v8 ad=3.973e+12p pd=2.798e+07u as=3.973e+12p ps=2.798e+07u w=1.37e+07u l=150000u
C0 in out 5.84fF
C1 out VDD 2.06fF
C2 en_b in 0.11fF
C3 in en 0.40fF
C4 en_b VDD 0.35fF
C5 VDD en 0.01fF
C6 en_b out 0.06fF
C7 out en 0.13fF
C8 en_b en 0.04fF
C9 in VDD 1.86fF
.ends


x2 clk GND GND VDD VDD net1 sky130_fd_sc_hd__inv_4
V2 VDD GND 1.8
V3 clk GND 1.8
V1 in GND DC 0.9
x1 in n1 clk net1 VDD VSS transmission_gate_flat
x3 __UNCONNECTED_PIN__0 out clk net1 VDD VSS transmission_gate_flat
C1 out GND 1p m=1
XM1 n1 net1 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 

.options savecurrents
.control
op
print v(n1)
write transmission_gate_tb.raw
.endc

.lib /farmshare/home/classes/ee/372/PDKs/open_pdks_1.0.310/sky130/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.inc /farmshare/home/classes/ee/372/PDKs/open_pdks_1.0.310/sky130/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice


.GLOBAL GND
.GLOBAL VDD
.end
