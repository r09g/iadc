magic
tech sky130A
magscale 1 2
timestamp 1652593120
<< nwell >>
rect -954 388 2224 810
<< pwell >>
rect -53 -91 1427 331
rect 668 -208 732 -96
<< nmos >>
rect 157 105 1217 135
<< pmos >>
rect -735 584 2005 614
<< ndiff >>
rect 157 181 1217 193
rect 157 147 169 181
rect 1205 147 1217 181
rect 157 135 1217 147
rect 157 93 1217 105
rect 157 59 169 93
rect 1205 59 1217 93
rect 157 47 1217 59
<< pdiff >>
rect -735 660 2005 672
rect -735 626 -723 660
rect 1993 626 2005 660
rect -735 614 2005 626
rect -735 572 2005 584
rect -735 538 -723 572
rect 1993 538 2005 572
rect -735 526 2005 538
<< ndiffc >>
rect 169 147 1205 181
rect 169 59 1205 93
<< pdiffc >>
rect -723 626 1993 660
rect -723 538 1993 572
<< psubdiff >>
rect -17 261 79 295
rect 1295 261 1391 295
rect -17 199 17 261
rect 1357 199 1391 261
rect -17 -21 17 41
rect 1357 -21 1391 41
rect -17 -55 79 -21
rect 1295 -55 1391 -21
<< nsubdiff >>
rect -918 740 -822 774
rect 2092 740 2188 774
rect -918 678 -884 740
rect 2154 678 2188 740
rect -918 458 -884 520
rect 2154 458 2188 520
rect -918 424 -822 458
rect 2092 424 2188 458
<< psubdiffcont >>
rect 79 261 1295 295
rect -17 41 17 199
rect 1357 41 1391 199
rect 79 -55 1295 -21
<< nsubdiffcont >>
rect -822 740 2092 774
rect -918 520 -884 678
rect 2154 520 2188 678
rect -822 424 2092 458
<< poly >>
rect -832 616 -766 632
rect -832 582 -816 616
rect -782 614 -766 616
rect 2036 616 2102 632
rect 2036 614 2052 616
rect -782 584 -735 614
rect 2005 584 2052 614
rect -782 582 -766 584
rect -832 566 -766 582
rect 2036 582 2052 584
rect 2086 582 2102 616
rect 2036 566 2102 582
rect 69 137 135 153
rect 69 103 85 137
rect 119 135 135 137
rect 1239 137 1305 153
rect 1239 135 1255 137
rect 119 105 157 135
rect 1217 105 1255 135
rect 119 103 135 105
rect 69 87 135 103
rect 1239 103 1255 105
rect 1289 103 1305 137
rect 1239 87 1305 103
<< polycont >>
rect -816 582 -782 616
rect 2052 582 2086 616
rect 85 103 119 137
rect 1255 103 1289 137
<< locali >>
rect -918 740 -822 774
rect 2092 740 2188 774
rect -918 678 -884 740
rect 2154 678 2188 740
rect -816 616 -782 632
rect -739 626 -723 660
rect 1993 626 2009 660
rect -816 566 -782 582
rect 2052 616 2086 632
rect -739 538 -723 572
rect 1993 538 2009 572
rect 2052 566 2086 582
rect -918 458 -884 520
rect 2154 458 2188 520
rect -918 424 -822 458
rect 2092 424 2188 458
rect -17 261 79 295
rect 1295 261 1391 295
rect -17 199 17 261
rect 1357 199 1391 261
rect 85 137 119 153
rect 153 147 169 181
rect 1205 147 1221 181
rect 85 87 119 103
rect 1255 137 1289 153
rect 153 59 169 93
rect 1205 59 1221 93
rect 1255 87 1289 103
rect -17 -21 17 41
rect 1357 -21 1391 41
rect -17 -55 79 -21
rect 1295 -55 1391 -21
<< viali >>
rect 540 740 858 774
rect -723 626 1993 660
rect -816 582 -782 616
rect 2052 582 2086 616
rect -723 538 1993 572
rect 169 147 1205 181
rect 85 103 119 137
rect 1255 103 1289 137
rect 169 59 1205 93
rect 538 -21 856 -20
rect 538 -54 856 -21
<< metal1 >>
rect 662 812 726 922
rect 1922 826 2318 890
rect 528 774 864 812
rect 528 740 540 774
rect 858 740 864 774
rect 528 698 864 740
rect 1922 666 1986 826
rect -735 660 2005 666
rect -1203 616 -776 628
rect -735 626 -723 660
rect 1993 626 2005 660
rect -735 620 2005 626
rect -1203 582 -816 616
rect -782 582 -776 616
rect -1203 570 -776 582
rect 2044 616 2102 634
rect 2044 582 2052 616
rect 2086 582 2102 616
rect -735 572 2005 578
rect -735 538 -723 572
rect 1993 538 2005 572
rect 2044 566 2102 582
rect -735 532 2005 538
rect 196 392 260 532
rect -1202 328 260 392
rect 196 187 260 328
rect 157 181 1217 187
rect 79 148 125 149
rect -1201 137 126 148
rect 157 147 169 181
rect 1205 147 1217 181
rect 157 141 1217 147
rect -1201 103 85 137
rect 119 103 126 137
rect -1201 90 126 103
rect 1248 137 1306 154
rect 1248 103 1255 137
rect 1289 103 1306 137
rect 1152 99 1216 100
rect 157 93 1217 99
rect 157 59 169 93
rect 1205 59 1217 93
rect 1248 86 1306 103
rect 157 53 1217 59
rect 532 -20 862 20
rect 532 -54 538 -20
rect 856 -54 862 -20
rect 532 -96 862 -54
rect 668 -208 732 -96
rect 1152 -98 1216 53
rect 2254 -98 2318 826
rect 1152 -162 2318 -98
<< labels >>
flabel metal1 -1182 120 -1182 120 1 FreeSans 800 0 0 0 en
port 3 n
flabel metal1 -1186 596 -1186 596 1 FreeSans 800 0 0 0 en_b
port 4 n
flabel metal1 -1186 358 -1186 358 1 FreeSans 800 0 0 0 in
port 1 n
flabel metal1 698 -180 698 -180 1 FreeSans 800 0 0 0 VSS
port 6 n
flabel metal1 694 866 694 866 1 FreeSans 800 0 0 0 VDD
port 5 n
flabel metal1 2288 346 2288 346 1 FreeSans 800 0 0 0 out
port 2 n
<< end >>
