magic
tech sky130A
magscale 1 2
timestamp 1654583101
<< error_p >>
rect -512 -184 -446 -176
rect -320 -184 -254 -176
rect -128 -184 -62 -176
rect 64 -184 130 -176
rect 256 -184 322 -176
rect 448 -184 514 -176
rect -512 -218 -496 -184
rect -320 -218 -304 -184
rect -128 -218 -112 -184
rect 64 -218 80 -184
rect 256 -218 272 -184
rect 448 -218 464 -184
rect -512 -226 -446 -218
rect -320 -226 -254 -218
rect -128 -226 -62 -218
rect 64 -226 130 -218
rect 256 -226 322 -218
rect 448 -226 514 -218
<< nwell >>
rect -646 -356 648 294
<< pmos >>
rect -446 -136 -416 136
rect -350 -136 -320 136
rect -254 -136 -224 136
rect -158 -136 -128 136
rect -62 -136 -32 136
rect 34 -136 64 136
rect 130 -136 160 136
rect 226 -136 256 136
rect 322 -136 352 136
rect 418 -136 448 136
<< pdiff >>
rect -508 119 -446 136
rect -508 85 -496 119
rect -462 85 -446 119
rect -508 51 -446 85
rect -508 17 -496 51
rect -462 17 -446 51
rect -508 -17 -446 17
rect -508 -51 -496 -17
rect -462 -51 -446 -17
rect -508 -85 -446 -51
rect -508 -119 -496 -85
rect -462 -119 -446 -85
rect -508 -136 -446 -119
rect -416 119 -350 136
rect -416 85 -400 119
rect -366 85 -350 119
rect -416 51 -350 85
rect -416 17 -400 51
rect -366 17 -350 51
rect -416 -17 -350 17
rect -416 -51 -400 -17
rect -366 -51 -350 -17
rect -416 -85 -350 -51
rect -416 -119 -400 -85
rect -366 -119 -350 -85
rect -416 -136 -350 -119
rect -320 119 -254 136
rect -320 85 -304 119
rect -270 85 -254 119
rect -320 51 -254 85
rect -320 17 -304 51
rect -270 17 -254 51
rect -320 -17 -254 17
rect -320 -51 -304 -17
rect -270 -51 -254 -17
rect -320 -85 -254 -51
rect -320 -119 -304 -85
rect -270 -119 -254 -85
rect -320 -136 -254 -119
rect -224 119 -158 136
rect -224 85 -208 119
rect -174 85 -158 119
rect -224 51 -158 85
rect -224 17 -208 51
rect -174 17 -158 51
rect -224 -17 -158 17
rect -224 -51 -208 -17
rect -174 -51 -158 -17
rect -224 -85 -158 -51
rect -224 -119 -208 -85
rect -174 -119 -158 -85
rect -224 -136 -158 -119
rect -128 119 -62 136
rect -128 85 -112 119
rect -78 85 -62 119
rect -128 51 -62 85
rect -128 17 -112 51
rect -78 17 -62 51
rect -128 -17 -62 17
rect -128 -51 -112 -17
rect -78 -51 -62 -17
rect -128 -85 -62 -51
rect -128 -119 -112 -85
rect -78 -119 -62 -85
rect -128 -136 -62 -119
rect -32 119 34 136
rect -32 85 -16 119
rect 18 85 34 119
rect -32 51 34 85
rect -32 17 -16 51
rect 18 17 34 51
rect -32 -17 34 17
rect -32 -51 -16 -17
rect 18 -51 34 -17
rect -32 -85 34 -51
rect -32 -119 -16 -85
rect 18 -119 34 -85
rect -32 -136 34 -119
rect 64 119 130 136
rect 64 85 80 119
rect 114 85 130 119
rect 64 51 130 85
rect 64 17 80 51
rect 114 17 130 51
rect 64 -17 130 17
rect 64 -51 80 -17
rect 114 -51 130 -17
rect 64 -85 130 -51
rect 64 -119 80 -85
rect 114 -119 130 -85
rect 64 -136 130 -119
rect 160 119 226 136
rect 160 85 176 119
rect 210 85 226 119
rect 160 51 226 85
rect 160 17 176 51
rect 210 17 226 51
rect 160 -17 226 17
rect 160 -51 176 -17
rect 210 -51 226 -17
rect 160 -85 226 -51
rect 160 -119 176 -85
rect 210 -119 226 -85
rect 160 -136 226 -119
rect 256 119 322 136
rect 256 85 272 119
rect 306 85 322 119
rect 256 51 322 85
rect 256 17 272 51
rect 306 17 322 51
rect 256 -17 322 17
rect 256 -51 272 -17
rect 306 -51 322 -17
rect 256 -85 322 -51
rect 256 -119 272 -85
rect 306 -119 322 -85
rect 256 -136 322 -119
rect 352 119 418 136
rect 352 85 368 119
rect 402 85 418 119
rect 352 51 418 85
rect 352 17 368 51
rect 402 17 418 51
rect 352 -17 418 17
rect 352 -51 368 -17
rect 402 -51 418 -17
rect 352 -85 418 -51
rect 352 -119 368 -85
rect 402 -119 418 -85
rect 352 -136 418 -119
rect 448 119 510 136
rect 448 85 464 119
rect 498 85 510 119
rect 448 51 510 85
rect 448 17 464 51
rect 498 17 510 51
rect 448 -17 510 17
rect 448 -51 464 -17
rect 498 -51 510 -17
rect 448 -85 510 -51
rect 448 -119 464 -85
rect 498 -119 510 -85
rect 448 -136 510 -119
<< pdiffc >>
rect -496 85 -462 119
rect -496 17 -462 51
rect -496 -51 -462 -17
rect -496 -119 -462 -85
rect -400 85 -366 119
rect -400 17 -366 51
rect -400 -51 -366 -17
rect -400 -119 -366 -85
rect -304 85 -270 119
rect -304 17 -270 51
rect -304 -51 -270 -17
rect -304 -119 -270 -85
rect -208 85 -174 119
rect -208 17 -174 51
rect -208 -51 -174 -17
rect -208 -119 -174 -85
rect -112 85 -78 119
rect -112 17 -78 51
rect -112 -51 -78 -17
rect -112 -119 -78 -85
rect -16 85 18 119
rect -16 17 18 51
rect -16 -51 18 -17
rect -16 -119 18 -85
rect 80 85 114 119
rect 80 17 114 51
rect 80 -51 114 -17
rect 80 -119 114 -85
rect 176 85 210 119
rect 176 17 210 51
rect 176 -51 210 -17
rect 176 -119 210 -85
rect 272 85 306 119
rect 272 17 306 51
rect 272 -51 306 -17
rect 272 -119 306 -85
rect 368 85 402 119
rect 368 17 402 51
rect 368 -51 402 -17
rect 368 -119 402 -85
rect 464 85 498 119
rect 464 17 498 51
rect 464 -51 498 -17
rect 464 -119 498 -85
<< nsubdiff >>
rect -610 224 -492 258
rect -458 224 -424 258
rect -390 224 -356 258
rect -322 224 -288 258
rect -254 224 -220 258
rect -186 224 -152 258
rect -118 224 -84 258
rect -50 224 -16 258
rect 18 224 52 258
rect 86 224 120 258
rect 154 224 188 258
rect 222 224 256 258
rect 290 224 324 258
rect 358 224 392 258
rect 426 224 460 258
rect 494 224 612 258
rect -610 156 -576 224
rect 578 156 612 224
rect -610 88 -576 122
rect -610 20 -576 54
rect -610 -48 -576 -14
rect -610 -116 -576 -82
rect 578 88 612 122
rect 578 20 612 54
rect 578 -48 612 -14
rect 578 -116 612 -82
rect -610 -184 -576 -150
rect -610 -286 -576 -218
rect 578 -184 612 -150
rect 578 -286 612 -218
rect -610 -320 -492 -286
rect -458 -320 -424 -286
rect -390 -320 -356 -286
rect -322 -320 -288 -286
rect -254 -320 -220 -286
rect -186 -320 -152 -286
rect -118 -320 -84 -286
rect -50 -320 -16 -286
rect 18 -320 52 -286
rect 86 -320 120 -286
rect 154 -320 188 -286
rect 222 -320 256 -286
rect 290 -320 324 -286
rect 358 -320 392 -286
rect 426 -320 460 -286
rect 494 -320 612 -286
<< nsubdiffcont >>
rect -492 224 -458 258
rect -424 224 -390 258
rect -356 224 -322 258
rect -288 224 -254 258
rect -220 224 -186 258
rect -152 224 -118 258
rect -84 224 -50 258
rect -16 224 18 258
rect 52 224 86 258
rect 120 224 154 258
rect 188 224 222 258
rect 256 224 290 258
rect 324 224 358 258
rect 392 224 426 258
rect 460 224 494 258
rect -610 122 -576 156
rect -610 54 -576 88
rect -610 -14 -576 20
rect -610 -82 -576 -48
rect -610 -150 -576 -116
rect 578 122 612 156
rect 578 54 612 88
rect 578 -14 612 20
rect 578 -82 612 -48
rect 578 -150 612 -116
rect -610 -218 -576 -184
rect 578 -218 612 -184
rect -492 -320 -458 -286
rect -424 -320 -390 -286
rect -356 -320 -322 -286
rect -288 -320 -254 -286
rect -220 -320 -186 -286
rect -152 -320 -118 -286
rect -84 -320 -50 -286
rect -16 -320 18 -286
rect 52 -320 86 -286
rect 120 -320 154 -286
rect 188 -320 222 -286
rect 256 -320 290 -286
rect 324 -320 358 -286
rect 392 -320 426 -286
rect 460 -320 494 -286
<< poly >>
rect -446 136 -416 162
rect -350 136 -320 162
rect -254 136 -224 162
rect -158 136 -128 162
rect -62 136 -32 162
rect 34 136 64 162
rect 130 136 160 162
rect 226 136 256 162
rect 322 136 352 162
rect 418 136 448 162
rect -446 -168 -416 -136
rect -350 -168 -320 -136
rect -254 -168 -224 -136
rect -158 -168 -128 -136
rect -62 -168 -32 -136
rect 34 -168 64 -136
rect 130 -168 160 -136
rect 226 -168 256 -136
rect 322 -168 352 -136
rect 418 -168 448 -136
rect -512 -184 514 -168
rect -512 -218 -496 -184
rect -462 -218 -304 -184
rect -270 -218 -112 -184
rect -78 -218 80 -184
rect 114 -218 272 -184
rect 306 -218 464 -184
rect 498 -218 514 -184
rect -512 -234 514 -218
<< polycont >>
rect -496 -218 -462 -184
rect -304 -218 -270 -184
rect -112 -218 -78 -184
rect 80 -218 114 -184
rect 272 -218 306 -184
rect 464 -218 498 -184
<< locali >>
rect -610 224 -492 258
rect -458 224 -424 258
rect -390 224 -356 258
rect -322 224 -288 258
rect -254 224 -220 258
rect -186 224 -152 258
rect -118 224 -84 258
rect -50 224 -16 258
rect 18 224 52 258
rect 86 224 120 258
rect 154 224 188 258
rect 222 224 256 258
rect 290 224 324 258
rect 358 224 392 258
rect 426 224 460 258
rect 494 224 612 258
rect -610 156 -576 224
rect 578 156 612 224
rect -610 88 -576 122
rect -610 20 -576 54
rect -610 -48 -576 -14
rect -610 -116 -576 -82
rect -496 119 -462 140
rect -496 51 -462 55
rect -496 -55 -462 -51
rect -496 -140 -462 -119
rect -400 119 -366 140
rect -400 51 -366 55
rect -400 -55 -366 -51
rect -400 -140 -366 -119
rect -304 119 -270 140
rect -304 51 -270 55
rect -304 -55 -270 -51
rect -304 -140 -270 -119
rect -208 119 -174 140
rect -208 51 -174 55
rect -208 -55 -174 -51
rect -208 -140 -174 -119
rect -112 119 -78 140
rect -112 51 -78 55
rect -112 -55 -78 -51
rect -112 -140 -78 -119
rect -16 119 18 140
rect -16 51 18 55
rect -16 -55 18 -51
rect -16 -140 18 -119
rect 80 119 114 140
rect 80 51 114 55
rect 80 -55 114 -51
rect 80 -140 114 -119
rect 176 119 210 140
rect 176 51 210 55
rect 176 -55 210 -51
rect 176 -140 210 -119
rect 272 119 306 140
rect 272 51 306 55
rect 272 -55 306 -51
rect 272 -140 306 -119
rect 368 119 402 140
rect 368 51 402 55
rect 368 -55 402 -51
rect 368 -140 402 -119
rect 464 119 498 140
rect 464 51 498 55
rect 464 -55 498 -51
rect 464 -140 498 -119
rect 578 88 612 122
rect 578 20 612 54
rect 578 -48 612 -14
rect 578 -116 612 -82
rect -610 -184 -576 -150
rect 578 -184 612 -150
rect -512 -218 -496 -184
rect -462 -218 -446 -184
rect -320 -218 -304 -184
rect -270 -218 -254 -184
rect -128 -218 -112 -184
rect -78 -218 -62 -184
rect 64 -218 80 -184
rect 114 -218 130 -184
rect 256 -218 272 -184
rect 306 -218 322 -184
rect 448 -218 464 -184
rect 498 -218 514 -184
rect -610 -286 -576 -218
rect 578 -286 612 -218
rect -610 -320 -492 -286
rect -458 -320 -424 -286
rect -390 -320 -356 -286
rect -322 -320 -288 -286
rect -254 -320 -220 -286
rect -186 -320 -152 -286
rect -118 -320 -84 -286
rect -50 -320 -16 -286
rect 18 -320 52 -286
rect 86 -320 120 -286
rect 154 -320 188 -286
rect 222 -320 256 -286
rect 290 -320 324 -286
rect 358 -320 392 -286
rect 426 -320 460 -286
rect 494 -320 612 -286
<< viali >>
rect -496 85 -462 89
rect -496 55 -462 85
rect -496 -17 -462 17
rect -496 -85 -462 -55
rect -496 -89 -462 -85
rect -400 85 -366 89
rect -400 55 -366 85
rect -400 -17 -366 17
rect -400 -85 -366 -55
rect -400 -89 -366 -85
rect -304 85 -270 89
rect -304 55 -270 85
rect -304 -17 -270 17
rect -304 -85 -270 -55
rect -304 -89 -270 -85
rect -208 85 -174 89
rect -208 55 -174 85
rect -208 -17 -174 17
rect -208 -85 -174 -55
rect -208 -89 -174 -85
rect -112 85 -78 89
rect -112 55 -78 85
rect -112 -17 -78 17
rect -112 -85 -78 -55
rect -112 -89 -78 -85
rect -16 85 18 89
rect -16 55 18 85
rect -16 -17 18 17
rect -16 -85 18 -55
rect -16 -89 18 -85
rect 80 85 114 89
rect 80 55 114 85
rect 80 -17 114 17
rect 80 -85 114 -55
rect 80 -89 114 -85
rect 176 85 210 89
rect 176 55 210 85
rect 176 -17 210 17
rect 176 -85 210 -55
rect 176 -89 210 -85
rect 272 85 306 89
rect 272 55 306 85
rect 272 -17 306 17
rect 272 -85 306 -55
rect 272 -89 306 -85
rect 368 85 402 89
rect 368 55 402 85
rect 368 -17 402 17
rect 368 -85 402 -55
rect 368 -89 402 -85
rect 464 85 498 89
rect 464 55 498 85
rect 464 -17 498 17
rect 464 -85 498 -55
rect 464 -89 498 -85
rect -496 -218 -462 -184
rect -304 -218 -270 -184
rect -112 -218 -78 -184
rect 80 -218 114 -184
rect 272 -218 306 -184
rect 464 -218 498 -184
<< metal1 >>
rect -502 89 -456 136
rect -502 55 -496 89
rect -462 55 -456 89
rect -502 17 -456 55
rect -502 -17 -496 17
rect -462 -17 -456 17
rect -502 -55 -456 -17
rect -502 -89 -496 -55
rect -462 -89 -456 -55
rect -502 -136 -456 -89
rect -406 89 -360 136
rect -406 55 -400 89
rect -366 55 -360 89
rect -406 17 -360 55
rect -406 -17 -400 17
rect -366 -17 -360 17
rect -406 -55 -360 -17
rect -406 -89 -400 -55
rect -366 -89 -360 -55
rect -406 -136 -360 -89
rect -310 89 -264 136
rect -310 55 -304 89
rect -270 55 -264 89
rect -310 17 -264 55
rect -310 -17 -304 17
rect -270 -17 -264 17
rect -310 -55 -264 -17
rect -310 -89 -304 -55
rect -270 -89 -264 -55
rect -310 -136 -264 -89
rect -214 89 -168 136
rect -214 55 -208 89
rect -174 55 -168 89
rect -214 17 -168 55
rect -214 -17 -208 17
rect -174 -17 -168 17
rect -214 -55 -168 -17
rect -214 -89 -208 -55
rect -174 -89 -168 -55
rect -214 -136 -168 -89
rect -118 89 -72 136
rect -118 55 -112 89
rect -78 55 -72 89
rect -118 17 -72 55
rect -118 -17 -112 17
rect -78 -17 -72 17
rect -118 -55 -72 -17
rect -118 -89 -112 -55
rect -78 -89 -72 -55
rect -118 -136 -72 -89
rect -22 89 24 136
rect -22 55 -16 89
rect 18 55 24 89
rect -22 17 24 55
rect -22 -17 -16 17
rect 18 -17 24 17
rect -22 -55 24 -17
rect -22 -89 -16 -55
rect 18 -89 24 -55
rect -22 -136 24 -89
rect 74 89 120 136
rect 74 55 80 89
rect 114 55 120 89
rect 74 17 120 55
rect 74 -17 80 17
rect 114 -17 120 17
rect 74 -55 120 -17
rect 74 -89 80 -55
rect 114 -89 120 -55
rect 74 -136 120 -89
rect 170 89 216 136
rect 170 55 176 89
rect 210 55 216 89
rect 170 17 216 55
rect 170 -17 176 17
rect 210 -17 216 17
rect 170 -55 216 -17
rect 170 -89 176 -55
rect 210 -89 216 -55
rect 170 -136 216 -89
rect 266 89 312 136
rect 266 55 272 89
rect 306 55 312 89
rect 266 17 312 55
rect 266 -17 272 17
rect 306 -17 312 17
rect 266 -55 312 -17
rect 266 -89 272 -55
rect 306 -89 312 -55
rect 266 -136 312 -89
rect 362 89 408 136
rect 362 55 368 89
rect 402 55 408 89
rect 362 17 408 55
rect 362 -17 368 17
rect 402 -17 408 17
rect 362 -55 408 -17
rect 362 -89 368 -55
rect 402 -89 408 -55
rect 362 -136 408 -89
rect 458 89 504 136
rect 458 55 464 89
rect 498 55 504 89
rect 458 17 504 55
rect 458 -17 464 17
rect 498 -17 504 17
rect 458 -55 504 -17
rect 458 -89 464 -55
rect 498 -89 504 -55
rect 458 -136 504 -89
rect -512 -184 -446 -176
rect -512 -218 -496 -184
rect -462 -218 -446 -184
rect -512 -226 -446 -218
rect -320 -184 -254 -176
rect -320 -218 -304 -184
rect -270 -218 -254 -184
rect -320 -226 -254 -218
rect -128 -184 -62 -176
rect -128 -218 -112 -184
rect -78 -218 -62 -184
rect -128 -226 -62 -218
rect 64 -184 130 -176
rect 64 -218 80 -184
rect 114 -218 130 -184
rect 64 -226 130 -218
rect 256 -184 322 -176
rect 256 -218 272 -184
rect 306 -218 322 -184
rect 256 -226 322 -218
rect 448 -184 514 -176
rect 448 -218 464 -184
rect 498 -218 514 -184
rect 448 -226 514 -218
<< properties >>
string FIXED_BBOX -594 -302 594 302
<< end >>
