* NGSPICE file created from esd_cell.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_g5v0d10v5_BRTJC6 a_n345_n500# a_1135_n588# a_n603_n588#
+ a_n1393_n588# a_n1609_n500# a_661_n588# a_n1135_n500# a_n977_n500# a_1293_n588#
+ a_n761_n588# a_n503_n500# a_n1551_n588# a_129_n500# a_n1293_n500# a_287_n500# a_n661_n500#
+ a_1451_n588# a_n1451_n500# a_919_n500# a_445_n500# a_1077_n500# a_29_n588# a_n129_n588#
+ a_603_n500# a_187_n588# a_1235_n500# a_n287_n588# a_761_n500# a_819_n588# a_345_n588#
+ a_n1077_n588# a_n29_n500# a_1393_n500# a_n919_n588# a_n1743_n722# a_n187_n500# a_977_n588#
+ a_n445_n588# a_503_n588# a_n1235_n588# a_1551_n500# a_n819_n500#
X0 a_n819_n500# a_n919_n588# a_n977_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X1 a_n661_n500# a_n761_n588# a_n819_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X2 a_919_n500# a_819_n588# a_761_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X3 a_n187_n500# a_n287_n588# a_n345_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X4 a_761_n500# a_661_n588# a_603_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X5 a_287_n500# a_187_n588# a_129_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X6 a_n1293_n500# a_n1393_n588# a_n1451_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X7 a_1393_n500# a_1293_n588# a_1235_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X8 a_n345_n500# a_n445_n588# a_n503_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X9 a_129_n500# a_29_n588# a_n29_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X10 a_445_n500# a_345_n588# a_287_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X11 a_n1451_n500# a_n1551_n588# a_n1609_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X12 a_1551_n500# a_1451_n588# a_1393_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X13 a_n977_n500# a_n1077_n588# a_n1135_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X14 a_n503_n500# a_n603_n588# a_n661_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X15 a_1077_n500# a_977_n588# a_919_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X16 a_n29_n500# a_n129_n588# a_n187_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X17 a_603_n500# a_503_n588# a_445_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X18 a_n1135_n500# a_n1235_n588# a_n1293_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X19 a_1235_n500# a_1135_n588# a_1077_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
C0 a_1393_n500# a_1551_n500# 0.56fF
C1 a_1235_n500# a_1551_n500# 0.24fF
C2 a_1551_n500# a_1077_n500# 0.15fF
C3 a_1393_n500# a_1235_n500# 0.56fF
C4 a_1393_n500# a_1077_n500# 0.24fF
C5 a_1235_n500# a_1077_n500# 0.56fF
C6 a_919_n500# a_1551_n500# 0.11fF
C7 a_1551_n500# a_603_n500# 0.07fF
C8 a_919_n500# a_1393_n500# 0.15fF
C9 a_919_n500# a_1235_n500# 0.24fF
C10 a_761_n500# a_1551_n500# 0.09fF
C11 a_919_n500# a_1077_n500# 0.56fF
C12 a_1393_n500# a_603_n500# 0.09fF
C13 a_1551_n500# a_445_n500# 0.06fF
C14 a_1235_n500# a_603_n500# 0.11fF
C15 a_1077_n500# a_603_n500# 0.15fF
C16 a_1393_n500# a_761_n500# 0.11fF
C17 a_1235_n500# a_761_n500# 0.15fF
C18 a_761_n500# a_1077_n500# 0.24fF
C19 a_1393_n500# a_445_n500# 0.07fF
C20 a_n29_n500# a_1551_n500# 0.04fF
C21 a_1551_n500# a_287_n500# 0.05fF
C22 a_1235_n500# a_445_n500# 0.09fF
C23 a_445_n500# a_1077_n500# 0.11fF
C24 a_1551_n500# a_129_n500# 0.05fF
C25 a_n29_n500# a_1393_n500# 0.05fF
C26 a_1393_n500# a_287_n500# 0.06fF
C27 a_n29_n500# a_1235_n500# 0.05fF
C28 a_1235_n500# a_287_n500# 0.07fF
C29 a_1393_n500# a_129_n500# 0.05fF
C30 a_n29_n500# a_1077_n500# 0.06fF
C31 a_1077_n500# a_287_n500# 0.09fF
C32 a_919_n500# a_603_n500# 0.24fF
C33 a_1235_n500# a_129_n500# 0.06fF
C34 a_129_n500# a_1077_n500# 0.07fF
C35 a_919_n500# a_761_n500# 0.56fF
C36 a_1393_n500# a_n187_n500# 0.04fF
C37 a_1235_n500# a_n345_n500# 0.04fF
C38 a_919_n500# a_445_n500# 0.15fF
C39 a_n345_n500# a_1077_n500# 0.05fF
C40 a_1235_n500# a_n187_n500# 0.05fF
C41 a_n187_n500# a_1077_n500# 0.05fF
C42 a_761_n500# a_603_n500# 0.56fF
C43 a_445_n500# a_603_n500# 0.56fF
C44 a_1077_n500# a_n503_n500# 0.04fF
C45 a_919_n500# a_n29_n500# 0.07fF
C46 a_919_n500# a_287_n500# 0.11fF
C47 a_761_n500# a_445_n500# 0.24fF
C48 a_919_n500# a_129_n500# 0.09fF
C49 a_287_n500# a_603_n500# 0.24fF
C50 a_n29_n500# a_603_n500# 0.11fF
C51 a_919_n500# a_n345_n500# 0.05fF
C52 a_919_n500# a_n187_n500# 0.06fF
C53 a_129_n500# a_603_n500# 0.15fF
C54 a_n29_n500# a_761_n500# 0.09fF
C55 a_761_n500# a_287_n500# 0.15fF
C56 a_761_n500# a_129_n500# 0.11fF
C57 a_445_n500# a_287_n500# 0.56fF
C58 a_n29_n500# a_445_n500# 0.15fF
C59 a_919_n500# a_n503_n500# 0.05fF
C60 a_n345_n500# a_603_n500# 0.07fF
C61 a_n187_n500# a_603_n500# 0.09fF
C62 a_445_n500# a_129_n500# 0.24fF
C63 a_761_n500# a_n345_n500# 0.06fF
C64 a_761_n500# a_n187_n500# 0.07fF
C65 a_n661_n500# a_919_n500# 0.04fF
C66 a_n29_n500# a_287_n500# 0.24fF
C67 a_603_n500# a_n503_n500# 0.06fF
C68 a_n345_n500# a_445_n500# 0.09fF
C69 a_445_n500# a_n187_n500# 0.11fF
C70 a_129_n500# a_287_n500# 0.56fF
C71 a_761_n500# a_n503_n500# 0.05fF
C72 a_n29_n500# a_129_n500# 0.56fF
C73 a_n661_n500# a_603_n500# 0.05fF
C74 a_445_n500# a_n503_n500# 0.07fF
C75 a_n345_n500# a_287_n500# 0.11fF
C76 a_n661_n500# a_761_n500# 0.05fF
C77 a_n29_n500# a_n345_n500# 0.24fF
C78 a_n29_n500# a_n187_n500# 0.56fF
C79 a_n187_n500# a_287_n500# 0.15fF
C80 a_n819_n500# a_603_n500# 0.05fF
C81 a_n345_n500# a_129_n500# 0.15fF
C82 a_761_n500# a_n819_n500# 0.04fF
C83 a_n187_n500# a_129_n500# 0.24fF
C84 a_n661_n500# a_445_n500# 0.06fF
C85 a_287_n500# a_n503_n500# 0.09fF
C86 a_n29_n500# a_n503_n500# 0.15fF
C87 a_445_n500# a_n819_n500# 0.05fF
C88 a_n345_n500# a_n187_n500# 0.56fF
C89 a_129_n500# a_n503_n500# 0.11fF
C90 a_n661_n500# a_287_n500# 0.07fF
C91 a_n977_n500# a_603_n500# 0.04fF
C92 a_n661_n500# a_n29_n500# 0.11fF
C93 a_n345_n500# a_n503_n500# 0.56fF
C94 a_287_n500# a_n819_n500# 0.06fF
C95 a_n661_n500# a_129_n500# 0.09fF
C96 a_n29_n500# a_n819_n500# 0.09fF
C97 a_n187_n500# a_n503_n500# 0.24fF
C98 a_445_n500# a_n1135_n500# 0.04fF
C99 a_129_n500# a_n819_n500# 0.07fF
C100 a_n977_n500# a_445_n500# 0.05fF
C101 a_n661_n500# a_n345_n500# 0.24fF
C102 a_n661_n500# a_n187_n500# 0.15fF
C103 a_n345_n500# a_n819_n500# 0.15fF
C104 a_n187_n500# a_n819_n500# 0.11fF
C105 a_287_n500# a_n1135_n500# 0.05fF
C106 a_n29_n500# a_n1135_n500# 0.06fF
C107 a_n977_n500# a_287_n500# 0.05fF
C108 a_n29_n500# a_n977_n500# 0.07fF
C109 a_n661_n500# a_n503_n500# 0.56fF
C110 a_129_n500# a_n1135_n500# 0.05fF
C111 a_n977_n500# a_129_n500# 0.06fF
C112 a_n819_n500# a_n503_n500# 0.24fF
C113 a_n345_n500# a_n1135_n500# 0.09fF
C114 a_n345_n500# a_n977_n500# 0.11fF
C115 a_n187_n500# a_n1135_n500# 0.07fF
C116 a_n977_n500# a_n187_n500# 0.09fF
C117 a_n661_n500# a_n819_n500# 0.56fF
C118 a_n1135_n500# a_n503_n500# 0.11fF
C119 a_n977_n500# a_n503_n500# 0.15fF
C120 a_n661_n500# a_n1135_n500# 0.15fF
C121 a_n661_n500# a_n977_n500# 0.24fF
C122 a_n1293_n500# a_287_n500# 0.04fF
C123 a_n29_n500# a_n1293_n500# 0.05fF
C124 a_n1451_n500# a_n29_n500# 0.05fF
C125 a_n819_n500# a_n1135_n500# 0.24fF
C126 a_n29_n500# a_n1609_n500# 0.04fF
C127 a_n977_n500# a_n819_n500# 0.56fF
C128 a_n1293_n500# a_129_n500# 0.05fF
C129 a_n1451_n500# a_129_n500# 0.04fF
C130 a_n345_n500# a_n1293_n500# 0.07fF
C131 a_n1451_n500# a_n345_n500# 0.06fF
C132 a_n1293_n500# a_n187_n500# 0.06fF
C133 a_n345_n500# a_n1609_n500# 0.05fF
C134 a_n1451_n500# a_n187_n500# 0.05fF
C135 a_n187_n500# a_n1609_n500# 0.05fF
C136 a_n977_n500# a_n1135_n500# 0.56fF
C137 a_n1293_n500# a_n503_n500# 0.09fF
C138 a_n1451_n500# a_n503_n500# 0.07fF
C139 a_n1609_n500# a_n503_n500# 0.06fF
C140 a_n661_n500# a_n1293_n500# 0.11fF
C141 a_n1451_n500# a_n661_n500# 0.09fF
C142 a_n661_n500# a_n1609_n500# 0.07fF
C143 a_n1293_n500# a_n819_n500# 0.15fF
C144 a_n1451_n500# a_n819_n500# 0.11fF
C145 a_n1609_n500# a_n819_n500# 0.09fF
C146 a_n1293_n500# a_n1135_n500# 0.56fF
C147 a_n1451_n500# a_n1135_n500# 0.24fF
C148 a_n1293_n500# a_n977_n500# 0.24fF
C149 a_n1451_n500# a_n977_n500# 0.15fF
C150 a_n1609_n500# a_n1135_n500# 0.15fF
C151 a_n977_n500# a_n1609_n500# 0.11fF
C152 a_n1451_n500# a_n1293_n500# 0.56fF
C153 a_n1293_n500# a_n1609_n500# 0.24fF
C154 a_n1451_n500# a_n1609_n500# 0.56fF
C155 a_1135_n588# a_1293_n588# 0.12fF
C156 a_1293_n588# a_1451_n588# 0.12fF
C157 a_1135_n588# a_1451_n588# 0.04fF
C158 a_1293_n588# a_977_n588# 0.04fF
C159 a_1135_n588# a_977_n588# 0.12fF
C160 a_977_n588# a_1451_n588# 0.02fF
C161 a_1293_n588# a_819_n588# 0.02fF
C162 a_1135_n588# a_819_n588# 0.04fF
C163 a_1293_n588# a_661_n588# 0.02fF
C164 a_1451_n588# a_819_n588# 0.02fF
C165 a_1135_n588# a_661_n588# 0.02fF
C166 a_661_n588# a_1451_n588# 0.01fF
C167 a_977_n588# a_819_n588# 0.12fF
C168 a_661_n588# a_977_n588# 0.04fF
C169 a_1293_n588# a_503_n588# 0.01fF
C170 a_661_n588# a_819_n588# 0.12fF
C171 a_1135_n588# a_503_n588# 0.02fF
C172 a_503_n588# a_1451_n588# 0.01fF
C173 a_1293_n588# a_345_n588# 0.01fF
C174 a_503_n588# a_977_n588# 0.02fF
C175 a_1135_n588# a_345_n588# 0.01fF
C176 a_345_n588# a_1451_n588# 0.01fF
C177 a_1293_n588# a_187_n588# 0.01fF
C178 a_345_n588# a_977_n588# 0.02fF
C179 a_29_n588# a_1293_n588# 0.01fF
C180 a_503_n588# a_819_n588# 0.04fF
C181 a_1293_n588# a_n287_n588# 0.01fF
C182 a_1135_n588# a_187_n588# 0.01fF
C183 a_29_n588# a_1135_n588# 0.01fF
C184 a_n129_n588# a_1293_n588# 0.01fF
C185 a_661_n588# a_503_n588# 0.12fF
C186 a_1135_n588# a_n287_n588# 0.01fF
C187 a_1451_n588# a_187_n588# 0.01fF
C188 a_29_n588# a_1451_n588# 0.01fF
C189 a_n445_n588# a_1135_n588# 0.01fF
C190 a_345_n588# a_819_n588# 0.02fF
C191 a_n129_n588# a_1135_n588# 0.01fF
C192 a_977_n588# a_187_n588# 0.01fF
C193 a_29_n588# a_977_n588# 0.01fF
C194 a_661_n588# a_345_n588# 0.04fF
C195 a_977_n588# a_n287_n588# 0.01fF
C196 a_n129_n588# a_1451_n588# 0.01fF
C197 a_n445_n588# a_977_n588# 0.01fF
C198 a_n129_n588# a_977_n588# 0.01fF
C199 a_187_n588# a_819_n588# 0.02fF
C200 a_29_n588# a_819_n588# 0.01fF
C201 a_n287_n588# a_819_n588# 0.01fF
C202 a_n603_n588# a_977_n588# 0.01fF
C203 a_661_n588# a_187_n588# 0.02fF
C204 a_n445_n588# a_819_n588# 0.01fF
C205 a_29_n588# a_661_n588# 0.02fF
C206 a_n129_n588# a_819_n588# 0.01fF
C207 a_661_n588# a_n287_n588# 0.01fF
C208 a_n445_n588# a_661_n588# 0.01fF
C209 a_n129_n588# a_661_n588# 0.01fF
C210 a_503_n588# a_345_n588# 0.12fF
C211 a_n603_n588# a_819_n588# 0.01fF
C212 a_n603_n588# a_661_n588# 0.01fF
C213 a_n761_n588# a_819_n588# 0.01fF
C214 a_503_n588# a_187_n588# 0.04fF
C215 a_29_n588# a_503_n588# 0.02fF
C216 a_503_n588# a_n287_n588# 0.01fF
C217 a_n761_n588# a_661_n588# 0.01fF
C218 a_n445_n588# a_503_n588# 0.01fF
C219 a_n919_n588# a_661_n588# 0.01fF
C220 a_n129_n588# a_503_n588# 0.02fF
C221 a_345_n588# a_187_n588# 0.12fF
C222 a_29_n588# a_345_n588# 0.04fF
C223 a_345_n588# a_n287_n588# 0.02fF
C224 a_n445_n588# a_345_n588# 0.01fF
C225 a_n603_n588# a_503_n588# 0.01fF
C226 a_n129_n588# a_345_n588# 0.02fF
C227 a_29_n588# a_187_n588# 0.12fF
C228 a_187_n588# a_n287_n588# 0.02fF
C229 a_503_n588# a_n1077_n588# 0.01fF
C230 a_n603_n588# a_345_n588# 0.01fF
C231 a_29_n588# a_n287_n588# 0.04fF
C232 a_n761_n588# a_503_n588# 0.01fF
C233 a_n445_n588# a_187_n588# 0.02fF
C234 a_n919_n588# a_503_n588# 0.01fF
C235 a_29_n588# a_n445_n588# 0.02fF
C236 a_n129_n588# a_187_n588# 0.04fF
C237 a_n445_n588# a_n287_n588# 0.12fF
C238 a_29_n588# a_n129_n588# 0.12fF
C239 a_n129_n588# a_n287_n588# 0.12fF
C240 a_345_n588# a_n1077_n588# 0.01fF
C241 a_n761_n588# a_345_n588# 0.01fF
C242 a_n445_n588# a_n129_n588# 0.04fF
C243 a_n603_n588# a_187_n588# 0.01fF
C244 a_29_n588# a_n603_n588# 0.02fF
C245 a_345_n588# a_n1235_n588# 0.01fF
C246 a_n919_n588# a_345_n588# 0.01fF
C247 a_n603_n588# a_n287_n588# 0.04fF
C248 a_n445_n588# a_n603_n588# 0.12fF
C249 a_n129_n588# a_n603_n588# 0.02fF
C250 a_n1077_n588# a_187_n588# 0.01fF
C251 a_n761_n588# a_187_n588# 0.01fF
C252 a_29_n588# a_n1077_n588# 0.01fF
C253 a_29_n588# a_n761_n588# 0.01fF
C254 a_n1077_n588# a_n287_n588# 0.01fF
C255 a_n919_n588# a_187_n588# 0.01fF
C256 a_n761_n588# a_n287_n588# 0.02fF
C257 a_187_n588# a_n1235_n588# 0.01fF
C258 a_29_n588# a_n919_n588# 0.01fF
C259 a_n445_n588# a_n1077_n588# 0.02fF
C260 a_29_n588# a_n1235_n588# 0.01fF
C261 a_n129_n588# a_n1077_n588# 0.01fF
C262 a_n445_n588# a_n761_n588# 0.04fF
C263 a_n287_n588# a_n1235_n588# 0.01fF
C264 a_n919_n588# a_n287_n588# 0.02fF
C265 a_n129_n588# a_n761_n588# 0.02fF
C266 a_n445_n588# a_n1235_n588# 0.01fF
C267 a_n919_n588# a_n445_n588# 0.02fF
C268 a_n129_n588# a_n1235_n588# 0.01fF
C269 a_n919_n588# a_n129_n588# 0.01fF
C270 a_n603_n588# a_n1077_n588# 0.02fF
C271 a_n761_n588# a_n603_n588# 0.12fF
C272 a_n603_n588# a_n1235_n588# 0.02fF
C273 a_n919_n588# a_n603_n588# 0.04fF
C274 a_n761_n588# a_n1077_n588# 0.04fF
C275 a_n1077_n588# a_n1235_n588# 0.12fF
C276 a_n919_n588# a_n1077_n588# 0.12fF
C277 a_n761_n588# a_n1235_n588# 0.02fF
C278 a_n919_n588# a_n761_n588# 0.12fF
C279 a_n919_n588# a_n1235_n588# 0.04fF
C280 a_n1393_n588# a_187_n588# 0.01fF
C281 a_29_n588# a_n1393_n588# 0.01fF
C282 a_n1393_n588# a_n287_n588# 0.01fF
C283 a_n445_n588# a_n1393_n588# 0.01fF
C284 a_n129_n588# a_n1393_n588# 0.01fF
C285 a_29_n588# a_n1551_n588# 0.01fF
C286 a_n1551_n588# a_n287_n588# 0.01fF
C287 a_n445_n588# a_n1551_n588# 0.01fF
C288 a_n1551_n588# a_n129_n588# 0.01fF
C289 a_n1393_n588# a_n603_n588# 0.01fF
C290 a_n1551_n588# a_n603_n588# 0.01fF
C291 a_n1393_n588# a_n1077_n588# 0.04fF
C292 a_n1393_n588# a_n761_n588# 0.02fF
C293 a_n1393_n588# a_n1235_n588# 0.12fF
C294 a_n919_n588# a_n1393_n588# 0.02fF
C295 a_n1551_n588# a_n1077_n588# 0.02fF
C296 a_n1551_n588# a_n761_n588# 0.01fF
C297 a_n919_n588# a_n1551_n588# 0.02fF
C298 a_n1551_n588# a_n1235_n588# 0.04fF
C299 a_n1551_n588# a_n1393_n588# 0.12fF
C300 a_1551_n500# a_n1743_n722# 0.30fF
C301 a_1393_n500# a_n1743_n722# 0.13fF
C302 a_1235_n500# a_n1743_n722# 0.09fF
C303 a_1077_n500# a_n1743_n722# 0.07fF
C304 a_919_n500# a_n1743_n722# 0.06fF
C305 a_761_n500# a_n1743_n722# 0.05fF
C306 a_603_n500# a_n1743_n722# 0.05fF
C307 a_445_n500# a_n1743_n722# 0.04fF
C308 a_287_n500# a_n1743_n722# 0.04fF
C309 a_129_n500# a_n1743_n722# 0.04fF
C310 a_n29_n500# a_n1743_n722# 0.02fF
C311 a_n187_n500# a_n1743_n722# 0.04fF
C312 a_n345_n500# a_n1743_n722# 0.04fF
C313 a_n503_n500# a_n1743_n722# 0.04fF
C314 a_n661_n500# a_n1743_n722# 0.05fF
C315 a_n819_n500# a_n1743_n722# 0.05fF
C316 a_n977_n500# a_n1743_n722# 0.06fF
C317 a_n1135_n500# a_n1743_n722# 0.07fF
C318 a_n1293_n500# a_n1743_n722# 0.09fF
C319 a_n1451_n500# a_n1743_n722# 0.13fF
C320 a_n1609_n500# a_n1743_n722# 0.30fF
C321 a_1451_n588# a_n1743_n722# 0.28fF
C322 a_1293_n588# a_n1743_n722# 0.23fF
C323 a_1135_n588# a_n1743_n722# 0.24fF
C324 a_977_n588# a_n1743_n722# 0.25fF
C325 a_819_n588# a_n1743_n722# 0.26fF
C326 a_661_n588# a_n1743_n722# 0.26fF
C327 a_503_n588# a_n1743_n722# 0.27fF
C328 a_345_n588# a_n1743_n722# 0.28fF
C329 a_187_n588# a_n1743_n722# 0.28fF
C330 a_29_n588# a_n1743_n722# 0.28fF
C331 a_n129_n588# a_n1743_n722# 0.28fF
C332 a_n287_n588# a_n1743_n722# 0.28fF
C333 a_n445_n588# a_n1743_n722# 0.28fF
C334 a_n603_n588# a_n1743_n722# 0.28fF
C335 a_n761_n588# a_n1743_n722# 0.28fF
C336 a_n919_n588# a_n1743_n722# 0.28fF
C337 a_n1077_n588# a_n1743_n722# 0.28fF
C338 a_n1235_n588# a_n1743_n722# 0.29fF
C339 a_n1393_n588# a_n1743_n722# 0.29fF
C340 a_n1551_n588# a_n1743_n722# 0.34fF
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_CADZ46 a_n345_n500# a_n1609_n500# a_n1135_n500#
+ a_29_n597# a_n977_n500# a_n129_n597# a_187_n597# a_n503_n500# a_129_n500# a_n1293_n500#
+ a_n287_n597# a_819_n597# a_n1077_n597# a_287_n500# a_n661_n500# a_345_n597# a_n919_n597#
+ a_n1451_n500# a_977_n597# a_n445_n597# a_919_n500# a_n1235_n597# a_445_n500# a_503_n597#
+ w_n1809_n797# a_n603_n597# a_1077_n500# a_1135_n597# a_661_n597# a_n1393_n597# a_603_n500#
+ a_1293_n597# a_n761_n597# a_1235_n500# a_n1551_n597# a_761_n500# a_n29_n500# a_1451_n597#
+ a_1393_n500# a_n187_n500# a_1551_n500# a_n819_n500# VSUBS
X0 a_n819_n500# a_n919_n597# a_n977_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X1 a_n661_n500# a_n761_n597# a_n819_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X2 a_919_n500# a_819_n597# a_761_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X3 a_n187_n500# a_n287_n597# a_n345_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X4 a_761_n500# a_661_n597# a_603_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X5 a_287_n500# a_187_n597# a_129_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X6 a_n1293_n500# a_n1393_n597# a_n1451_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X7 a_1393_n500# a_1293_n597# a_1235_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X8 a_n345_n500# a_n445_n597# a_n503_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X9 a_129_n500# a_29_n597# a_n29_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X10 a_445_n500# a_345_n597# a_287_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X11 a_n1451_n500# a_n1551_n597# a_n1609_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X12 a_1551_n500# a_1451_n597# a_1393_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X13 a_n977_n500# a_n1077_n597# a_n1135_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X14 a_1077_n500# a_977_n597# a_919_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X15 a_n503_n500# a_n603_n597# a_n661_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X16 a_n29_n500# a_n129_n597# a_n187_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X17 a_603_n500# a_503_n597# a_445_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X18 a_n1135_n500# a_n1235_n597# a_n1293_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X19 a_1235_n500# a_1135_n597# a_1077_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
C0 a_1393_n500# a_1551_n500# 0.56fF
C1 w_n1809_n797# a_1551_n500# 0.30fF
C2 w_n1809_n797# a_1393_n500# 0.13fF
C3 w_n1809_n797# a_n1551_n597# 0.30fF
C4 w_n1809_n797# a_n1393_n597# 0.25fF
C5 a_n1551_n597# a_n1393_n597# 0.12fF
C6 a_n1235_n597# w_n1809_n797# 0.24fF
C7 a_n1235_n597# a_n1551_n597# 0.04fF
C8 a_n1235_n597# a_n1393_n597# 0.12fF
C9 w_n1809_n797# a_n919_n597# 0.24fF
C10 a_n1551_n597# a_n919_n597# 0.02fF
C11 a_n1393_n597# a_n919_n597# 0.02fF
C12 w_n1809_n797# a_n1077_n597# 0.24fF
C13 a_n1551_n597# a_n1077_n597# 0.02fF
C14 a_n1077_n597# a_n1393_n597# 0.04fF
C15 w_n1809_n797# a_n761_n597# 0.24fF
C16 a_n761_n597# a_n1393_n597# 0.02fF
C17 a_n1551_n597# a_n761_n597# 0.01fF
C18 w_n1809_n797# a_n603_n597# 0.24fF
C19 a_n287_n597# w_n1809_n797# 0.24fF
C20 a_n1551_n597# a_n603_n597# 0.01fF
C21 a_n287_n597# a_n1551_n597# 0.01fF
C22 a_n1393_n597# a_n603_n597# 0.01fF
C23 w_n1809_n797# a_n445_n597# 0.24fF
C24 a_n287_n597# a_n1393_n597# 0.01fF
C25 a_n1235_n597# a_n919_n597# 0.04fF
C26 a_n1551_n597# a_n445_n597# 0.01fF
C27 a_n445_n597# a_n1393_n597# 0.01fF
C28 a_n1235_n597# a_n1077_n597# 0.12fF
C29 w_n1809_n797# a_29_n597# 0.24fF
C30 w_n1809_n797# a_n129_n597# 0.24fF
C31 a_n1551_n597# a_29_n597# 0.01fF
C32 a_29_n597# a_n1393_n597# 0.01fF
C33 a_n1235_n597# a_n761_n597# 0.02fF
C34 a_n1551_n597# a_n129_n597# 0.01fF
C35 a_n129_n597# a_n1393_n597# 0.01fF
C36 a_n1077_n597# a_n919_n597# 0.12fF
C37 w_n1809_n797# a_187_n597# 0.24fF
C38 a_n1235_n597# a_n287_n597# 0.01fF
C39 a_n761_n597# a_n919_n597# 0.12fF
C40 a_n1393_n597# a_187_n597# 0.01fF
C41 a_n1235_n597# a_n603_n597# 0.02fF
C42 a_345_n597# w_n1809_n797# 0.23fF
C43 a_n1077_n597# a_n761_n597# 0.04fF
C44 a_n1235_n597# a_n445_n597# 0.01fF
C45 w_n1809_n797# a_503_n597# 0.23fF
C46 a_n603_n597# a_n919_n597# 0.04fF
C47 a_n287_n597# a_n919_n597# 0.02fF
C48 a_n1235_n597# a_29_n597# 0.01fF
C49 a_n1077_n597# a_n603_n597# 0.02fF
C50 a_n445_n597# a_n919_n597# 0.02fF
C51 a_n1235_n597# a_n129_n597# 0.01fF
C52 a_n287_n597# a_n1077_n597# 0.01fF
C53 a_n1077_n597# a_n445_n597# 0.02fF
C54 a_n761_n597# a_n603_n597# 0.12fF
C55 a_29_n597# a_n919_n597# 0.01fF
C56 a_n287_n597# a_n761_n597# 0.02fF
C57 a_n1235_n597# a_187_n597# 0.01fF
C58 w_n1809_n797# a_819_n597# 0.21fF
C59 a_n129_n597# a_n919_n597# 0.01fF
C60 w_n1809_n797# a_661_n597# 0.22fF
C61 a_n761_n597# a_n445_n597# 0.04fF
C62 a_n1077_n597# a_29_n597# 0.01fF
C63 a_n1077_n597# a_n129_n597# 0.01fF
C64 a_345_n597# a_n1235_n597# 0.01fF
C65 a_n287_n597# a_n603_n597# 0.04fF
C66 a_n919_n597# a_187_n597# 0.01fF
C67 a_29_n597# a_n761_n597# 0.01fF
C68 a_n761_n597# a_n129_n597# 0.02fF
C69 a_n445_n597# a_n603_n597# 0.12fF
C70 a_n1077_n597# a_187_n597# 0.01fF
C71 a_n287_n597# a_n445_n597# 0.12fF
C72 a_345_n597# a_n919_n597# 0.01fF
C73 a_n761_n597# a_187_n597# 0.01fF
C74 a_29_n597# a_n603_n597# 0.02fF
C75 a_345_n597# a_n1077_n597# 0.01fF
C76 a_n287_n597# a_29_n597# 0.04fF
C77 a_n129_n597# a_n603_n597# 0.02fF
C78 a_503_n597# a_n919_n597# 0.01fF
C79 a_n287_n597# a_n129_n597# 0.12fF
C80 a_29_n597# a_n445_n597# 0.02fF
C81 a_n1077_n597# a_503_n597# 0.01fF
C82 a_345_n597# a_n761_n597# 0.01fF
C83 a_n129_n597# a_n445_n597# 0.04fF
C84 a_n603_n597# a_187_n597# 0.01fF
C85 a_n287_n597# a_187_n597# 0.02fF
C86 w_n1809_n797# a_977_n597# 0.20fF
C87 a_1135_n597# w_n1809_n797# 0.20fF
C88 a_n761_n597# a_503_n597# 0.01fF
C89 a_n445_n597# a_187_n597# 0.02fF
C90 a_29_n597# a_n129_n597# 0.12fF
C91 w_n1809_n797# a_1293_n597# 0.19fF
C92 a_345_n597# a_n603_n597# 0.01fF
C93 a_661_n597# a_n919_n597# 0.01fF
C94 a_345_n597# a_n287_n597# 0.02fF
C95 a_29_n597# a_187_n597# 0.12fF
C96 a_n603_n597# a_503_n597# 0.01fF
C97 a_345_n597# a_n445_n597# 0.01fF
C98 w_n1809_n797# a_n1609_n500# 0.30fF
C99 a_n129_n597# a_187_n597# 0.04fF
C100 a_n287_n597# a_503_n597# 0.01fF
C101 a_n445_n597# a_503_n597# 0.01fF
C102 a_n761_n597# a_819_n597# 0.01fF
C103 w_n1809_n797# a_n1451_n500# 0.13fF
C104 a_661_n597# a_n761_n597# 0.01fF
C105 a_345_n597# a_29_n597# 0.04fF
C106 w_n1809_n797# a_1451_n597# 0.24fF
C107 a_345_n597# a_n129_n597# 0.02fF
C108 a_29_n597# a_503_n597# 0.02fF
C109 w_n1809_n797# a_n1293_n500# 0.09fF
C110 a_n129_n597# a_503_n597# 0.02fF
C111 a_n603_n597# a_819_n597# 0.01fF
C112 a_n287_n597# a_819_n597# 0.01fF
C113 a_661_n597# a_n603_n597# 0.01fF
C114 a_345_n597# a_187_n597# 0.12fF
C115 a_n287_n597# a_661_n597# 0.01fF
C116 a_n445_n597# a_819_n597# 0.01fF
C117 a_661_n597# a_n445_n597# 0.01fF
C118 a_503_n597# a_187_n597# 0.04fF
C119 w_n1809_n797# a_n1135_n500# 0.07fF
C120 w_n1809_n797# a_n977_n500# 0.06fF
C121 a_29_n597# a_819_n597# 0.01fF
C122 a_29_n597# a_661_n597# 0.02fF
C123 a_n129_n597# a_819_n597# 0.01fF
C124 a_661_n597# a_n129_n597# 0.01fF
C125 a_345_n597# a_503_n597# 0.12fF
C126 a_661_n597# a_187_n597# 0.02fF
C127 a_819_n597# a_187_n597# 0.02fF
C128 a_345_n597# a_819_n597# 0.02fF
C129 a_345_n597# a_661_n597# 0.04fF
C130 a_977_n597# a_n603_n597# 0.01fF
C131 w_n1809_n797# a_n819_n500# 0.05fF
C132 a_n287_n597# a_977_n597# 0.01fF
C133 a_1135_n597# a_n287_n597# 0.01fF
C134 a_503_n597# a_819_n597# 0.04fF
C135 a_n287_n597# a_1293_n597# 0.01fF
C136 a_661_n597# a_503_n597# 0.12fF
C137 a_977_n597# a_n445_n597# 0.01fF
C138 a_1551_n500# a_n29_n500# 0.04fF
C139 a_1135_n597# a_n445_n597# 0.01fF
C140 w_n1809_n797# a_n661_n500# 0.05fF
C141 a_129_n500# a_1551_n500# 0.05fF
C142 a_29_n597# a_977_n597# 0.01fF
C143 a_977_n597# a_n129_n597# 0.01fF
C144 a_1135_n597# a_29_n597# 0.01fF
C145 a_29_n597# a_1293_n597# 0.01fF
C146 a_1135_n597# a_n129_n597# 0.01fF
C147 a_1393_n500# a_n29_n500# 0.05fF
C148 a_n129_n597# a_1293_n597# 0.01fF
C149 a_287_n500# a_1551_n500# 0.05fF
C150 w_n1809_n797# a_n503_n500# 0.04fF
C151 a_661_n597# a_819_n597# 0.12fF
C152 a_129_n500# a_1393_n500# 0.05fF
C153 a_n345_n500# w_n1809_n797# 0.04fF
C154 a_977_n597# a_187_n597# 0.01fF
C155 w_n1809_n797# a_n29_n500# 0.02fF
C156 a_n187_n500# a_1393_n500# 0.04fF
C157 a_1135_n597# a_187_n597# 0.01fF
C158 a_129_n500# w_n1809_n797# 0.04fF
C159 a_1551_n500# a_761_n500# 0.09fF
C160 a_1293_n597# a_187_n597# 0.01fF
C161 w_n1809_n797# a_n187_n500# 0.04fF
C162 a_445_n500# a_1551_n500# 0.06fF
C163 a_1393_n500# a_287_n500# 0.06fF
C164 a_345_n597# a_977_n597# 0.02fF
C165 a_1551_n500# a_919_n500# 0.11fF
C166 a_603_n500# a_1551_n500# 0.07fF
C167 a_29_n597# a_1451_n597# 0.01fF
C168 a_1135_n597# a_345_n597# 0.01fF
C169 a_345_n597# a_1293_n597# 0.01fF
C170 a_n129_n597# a_1451_n597# 0.01fF
C171 w_n1809_n797# a_287_n500# 0.04fF
C172 a_977_n597# a_503_n597# 0.02fF
C173 a_1135_n597# a_503_n597# 0.02fF
C174 a_1393_n500# a_761_n500# 0.11fF
C175 a_1293_n597# a_503_n597# 0.01fF
C176 a_1393_n500# a_445_n500# 0.07fF
C177 a_1451_n597# a_187_n597# 0.01fF
C178 w_n1809_n797# a_761_n500# 0.05fF
C179 a_1393_n500# a_919_n500# 0.15fF
C180 a_603_n500# a_1393_n500# 0.09fF
C181 w_n1809_n797# a_445_n500# 0.04fF
C182 a_603_n500# w_n1809_n797# 0.05fF
C183 w_n1809_n797# a_919_n500# 0.06fF
C184 a_977_n597# a_819_n597# 0.12fF
C185 a_345_n597# a_1451_n597# 0.01fF
C186 a_977_n597# a_661_n597# 0.04fF
C187 a_1135_n597# a_819_n597# 0.04fF
C188 a_1135_n597# a_661_n597# 0.02fF
C189 a_1293_n597# a_819_n597# 0.02fF
C190 a_661_n597# a_1293_n597# 0.02fF
C191 a_1451_n597# a_503_n597# 0.01fF
C192 a_1077_n500# a_1551_n500# 0.15fF
C193 a_1451_n597# a_819_n597# 0.02fF
C194 a_1235_n500# a_1551_n500# 0.24fF
C195 a_661_n597# a_1451_n597# 0.01fF
C196 a_1393_n500# a_1077_n500# 0.24fF
C197 w_n1809_n797# a_1077_n500# 0.07fF
C198 a_1235_n500# a_1393_n500# 0.56fF
C199 a_1135_n597# a_977_n597# 0.12fF
C200 a_977_n597# a_1293_n597# 0.04fF
C201 a_1235_n500# w_n1809_n797# 0.09fF
C202 a_1135_n597# a_1293_n597# 0.12fF
C203 a_977_n597# a_1451_n597# 0.02fF
C204 a_1135_n597# a_1451_n597# 0.04fF
C205 a_1293_n597# a_1451_n597# 0.12fF
C206 a_n1451_n500# a_n1609_n500# 0.56fF
C207 a_n1609_n500# a_n1293_n500# 0.24fF
C208 a_n1451_n500# a_n1293_n500# 0.56fF
C209 a_n1609_n500# a_n1135_n500# 0.15fF
C210 a_n1451_n500# a_n1135_n500# 0.24fF
C211 a_n1609_n500# a_n977_n500# 0.11fF
C212 a_n1451_n500# a_n977_n500# 0.15fF
C213 a_n1293_n500# a_n1135_n500# 0.56fF
C214 a_n977_n500# a_n1293_n500# 0.24fF
C215 a_n977_n500# a_n1135_n500# 0.56fF
C216 a_n1609_n500# a_n819_n500# 0.09fF
C217 a_n1451_n500# a_n819_n500# 0.11fF
C218 a_n1609_n500# a_n661_n500# 0.07fF
C219 a_n1451_n500# a_n661_n500# 0.09fF
C220 a_n819_n500# a_n1293_n500# 0.15fF
C221 a_n661_n500# a_n1293_n500# 0.11fF
C222 a_n1609_n500# a_n503_n500# 0.06fF
C223 a_n819_n500# a_n1135_n500# 0.24fF
C224 a_n345_n500# a_n1609_n500# 0.05fF
C225 a_n1609_n500# a_n29_n500# 0.04fF
C226 a_n1451_n500# a_n503_n500# 0.07fF
C227 a_n345_n500# a_n1451_n500# 0.06fF
C228 a_n977_n500# a_n819_n500# 0.56fF
C229 a_n187_n500# a_n1609_n500# 0.05fF
C230 a_n1451_n500# a_n29_n500# 0.05fF
C231 a_129_n500# a_n1451_n500# 0.04fF
C232 a_n661_n500# a_n1135_n500# 0.15fF
C233 a_n187_n500# a_n1451_n500# 0.05fF
C234 a_n1293_n500# a_n503_n500# 0.09fF
C235 a_n345_n500# a_n1293_n500# 0.07fF
C236 a_n977_n500# a_n661_n500# 0.24fF
C237 a_n1293_n500# a_n29_n500# 0.05fF
C238 a_129_n500# a_n1293_n500# 0.05fF
C239 a_n187_n500# a_n1293_n500# 0.06fF
C240 a_n503_n500# a_n1135_n500# 0.11fF
C241 a_n345_n500# a_n1135_n500# 0.09fF
C242 a_n29_n500# a_n1135_n500# 0.06fF
C243 a_n977_n500# a_n503_n500# 0.15fF
C244 a_287_n500# a_n1293_n500# 0.04fF
C245 a_n345_n500# a_n977_n500# 0.11fF
C246 a_129_n500# a_n1135_n500# 0.05fF
C247 a_n187_n500# a_n1135_n500# 0.07fF
C248 a_n977_n500# a_n29_n500# 0.07fF
C249 a_129_n500# a_n977_n500# 0.06fF
C250 a_n187_n500# a_n977_n500# 0.09fF
C251 a_n819_n500# a_n661_n500# 0.56fF
C252 a_287_n500# a_n1135_n500# 0.05fF
C253 a_287_n500# a_n977_n500# 0.05fF
C254 a_445_n500# a_n1135_n500# 0.04fF
C255 a_n819_n500# a_n503_n500# 0.24fF
C256 a_n345_n500# a_n819_n500# 0.15fF
C257 a_n819_n500# a_n29_n500# 0.09fF
C258 a_445_n500# a_n977_n500# 0.05fF
C259 a_129_n500# a_n819_n500# 0.07fF
C260 a_603_n500# a_n977_n500# 0.04fF
C261 a_n187_n500# a_n819_n500# 0.11fF
C262 a_n661_n500# a_n503_n500# 0.56fF
C263 a_n345_n500# a_n661_n500# 0.24fF
C264 a_n661_n500# a_n29_n500# 0.11fF
C265 a_287_n500# a_n819_n500# 0.06fF
C266 a_129_n500# a_n661_n500# 0.09fF
C267 a_n187_n500# a_n661_n500# 0.15fF
C268 a_n345_n500# a_n503_n500# 0.56fF
C269 a_n503_n500# a_n29_n500# 0.15fF
C270 a_287_n500# a_n661_n500# 0.07fF
C271 a_n819_n500# a_761_n500# 0.04fF
C272 a_n345_n500# a_n29_n500# 0.24fF
C273 a_445_n500# a_n819_n500# 0.05fF
C274 a_129_n500# a_n503_n500# 0.11fF
C275 a_n187_n500# a_n503_n500# 0.24fF
C276 a_603_n500# a_n819_n500# 0.05fF
C277 a_n345_n500# a_129_n500# 0.15fF
C278 a_n345_n500# a_n187_n500# 0.56fF
C279 a_129_n500# a_n29_n500# 0.56fF
C280 a_n187_n500# a_n29_n500# 0.56fF
C281 a_n661_n500# a_761_n500# 0.05fF
C282 a_445_n500# a_n661_n500# 0.06fF
C283 a_129_n500# a_n187_n500# 0.24fF
C284 a_287_n500# a_n503_n500# 0.09fF
C285 a_n661_n500# a_919_n500# 0.04fF
C286 a_n345_n500# a_287_n500# 0.11fF
C287 a_603_n500# a_n661_n500# 0.05fF
C288 a_287_n500# a_n29_n500# 0.24fF
C289 a_129_n500# a_287_n500# 0.56fF
C290 a_n187_n500# a_287_n500# 0.15fF
C291 a_761_n500# a_n503_n500# 0.05fF
C292 a_445_n500# a_n503_n500# 0.07fF
C293 a_n345_n500# a_761_n500# 0.06fF
C294 a_n345_n500# a_445_n500# 0.09fF
C295 a_761_n500# a_n29_n500# 0.09fF
C296 a_603_n500# a_n503_n500# 0.06fF
C297 a_445_n500# a_n29_n500# 0.15fF
C298 a_n345_n500# a_603_n500# 0.07fF
C299 a_129_n500# a_761_n500# 0.11fF
C300 a_n503_n500# a_919_n500# 0.05fF
C301 a_129_n500# a_445_n500# 0.24fF
C302 a_n187_n500# a_761_n500# 0.07fF
C303 a_n345_n500# a_919_n500# 0.05fF
C304 a_n29_n500# a_919_n500# 0.07fF
C305 a_603_n500# a_n29_n500# 0.11fF
C306 a_n187_n500# a_445_n500# 0.11fF
C307 a_129_n500# a_919_n500# 0.09fF
C308 a_603_n500# a_129_n500# 0.15fF
C309 a_n187_n500# a_919_n500# 0.06fF
C310 a_603_n500# a_n187_n500# 0.09fF
C311 a_287_n500# a_761_n500# 0.15fF
C312 a_445_n500# a_287_n500# 0.56fF
C313 a_603_n500# a_287_n500# 0.24fF
C314 a_287_n500# a_919_n500# 0.11fF
C315 a_445_n500# a_761_n500# 0.24fF
C316 a_761_n500# a_919_n500# 0.56fF
C317 a_603_n500# a_761_n500# 0.56fF
C318 a_603_n500# a_445_n500# 0.56fF
C319 a_445_n500# a_919_n500# 0.15fF
C320 a_603_n500# a_919_n500# 0.24fF
C321 a_1077_n500# a_n503_n500# 0.04fF
C322 a_n345_n500# a_1077_n500# 0.05fF
C323 a_1077_n500# a_n29_n500# 0.06fF
C324 a_129_n500# a_1077_n500# 0.07fF
C325 a_n187_n500# a_1077_n500# 0.05fF
C326 a_n345_n500# a_1235_n500# 0.04fF
C327 a_1235_n500# a_n29_n500# 0.05fF
C328 a_129_n500# a_1235_n500# 0.06fF
C329 a_1235_n500# a_n187_n500# 0.05fF
C330 a_1077_n500# a_287_n500# 0.09fF
C331 a_1235_n500# a_287_n500# 0.07fF
C332 a_1077_n500# a_761_n500# 0.24fF
C333 a_1077_n500# a_445_n500# 0.11fF
C334 a_603_n500# a_1077_n500# 0.15fF
C335 a_1077_n500# a_919_n500# 0.56fF
C336 a_1235_n500# a_761_n500# 0.15fF
C337 a_1235_n500# a_445_n500# 0.09fF
C338 a_603_n500# a_1235_n500# 0.11fF
C339 a_1235_n500# a_919_n500# 0.24fF
C340 a_1235_n500# a_1077_n500# 0.56fF
C341 w_n1809_n797# VSUBS 17.30fF
.ends

.subckt esd_cell esd VDD VSS
Xsky130_fd_pr__nfet_g5v0d10v5_BRTJC6_0 VSS VSS VSS VSS VSS VSS esd VSS VSS VSS esd
+ VSS esd VSS VSS VSS VSS esd VSS esd esd VSS VSS VSS VSS VSS VSS esd VSS VSS VSS
+ VSS esd VSS VSS esd VSS VSS VSS VSS VSS esd sky130_fd_pr__nfet_g5v0d10v5_BRTJC6
Xsky130_fd_pr__pfet_g5v0d10v5_CADZ46_0 VDD VDD esd VDD VDD VDD VDD esd esd VDD VDD
+ VDD VDD VDD VDD VDD VDD esd VDD VDD VDD VDD esd VDD VDD VDD esd VDD VDD VDD VDD
+ VDD VDD VDD VDD esd VDD VDD esd esd VDD esd VSS sky130_fd_pr__pfet_g5v0d10v5_CADZ46
C0 esd VDD 7.39fF
C1 VDD VSS -181.47fF
C2 esd VSS 8.04fF
.ends

