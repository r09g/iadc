magic
tech sky130A
magscale 1 2
timestamp 1654727055
<< nwell >>
rect -2386 -1864 -1092 -530
rect -589 -1479 -145 -913
rect 285 -1180 3100 -530
rect 285 -2514 3100 -1864
<< pwell >>
rect 1553 -68 1809 -66
rect -2386 -530 -1092 -68
rect 285 -530 3100 -68
rect -430 -669 -396 -635
rect -417 -673 -396 -669
rect -548 -700 -462 -690
rect -417 -700 -231 -673
rect -548 -855 -231 -700
rect 1553 -1402 1809 -1400
rect -548 -1692 -231 -1537
rect -548 -1693 -429 -1692
rect -548 -1702 -462 -1693
rect -417 -1719 -231 -1692
rect -417 -1723 -396 -1719
rect -430 -1757 -396 -1723
rect -2386 -2326 -1092 -1864
rect 285 -1864 3100 -1402
<< nmos >>
rect -2186 -382 -2156 -278
rect -2090 -382 -2060 -278
rect -1994 -382 -1964 -278
rect -1898 -382 -1868 -278
rect -1802 -382 -1772 -278
rect -1706 -382 -1676 -278
rect -1610 -382 -1580 -278
rect -1514 -382 -1484 -278
rect -1418 -382 -1388 -278
rect -1322 -382 -1292 -278
rect 485 -382 515 -278
rect 581 -382 611 -278
rect 677 -382 707 -278
rect 773 -382 803 -278
rect 869 -382 899 -278
rect 965 -382 995 -278
rect 1061 -382 1091 -278
rect 1157 -382 1187 -278
rect 1253 -382 1283 -278
rect 1349 -382 1379 -278
rect 1661 -384 1691 -284
rect 2006 -382 2036 -278
rect 2102 -382 2132 -278
rect 2198 -382 2228 -278
rect 2294 -382 2324 -278
rect 2390 -382 2420 -278
rect 2486 -382 2516 -278
rect 2582 -382 2612 -278
rect 2678 -382 2708 -278
rect 2774 -382 2804 -278
rect 2870 -382 2900 -278
rect 485 -1716 515 -1612
rect 581 -1716 611 -1612
rect 677 -1716 707 -1612
rect 773 -1716 803 -1612
rect 869 -1716 899 -1612
rect 965 -1716 995 -1612
rect 1061 -1716 1091 -1612
rect 1157 -1716 1187 -1612
rect 1253 -1716 1283 -1612
rect 1349 -1716 1379 -1612
rect 1661 -1718 1691 -1618
rect 2006 -1716 2036 -1612
rect 2102 -1716 2132 -1612
rect 2198 -1716 2228 -1612
rect 2294 -1716 2324 -1612
rect 2390 -1716 2420 -1612
rect 2486 -1716 2516 -1612
rect 2582 -1716 2612 -1612
rect 2678 -1716 2708 -1612
rect 2774 -1716 2804 -1612
rect 2870 -1716 2900 -1612
rect -2186 -2116 -2156 -2012
rect -2090 -2116 -2060 -2012
rect -1994 -2116 -1964 -2012
rect -1898 -2116 -1868 -2012
rect -1802 -2116 -1772 -2012
rect -1706 -2116 -1676 -2012
rect -1610 -2116 -1580 -2012
rect -1514 -2116 -1484 -2012
rect -1418 -2116 -1388 -2012
rect -1322 -2116 -1292 -2012
<< scnmos >>
rect -339 -829 -309 -699
rect -339 -1693 -309 -1563
<< pmos >>
rect -2186 -960 -2156 -688
rect -2090 -960 -2060 -688
rect -1994 -960 -1964 -688
rect -1898 -960 -1868 -688
rect -1802 -960 -1772 -688
rect -1706 -960 -1676 -688
rect -1610 -960 -1580 -688
rect -1514 -960 -1484 -688
rect -1418 -960 -1388 -688
rect -1322 -960 -1292 -688
rect 485 -960 515 -688
rect 581 -960 611 -688
rect 677 -960 707 -688
rect 773 -960 803 -688
rect 869 -960 899 -688
rect 965 -960 995 -688
rect 1061 -960 1091 -688
rect 1157 -960 1187 -688
rect 1253 -960 1283 -688
rect 1349 -960 1379 -688
rect 2006 -960 2036 -688
rect 2102 -960 2132 -688
rect 2198 -960 2228 -688
rect 2294 -960 2324 -688
rect 2390 -960 2420 -688
rect 2486 -960 2516 -688
rect 2582 -960 2612 -688
rect 2678 -960 2708 -688
rect 2774 -960 2804 -688
rect 2870 -960 2900 -688
rect -2186 -1706 -2156 -1434
rect -2090 -1706 -2060 -1434
rect -1994 -1706 -1964 -1434
rect -1898 -1706 -1868 -1434
rect -1802 -1706 -1772 -1434
rect -1706 -1706 -1676 -1434
rect -1610 -1706 -1580 -1434
rect -1514 -1706 -1484 -1434
rect -1418 -1706 -1388 -1434
rect -1322 -1706 -1292 -1434
rect 485 -2294 515 -2022
rect 581 -2294 611 -2022
rect 677 -2294 707 -2022
rect 773 -2294 803 -2022
rect 869 -2294 899 -2022
rect 965 -2294 995 -2022
rect 1061 -2294 1091 -2022
rect 1157 -2294 1187 -2022
rect 1253 -2294 1283 -2022
rect 1349 -2294 1379 -2022
rect 2006 -2294 2036 -2022
rect 2102 -2294 2132 -2022
rect 2198 -2294 2228 -2022
rect 2294 -2294 2324 -2022
rect 2390 -2294 2420 -2022
rect 2486 -2294 2516 -2022
rect 2582 -2294 2612 -2022
rect 2678 -2294 2708 -2022
rect 2774 -2294 2804 -2022
rect 2870 -2294 2900 -2022
<< scpmoshvt >>
rect -339 -1149 -309 -949
rect -339 -1443 -309 -1243
<< ndiff >>
rect -2248 -290 -2186 -278
rect -2248 -370 -2236 -290
rect -2202 -370 -2186 -290
rect -2248 -382 -2186 -370
rect -2156 -290 -2090 -278
rect -2156 -370 -2140 -290
rect -2106 -370 -2090 -290
rect -2156 -382 -2090 -370
rect -2060 -290 -1994 -278
rect -2060 -370 -2044 -290
rect -2010 -370 -1994 -290
rect -2060 -382 -1994 -370
rect -1964 -290 -1898 -278
rect -1964 -370 -1948 -290
rect -1914 -370 -1898 -290
rect -1964 -382 -1898 -370
rect -1868 -290 -1802 -278
rect -1868 -370 -1852 -290
rect -1818 -370 -1802 -290
rect -1868 -382 -1802 -370
rect -1772 -290 -1706 -278
rect -1772 -370 -1756 -290
rect -1722 -370 -1706 -290
rect -1772 -382 -1706 -370
rect -1676 -290 -1610 -278
rect -1676 -370 -1660 -290
rect -1626 -370 -1610 -290
rect -1676 -382 -1610 -370
rect -1580 -290 -1514 -278
rect -1580 -370 -1564 -290
rect -1530 -370 -1514 -290
rect -1580 -382 -1514 -370
rect -1484 -290 -1418 -278
rect -1484 -370 -1468 -290
rect -1434 -370 -1418 -290
rect -1484 -382 -1418 -370
rect -1388 -290 -1322 -278
rect -1388 -370 -1372 -290
rect -1338 -370 -1322 -290
rect -1388 -382 -1322 -370
rect -1292 -290 -1230 -278
rect -1292 -370 -1276 -290
rect -1242 -370 -1230 -290
rect -1292 -382 -1230 -370
rect 423 -290 485 -278
rect 423 -370 435 -290
rect 469 -370 485 -290
rect 423 -382 485 -370
rect 515 -290 581 -278
rect 515 -370 531 -290
rect 565 -370 581 -290
rect 515 -382 581 -370
rect 611 -290 677 -278
rect 611 -370 627 -290
rect 661 -370 677 -290
rect 611 -382 677 -370
rect 707 -290 773 -278
rect 707 -370 723 -290
rect 757 -370 773 -290
rect 707 -382 773 -370
rect 803 -290 869 -278
rect 803 -370 819 -290
rect 853 -370 869 -290
rect 803 -382 869 -370
rect 899 -290 965 -278
rect 899 -370 915 -290
rect 949 -370 965 -290
rect 899 -382 965 -370
rect 995 -290 1061 -278
rect 995 -370 1011 -290
rect 1045 -370 1061 -290
rect 995 -382 1061 -370
rect 1091 -290 1157 -278
rect 1091 -370 1107 -290
rect 1141 -370 1157 -290
rect 1091 -382 1157 -370
rect 1187 -290 1253 -278
rect 1187 -370 1203 -290
rect 1237 -370 1253 -290
rect 1187 -382 1253 -370
rect 1283 -290 1349 -278
rect 1283 -370 1299 -290
rect 1333 -370 1349 -290
rect 1283 -382 1349 -370
rect 1379 -290 1441 -278
rect 1379 -370 1395 -290
rect 1429 -370 1441 -290
rect 1379 -382 1441 -370
rect 1603 -296 1661 -284
rect 1603 -372 1615 -296
rect 1649 -372 1661 -296
rect 1603 -384 1661 -372
rect 1691 -296 1749 -284
rect 1691 -372 1703 -296
rect 1737 -372 1749 -296
rect 1691 -384 1749 -372
rect 1944 -290 2006 -278
rect 1944 -370 1956 -290
rect 1990 -370 2006 -290
rect 1944 -382 2006 -370
rect 2036 -290 2102 -278
rect 2036 -370 2052 -290
rect 2086 -370 2102 -290
rect 2036 -382 2102 -370
rect 2132 -290 2198 -278
rect 2132 -370 2148 -290
rect 2182 -370 2198 -290
rect 2132 -382 2198 -370
rect 2228 -290 2294 -278
rect 2228 -370 2244 -290
rect 2278 -370 2294 -290
rect 2228 -382 2294 -370
rect 2324 -290 2390 -278
rect 2324 -370 2340 -290
rect 2374 -370 2390 -290
rect 2324 -382 2390 -370
rect 2420 -290 2486 -278
rect 2420 -370 2436 -290
rect 2470 -370 2486 -290
rect 2420 -382 2486 -370
rect 2516 -290 2582 -278
rect 2516 -370 2532 -290
rect 2566 -370 2582 -290
rect 2516 -382 2582 -370
rect 2612 -290 2678 -278
rect 2612 -370 2628 -290
rect 2662 -370 2678 -290
rect 2612 -382 2678 -370
rect 2708 -290 2774 -278
rect 2708 -370 2724 -290
rect 2758 -370 2774 -290
rect 2708 -382 2774 -370
rect 2804 -290 2870 -278
rect 2804 -370 2820 -290
rect 2854 -370 2870 -290
rect 2804 -382 2870 -370
rect 2900 -290 2962 -278
rect 2900 -370 2916 -290
rect 2950 -370 2962 -290
rect 2900 -382 2962 -370
rect -391 -715 -339 -699
rect -391 -749 -383 -715
rect -349 -749 -339 -715
rect -391 -783 -339 -749
rect -391 -817 -383 -783
rect -349 -817 -339 -783
rect -391 -829 -339 -817
rect -309 -715 -257 -699
rect -309 -749 -299 -715
rect -265 -749 -257 -715
rect -309 -783 -257 -749
rect -309 -817 -299 -783
rect -265 -817 -257 -783
rect -309 -829 -257 -817
rect -391 -1575 -339 -1563
rect -391 -1609 -383 -1575
rect -349 -1609 -339 -1575
rect -391 -1643 -339 -1609
rect -391 -1677 -383 -1643
rect -349 -1677 -339 -1643
rect -391 -1693 -339 -1677
rect -309 -1575 -257 -1563
rect -309 -1609 -299 -1575
rect -265 -1609 -257 -1575
rect -309 -1643 -257 -1609
rect -309 -1677 -299 -1643
rect -265 -1677 -257 -1643
rect -309 -1693 -257 -1677
rect 423 -1624 485 -1612
rect 423 -1704 435 -1624
rect 469 -1704 485 -1624
rect 423 -1716 485 -1704
rect 515 -1624 581 -1612
rect 515 -1704 531 -1624
rect 565 -1704 581 -1624
rect 515 -1716 581 -1704
rect 611 -1624 677 -1612
rect 611 -1704 627 -1624
rect 661 -1704 677 -1624
rect 611 -1716 677 -1704
rect 707 -1624 773 -1612
rect 707 -1704 723 -1624
rect 757 -1704 773 -1624
rect 707 -1716 773 -1704
rect 803 -1624 869 -1612
rect 803 -1704 819 -1624
rect 853 -1704 869 -1624
rect 803 -1716 869 -1704
rect 899 -1624 965 -1612
rect 899 -1704 915 -1624
rect 949 -1704 965 -1624
rect 899 -1716 965 -1704
rect 995 -1624 1061 -1612
rect 995 -1704 1011 -1624
rect 1045 -1704 1061 -1624
rect 995 -1716 1061 -1704
rect 1091 -1624 1157 -1612
rect 1091 -1704 1107 -1624
rect 1141 -1704 1157 -1624
rect 1091 -1716 1157 -1704
rect 1187 -1624 1253 -1612
rect 1187 -1704 1203 -1624
rect 1237 -1704 1253 -1624
rect 1187 -1716 1253 -1704
rect 1283 -1624 1349 -1612
rect 1283 -1704 1299 -1624
rect 1333 -1704 1349 -1624
rect 1283 -1716 1349 -1704
rect 1379 -1624 1441 -1612
rect 1379 -1704 1395 -1624
rect 1429 -1704 1441 -1624
rect 1379 -1716 1441 -1704
rect 1603 -1630 1661 -1618
rect 1603 -1706 1615 -1630
rect 1649 -1706 1661 -1630
rect 1603 -1718 1661 -1706
rect 1691 -1630 1749 -1618
rect 1691 -1706 1703 -1630
rect 1737 -1706 1749 -1630
rect 1691 -1718 1749 -1706
rect 1944 -1624 2006 -1612
rect 1944 -1704 1956 -1624
rect 1990 -1704 2006 -1624
rect 1944 -1716 2006 -1704
rect 2036 -1624 2102 -1612
rect 2036 -1704 2052 -1624
rect 2086 -1704 2102 -1624
rect 2036 -1716 2102 -1704
rect 2132 -1624 2198 -1612
rect 2132 -1704 2148 -1624
rect 2182 -1704 2198 -1624
rect 2132 -1716 2198 -1704
rect 2228 -1624 2294 -1612
rect 2228 -1704 2244 -1624
rect 2278 -1704 2294 -1624
rect 2228 -1716 2294 -1704
rect 2324 -1624 2390 -1612
rect 2324 -1704 2340 -1624
rect 2374 -1704 2390 -1624
rect 2324 -1716 2390 -1704
rect 2420 -1624 2486 -1612
rect 2420 -1704 2436 -1624
rect 2470 -1704 2486 -1624
rect 2420 -1716 2486 -1704
rect 2516 -1624 2582 -1612
rect 2516 -1704 2532 -1624
rect 2566 -1704 2582 -1624
rect 2516 -1716 2582 -1704
rect 2612 -1624 2678 -1612
rect 2612 -1704 2628 -1624
rect 2662 -1704 2678 -1624
rect 2612 -1716 2678 -1704
rect 2708 -1624 2774 -1612
rect 2708 -1704 2724 -1624
rect 2758 -1704 2774 -1624
rect 2708 -1716 2774 -1704
rect 2804 -1624 2870 -1612
rect 2804 -1704 2820 -1624
rect 2854 -1704 2870 -1624
rect 2804 -1716 2870 -1704
rect 2900 -1624 2962 -1612
rect 2900 -1704 2916 -1624
rect 2950 -1704 2962 -1624
rect 2900 -1716 2962 -1704
rect -2248 -2024 -2186 -2012
rect -2248 -2104 -2236 -2024
rect -2202 -2104 -2186 -2024
rect -2248 -2116 -2186 -2104
rect -2156 -2024 -2090 -2012
rect -2156 -2104 -2140 -2024
rect -2106 -2104 -2090 -2024
rect -2156 -2116 -2090 -2104
rect -2060 -2024 -1994 -2012
rect -2060 -2104 -2044 -2024
rect -2010 -2104 -1994 -2024
rect -2060 -2116 -1994 -2104
rect -1964 -2024 -1898 -2012
rect -1964 -2104 -1948 -2024
rect -1914 -2104 -1898 -2024
rect -1964 -2116 -1898 -2104
rect -1868 -2024 -1802 -2012
rect -1868 -2104 -1852 -2024
rect -1818 -2104 -1802 -2024
rect -1868 -2116 -1802 -2104
rect -1772 -2024 -1706 -2012
rect -1772 -2104 -1756 -2024
rect -1722 -2104 -1706 -2024
rect -1772 -2116 -1706 -2104
rect -1676 -2024 -1610 -2012
rect -1676 -2104 -1660 -2024
rect -1626 -2104 -1610 -2024
rect -1676 -2116 -1610 -2104
rect -1580 -2024 -1514 -2012
rect -1580 -2104 -1564 -2024
rect -1530 -2104 -1514 -2024
rect -1580 -2116 -1514 -2104
rect -1484 -2024 -1418 -2012
rect -1484 -2104 -1468 -2024
rect -1434 -2104 -1418 -2024
rect -1484 -2116 -1418 -2104
rect -1388 -2024 -1322 -2012
rect -1388 -2104 -1372 -2024
rect -1338 -2104 -1322 -2024
rect -1388 -2116 -1322 -2104
rect -1292 -2024 -1230 -2012
rect -1292 -2104 -1276 -2024
rect -1242 -2104 -1230 -2024
rect -1292 -2116 -1230 -2104
<< pdiff >>
rect -2248 -700 -2186 -688
rect -2248 -948 -2236 -700
rect -2202 -948 -2186 -700
rect -2248 -960 -2186 -948
rect -2156 -700 -2090 -688
rect -2156 -948 -2140 -700
rect -2106 -948 -2090 -700
rect -2156 -960 -2090 -948
rect -2060 -700 -1994 -688
rect -2060 -948 -2044 -700
rect -2010 -948 -1994 -700
rect -2060 -960 -1994 -948
rect -1964 -700 -1898 -688
rect -1964 -948 -1948 -700
rect -1914 -948 -1898 -700
rect -1964 -960 -1898 -948
rect -1868 -700 -1802 -688
rect -1868 -948 -1852 -700
rect -1818 -948 -1802 -700
rect -1868 -960 -1802 -948
rect -1772 -700 -1706 -688
rect -1772 -948 -1756 -700
rect -1722 -948 -1706 -700
rect -1772 -960 -1706 -948
rect -1676 -700 -1610 -688
rect -1676 -948 -1660 -700
rect -1626 -948 -1610 -700
rect -1676 -960 -1610 -948
rect -1580 -700 -1514 -688
rect -1580 -948 -1564 -700
rect -1530 -948 -1514 -700
rect -1580 -960 -1514 -948
rect -1484 -700 -1418 -688
rect -1484 -948 -1468 -700
rect -1434 -948 -1418 -700
rect -1484 -960 -1418 -948
rect -1388 -700 -1322 -688
rect -1388 -948 -1372 -700
rect -1338 -948 -1322 -700
rect -1388 -960 -1322 -948
rect -1292 -700 -1230 -688
rect -1292 -948 -1276 -700
rect -1242 -948 -1230 -700
rect -1292 -960 -1230 -948
rect -391 -967 -339 -949
rect -391 -1001 -383 -967
rect -349 -1001 -339 -967
rect -391 -1035 -339 -1001
rect -391 -1069 -383 -1035
rect -349 -1069 -339 -1035
rect -391 -1103 -339 -1069
rect -391 -1137 -383 -1103
rect -349 -1137 -339 -1103
rect -391 -1149 -339 -1137
rect -309 -967 -257 -949
rect -309 -1001 -299 -967
rect -265 -1001 -257 -967
rect -309 -1035 -257 -1001
rect -309 -1069 -299 -1035
rect -265 -1069 -257 -1035
rect -309 -1103 -257 -1069
rect -309 -1137 -299 -1103
rect -265 -1137 -257 -1103
rect -309 -1149 -257 -1137
rect 423 -700 485 -688
rect 423 -948 435 -700
rect 469 -948 485 -700
rect 423 -960 485 -948
rect 515 -700 581 -688
rect 515 -948 531 -700
rect 565 -948 581 -700
rect 515 -960 581 -948
rect 611 -700 677 -688
rect 611 -948 627 -700
rect 661 -948 677 -700
rect 611 -960 677 -948
rect 707 -700 773 -688
rect 707 -948 723 -700
rect 757 -948 773 -700
rect 707 -960 773 -948
rect 803 -700 869 -688
rect 803 -948 819 -700
rect 853 -948 869 -700
rect 803 -960 869 -948
rect 899 -700 965 -688
rect 899 -948 915 -700
rect 949 -948 965 -700
rect 899 -960 965 -948
rect 995 -700 1061 -688
rect 995 -948 1011 -700
rect 1045 -948 1061 -700
rect 995 -960 1061 -948
rect 1091 -700 1157 -688
rect 1091 -948 1107 -700
rect 1141 -948 1157 -700
rect 1091 -960 1157 -948
rect 1187 -700 1253 -688
rect 1187 -948 1203 -700
rect 1237 -948 1253 -700
rect 1187 -960 1253 -948
rect 1283 -700 1349 -688
rect 1283 -948 1299 -700
rect 1333 -948 1349 -700
rect 1283 -960 1349 -948
rect 1379 -700 1441 -688
rect 1379 -948 1395 -700
rect 1429 -948 1441 -700
rect 1379 -960 1441 -948
rect 1944 -700 2006 -688
rect 1944 -948 1956 -700
rect 1990 -948 2006 -700
rect 1944 -960 2006 -948
rect 2036 -700 2102 -688
rect 2036 -948 2052 -700
rect 2086 -948 2102 -700
rect 2036 -960 2102 -948
rect 2132 -700 2198 -688
rect 2132 -948 2148 -700
rect 2182 -948 2198 -700
rect 2132 -960 2198 -948
rect 2228 -700 2294 -688
rect 2228 -948 2244 -700
rect 2278 -948 2294 -700
rect 2228 -960 2294 -948
rect 2324 -700 2390 -688
rect 2324 -948 2340 -700
rect 2374 -948 2390 -700
rect 2324 -960 2390 -948
rect 2420 -700 2486 -688
rect 2420 -948 2436 -700
rect 2470 -948 2486 -700
rect 2420 -960 2486 -948
rect 2516 -700 2582 -688
rect 2516 -948 2532 -700
rect 2566 -948 2582 -700
rect 2516 -960 2582 -948
rect 2612 -700 2678 -688
rect 2612 -948 2628 -700
rect 2662 -948 2678 -700
rect 2612 -960 2678 -948
rect 2708 -700 2774 -688
rect 2708 -948 2724 -700
rect 2758 -948 2774 -700
rect 2708 -960 2774 -948
rect 2804 -700 2870 -688
rect 2804 -948 2820 -700
rect 2854 -948 2870 -700
rect 2804 -960 2870 -948
rect 2900 -700 2962 -688
rect 2900 -948 2916 -700
rect 2950 -948 2962 -700
rect 2900 -960 2962 -948
rect -391 -1255 -339 -1243
rect -2248 -1446 -2186 -1434
rect -2248 -1694 -2236 -1446
rect -2202 -1694 -2186 -1446
rect -2248 -1706 -2186 -1694
rect -2156 -1446 -2090 -1434
rect -2156 -1694 -2140 -1446
rect -2106 -1694 -2090 -1446
rect -2156 -1706 -2090 -1694
rect -2060 -1446 -1994 -1434
rect -2060 -1694 -2044 -1446
rect -2010 -1694 -1994 -1446
rect -2060 -1706 -1994 -1694
rect -1964 -1446 -1898 -1434
rect -1964 -1694 -1948 -1446
rect -1914 -1694 -1898 -1446
rect -1964 -1706 -1898 -1694
rect -1868 -1446 -1802 -1434
rect -1868 -1694 -1852 -1446
rect -1818 -1694 -1802 -1446
rect -1868 -1706 -1802 -1694
rect -1772 -1446 -1706 -1434
rect -1772 -1694 -1756 -1446
rect -1722 -1694 -1706 -1446
rect -1772 -1706 -1706 -1694
rect -1676 -1446 -1610 -1434
rect -1676 -1694 -1660 -1446
rect -1626 -1694 -1610 -1446
rect -1676 -1706 -1610 -1694
rect -1580 -1446 -1514 -1434
rect -1580 -1694 -1564 -1446
rect -1530 -1694 -1514 -1446
rect -1580 -1706 -1514 -1694
rect -1484 -1446 -1418 -1434
rect -1484 -1694 -1468 -1446
rect -1434 -1694 -1418 -1446
rect -1484 -1706 -1418 -1694
rect -1388 -1446 -1322 -1434
rect -1388 -1694 -1372 -1446
rect -1338 -1694 -1322 -1446
rect -1388 -1706 -1322 -1694
rect -1292 -1446 -1230 -1434
rect -1292 -1694 -1276 -1446
rect -1242 -1694 -1230 -1446
rect -1292 -1706 -1230 -1694
rect -391 -1289 -383 -1255
rect -349 -1289 -339 -1255
rect -391 -1323 -339 -1289
rect -391 -1357 -383 -1323
rect -349 -1357 -339 -1323
rect -391 -1391 -339 -1357
rect -391 -1425 -383 -1391
rect -349 -1425 -339 -1391
rect -391 -1443 -339 -1425
rect -309 -1255 -257 -1243
rect -309 -1289 -299 -1255
rect -265 -1289 -257 -1255
rect -309 -1323 -257 -1289
rect -309 -1357 -299 -1323
rect -265 -1357 -257 -1323
rect -309 -1391 -257 -1357
rect -309 -1425 -299 -1391
rect -265 -1425 -257 -1391
rect -309 -1443 -257 -1425
rect 423 -2034 485 -2022
rect 423 -2282 435 -2034
rect 469 -2282 485 -2034
rect 423 -2294 485 -2282
rect 515 -2034 581 -2022
rect 515 -2282 531 -2034
rect 565 -2282 581 -2034
rect 515 -2294 581 -2282
rect 611 -2034 677 -2022
rect 611 -2282 627 -2034
rect 661 -2282 677 -2034
rect 611 -2294 677 -2282
rect 707 -2034 773 -2022
rect 707 -2282 723 -2034
rect 757 -2282 773 -2034
rect 707 -2294 773 -2282
rect 803 -2034 869 -2022
rect 803 -2282 819 -2034
rect 853 -2282 869 -2034
rect 803 -2294 869 -2282
rect 899 -2034 965 -2022
rect 899 -2282 915 -2034
rect 949 -2282 965 -2034
rect 899 -2294 965 -2282
rect 995 -2034 1061 -2022
rect 995 -2282 1011 -2034
rect 1045 -2282 1061 -2034
rect 995 -2294 1061 -2282
rect 1091 -2034 1157 -2022
rect 1091 -2282 1107 -2034
rect 1141 -2282 1157 -2034
rect 1091 -2294 1157 -2282
rect 1187 -2034 1253 -2022
rect 1187 -2282 1203 -2034
rect 1237 -2282 1253 -2034
rect 1187 -2294 1253 -2282
rect 1283 -2034 1349 -2022
rect 1283 -2282 1299 -2034
rect 1333 -2282 1349 -2034
rect 1283 -2294 1349 -2282
rect 1379 -2034 1441 -2022
rect 1379 -2282 1395 -2034
rect 1429 -2282 1441 -2034
rect 1379 -2294 1441 -2282
rect 1944 -2034 2006 -2022
rect 1944 -2282 1956 -2034
rect 1990 -2282 2006 -2034
rect 1944 -2294 2006 -2282
rect 2036 -2034 2102 -2022
rect 2036 -2282 2052 -2034
rect 2086 -2282 2102 -2034
rect 2036 -2294 2102 -2282
rect 2132 -2034 2198 -2022
rect 2132 -2282 2148 -2034
rect 2182 -2282 2198 -2034
rect 2132 -2294 2198 -2282
rect 2228 -2034 2294 -2022
rect 2228 -2282 2244 -2034
rect 2278 -2282 2294 -2034
rect 2228 -2294 2294 -2282
rect 2324 -2034 2390 -2022
rect 2324 -2282 2340 -2034
rect 2374 -2282 2390 -2034
rect 2324 -2294 2390 -2282
rect 2420 -2034 2486 -2022
rect 2420 -2282 2436 -2034
rect 2470 -2282 2486 -2034
rect 2420 -2294 2486 -2282
rect 2516 -2034 2582 -2022
rect 2516 -2282 2532 -2034
rect 2566 -2282 2582 -2034
rect 2516 -2294 2582 -2282
rect 2612 -2034 2678 -2022
rect 2612 -2282 2628 -2034
rect 2662 -2282 2678 -2034
rect 2612 -2294 2678 -2282
rect 2708 -2034 2774 -2022
rect 2708 -2282 2724 -2034
rect 2758 -2282 2774 -2034
rect 2708 -2294 2774 -2282
rect 2804 -2034 2870 -2022
rect 2804 -2282 2820 -2034
rect 2854 -2282 2870 -2034
rect 2804 -2294 2870 -2282
rect 2900 -2034 2962 -2022
rect 2900 -2282 2916 -2034
rect 2950 -2282 2962 -2034
rect 2900 -2294 2962 -2282
<< ndiffc >>
rect -2236 -370 -2202 -290
rect -2140 -370 -2106 -290
rect -2044 -370 -2010 -290
rect -1948 -370 -1914 -290
rect -1852 -370 -1818 -290
rect -1756 -370 -1722 -290
rect -1660 -370 -1626 -290
rect -1564 -370 -1530 -290
rect -1468 -370 -1434 -290
rect -1372 -370 -1338 -290
rect -1276 -370 -1242 -290
rect 435 -370 469 -290
rect 531 -370 565 -290
rect 627 -370 661 -290
rect 723 -370 757 -290
rect 819 -370 853 -290
rect 915 -370 949 -290
rect 1011 -370 1045 -290
rect 1107 -370 1141 -290
rect 1203 -370 1237 -290
rect 1299 -370 1333 -290
rect 1395 -370 1429 -290
rect 1615 -372 1649 -296
rect 1703 -372 1737 -296
rect 1956 -370 1990 -290
rect 2052 -370 2086 -290
rect 2148 -370 2182 -290
rect 2244 -370 2278 -290
rect 2340 -370 2374 -290
rect 2436 -370 2470 -290
rect 2532 -370 2566 -290
rect 2628 -370 2662 -290
rect 2724 -370 2758 -290
rect 2820 -370 2854 -290
rect 2916 -370 2950 -290
rect -383 -749 -349 -715
rect -383 -817 -349 -783
rect -299 -749 -265 -715
rect -299 -817 -265 -783
rect -383 -1609 -349 -1575
rect -383 -1677 -349 -1643
rect -299 -1609 -265 -1575
rect -299 -1677 -265 -1643
rect 435 -1704 469 -1624
rect 531 -1704 565 -1624
rect 627 -1704 661 -1624
rect 723 -1704 757 -1624
rect 819 -1704 853 -1624
rect 915 -1704 949 -1624
rect 1011 -1704 1045 -1624
rect 1107 -1704 1141 -1624
rect 1203 -1704 1237 -1624
rect 1299 -1704 1333 -1624
rect 1395 -1704 1429 -1624
rect 1615 -1706 1649 -1630
rect 1703 -1706 1737 -1630
rect 1956 -1704 1990 -1624
rect 2052 -1704 2086 -1624
rect 2148 -1704 2182 -1624
rect 2244 -1704 2278 -1624
rect 2340 -1704 2374 -1624
rect 2436 -1704 2470 -1624
rect 2532 -1704 2566 -1624
rect 2628 -1704 2662 -1624
rect 2724 -1704 2758 -1624
rect 2820 -1704 2854 -1624
rect 2916 -1704 2950 -1624
rect -2236 -2104 -2202 -2024
rect -2140 -2104 -2106 -2024
rect -2044 -2104 -2010 -2024
rect -1948 -2104 -1914 -2024
rect -1852 -2104 -1818 -2024
rect -1756 -2104 -1722 -2024
rect -1660 -2104 -1626 -2024
rect -1564 -2104 -1530 -2024
rect -1468 -2104 -1434 -2024
rect -1372 -2104 -1338 -2024
rect -1276 -2104 -1242 -2024
<< pdiffc >>
rect -2236 -948 -2202 -700
rect -2140 -948 -2106 -700
rect -2044 -948 -2010 -700
rect -1948 -948 -1914 -700
rect -1852 -948 -1818 -700
rect -1756 -948 -1722 -700
rect -1660 -948 -1626 -700
rect -1564 -948 -1530 -700
rect -1468 -948 -1434 -700
rect -1372 -948 -1338 -700
rect -1276 -948 -1242 -700
rect -383 -1001 -349 -967
rect -383 -1069 -349 -1035
rect -383 -1137 -349 -1103
rect -299 -1001 -265 -967
rect -299 -1069 -265 -1035
rect -299 -1137 -265 -1103
rect 435 -948 469 -700
rect 531 -948 565 -700
rect 627 -948 661 -700
rect 723 -948 757 -700
rect 819 -948 853 -700
rect 915 -948 949 -700
rect 1011 -948 1045 -700
rect 1107 -948 1141 -700
rect 1203 -948 1237 -700
rect 1299 -948 1333 -700
rect 1395 -948 1429 -700
rect 1956 -948 1990 -700
rect 2052 -948 2086 -700
rect 2148 -948 2182 -700
rect 2244 -948 2278 -700
rect 2340 -948 2374 -700
rect 2436 -948 2470 -700
rect 2532 -948 2566 -700
rect 2628 -948 2662 -700
rect 2724 -948 2758 -700
rect 2820 -948 2854 -700
rect 2916 -948 2950 -700
rect -2236 -1694 -2202 -1446
rect -2140 -1694 -2106 -1446
rect -2044 -1694 -2010 -1446
rect -1948 -1694 -1914 -1446
rect -1852 -1694 -1818 -1446
rect -1756 -1694 -1722 -1446
rect -1660 -1694 -1626 -1446
rect -1564 -1694 -1530 -1446
rect -1468 -1694 -1434 -1446
rect -1372 -1694 -1338 -1446
rect -1276 -1694 -1242 -1446
rect -383 -1289 -349 -1255
rect -383 -1357 -349 -1323
rect -383 -1425 -349 -1391
rect -299 -1289 -265 -1255
rect -299 -1357 -265 -1323
rect -299 -1425 -265 -1391
rect 435 -2282 469 -2034
rect 531 -2282 565 -2034
rect 627 -2282 661 -2034
rect 723 -2282 757 -2034
rect 819 -2282 853 -2034
rect 915 -2282 949 -2034
rect 1011 -2282 1045 -2034
rect 1107 -2282 1141 -2034
rect 1203 -2282 1237 -2034
rect 1299 -2282 1333 -2034
rect 1395 -2282 1429 -2034
rect 1956 -2282 1990 -2034
rect 2052 -2282 2086 -2034
rect 2148 -2282 2182 -2034
rect 2244 -2282 2278 -2034
rect 2340 -2282 2374 -2034
rect 2436 -2282 2470 -2034
rect 2532 -2282 2566 -2034
rect 2628 -2282 2662 -2034
rect 2724 -2282 2758 -2034
rect 2820 -2282 2854 -2034
rect 2916 -2282 2950 -2034
<< psubdiff >>
rect -2350 -138 -2254 -104
rect -1224 -138 -1128 -104
rect -2350 -200 -2316 -138
rect -1162 -200 -1128 -138
rect -2350 -460 -2316 -398
rect -1162 -460 -1128 -398
rect -2350 -494 -2254 -460
rect -1224 -494 -1128 -460
rect 321 -138 417 -104
rect 1447 -138 1543 -104
rect 321 -200 355 -138
rect 1509 -200 1543 -138
rect 321 -460 355 -398
rect 1842 -138 1938 -104
rect 2968 -138 3064 -104
rect 1842 -200 1876 -138
rect 1509 -460 1543 -398
rect 3030 -200 3064 -138
rect 321 -494 417 -460
rect 1447 -494 1543 -460
rect 1842 -460 1876 -398
rect 3030 -460 3064 -398
rect 1842 -494 1938 -460
rect 2968 -494 3064 -460
rect -522 -763 -488 -716
rect -522 -821 -488 -797
rect 321 -1472 417 -1438
rect 1447 -1472 1543 -1438
rect 321 -1534 355 -1472
rect -522 -1595 -488 -1571
rect -522 -1676 -488 -1629
rect 1509 -1534 1543 -1472
rect 321 -1794 355 -1732
rect 1842 -1472 1938 -1438
rect 2968 -1472 3064 -1438
rect 1842 -1534 1876 -1472
rect 1509 -1794 1543 -1732
rect 3030 -1534 3064 -1472
rect 321 -1828 417 -1794
rect 1447 -1828 1543 -1794
rect 1842 -1794 1876 -1732
rect 3030 -1794 3064 -1732
rect 1842 -1828 1938 -1794
rect 2968 -1828 3064 -1794
rect -2350 -1934 -2254 -1900
rect -1224 -1934 -1128 -1900
rect -2350 -1996 -2316 -1934
rect -1162 -1996 -1128 -1934
rect -2350 -2256 -2316 -2194
rect -1162 -2256 -1128 -2194
rect -2350 -2290 -2254 -2256
rect -1224 -2290 -1128 -2256
<< nsubdiff >>
rect -2350 -600 -2254 -566
rect -1224 -600 -1128 -566
rect -2350 -662 -2316 -600
rect -1162 -662 -1128 -600
rect -2350 -1110 -2316 -1048
rect 321 -600 417 -566
rect 1447 -600 1543 -566
rect 321 -662 355 -600
rect 1509 -662 1543 -600
rect -1162 -1110 -1128 -1048
rect -2350 -1144 -2254 -1110
rect -1224 -1144 -1128 -1110
rect -522 -981 -488 -957
rect -522 -1074 -488 -1015
rect -522 -1132 -488 -1108
rect 321 -1110 355 -1048
rect 1509 -1110 1543 -1048
rect 321 -1144 417 -1110
rect 1447 -1144 1543 -1110
rect 1842 -600 1938 -566
rect 2968 -600 3064 -566
rect 1842 -662 1876 -600
rect 3030 -662 3064 -600
rect 1842 -1110 1876 -1048
rect 3030 -1110 3064 -1048
rect 1842 -1144 1938 -1110
rect 2968 -1144 3064 -1110
rect -2350 -1284 -2254 -1250
rect -1224 -1284 -1128 -1250
rect -2350 -1346 -2316 -1284
rect -1162 -1346 -1128 -1284
rect -522 -1284 -488 -1260
rect -522 -1377 -488 -1318
rect -522 -1435 -488 -1411
rect -2350 -1794 -2316 -1732
rect -1162 -1794 -1128 -1732
rect -2350 -1828 -2254 -1794
rect -1224 -1828 -1128 -1794
rect 321 -1934 417 -1900
rect 1447 -1934 1543 -1900
rect 321 -1996 355 -1934
rect 1509 -1996 1543 -1934
rect 321 -2444 355 -2382
rect 1509 -2444 1543 -2382
rect 321 -2478 417 -2444
rect 1447 -2478 1543 -2444
rect 1842 -1934 1938 -1900
rect 2968 -1934 3064 -1900
rect 1842 -1996 1876 -1934
rect 3030 -1996 3064 -1934
rect 1842 -2444 1876 -2382
rect 3030 -2444 3064 -2382
rect 1842 -2478 1938 -2444
rect 2968 -2478 3064 -2444
<< psubdiffcont >>
rect -2254 -138 -1224 -104
rect -2350 -398 -2316 -200
rect -1162 -398 -1128 -200
rect -2254 -494 -1224 -460
rect 417 -138 1447 -104
rect 321 -398 355 -200
rect 1509 -398 1543 -200
rect 1938 -138 2968 -104
rect 1842 -398 1876 -200
rect 417 -494 1447 -460
rect 3030 -398 3064 -200
rect 1938 -494 2968 -460
rect -522 -797 -488 -763
rect 417 -1472 1447 -1438
rect -522 -1629 -488 -1595
rect 321 -1732 355 -1534
rect 1509 -1732 1543 -1534
rect 1938 -1472 2968 -1438
rect 1842 -1732 1876 -1534
rect 417 -1828 1447 -1794
rect 3030 -1732 3064 -1534
rect 1938 -1828 2968 -1794
rect -2254 -1934 -1224 -1900
rect -2350 -2194 -2316 -1996
rect -1162 -2194 -1128 -1996
rect -2254 -2290 -1224 -2256
<< nsubdiffcont >>
rect -2254 -600 -1224 -566
rect -2350 -1048 -2316 -662
rect -1162 -1048 -1128 -662
rect 417 -600 1447 -566
rect -2254 -1144 -1224 -1110
rect -522 -1015 -488 -981
rect -522 -1108 -488 -1074
rect 321 -1048 355 -662
rect 1509 -1048 1543 -662
rect 417 -1144 1447 -1110
rect 1938 -600 2968 -566
rect 1842 -1048 1876 -662
rect 3030 -1048 3064 -662
rect 1938 -1144 2968 -1110
rect -2254 -1284 -1224 -1250
rect -2350 -1732 -2316 -1346
rect -1162 -1732 -1128 -1346
rect -522 -1318 -488 -1284
rect -522 -1411 -488 -1377
rect -2254 -1828 -1224 -1794
rect 417 -1934 1447 -1900
rect 321 -2382 355 -1996
rect 1509 -2382 1543 -1996
rect 417 -2478 1447 -2444
rect 1938 -1934 2968 -1900
rect 1842 -2382 1876 -1996
rect 3030 -2382 3064 -1996
rect 1938 -2478 2968 -2444
<< poly >>
rect -2252 -197 -1226 -181
rect -2252 -231 -2236 -197
rect -2202 -231 -2044 -197
rect -2010 -231 -1852 -197
rect -1818 -231 -1660 -197
rect -1626 -231 -1468 -197
rect -1434 -231 -1276 -197
rect -1242 -231 -1226 -197
rect -2252 -247 -1226 -231
rect -2186 -278 -2156 -247
rect -2090 -278 -2060 -247
rect -1994 -278 -1964 -247
rect -1898 -278 -1868 -247
rect -1802 -278 -1772 -247
rect -1706 -278 -1676 -247
rect -1610 -278 -1580 -247
rect -1514 -278 -1484 -247
rect -1418 -278 -1388 -247
rect -1322 -278 -1292 -247
rect -2186 -408 -2156 -382
rect -2090 -408 -2060 -382
rect -1994 -408 -1964 -382
rect -1898 -408 -1868 -382
rect -1802 -408 -1772 -382
rect -1706 -408 -1676 -382
rect -1610 -408 -1580 -382
rect -1514 -408 -1484 -382
rect -1418 -408 -1388 -382
rect -1322 -408 -1292 -382
rect 419 -197 1445 -181
rect 419 -231 435 -197
rect 469 -231 627 -197
rect 661 -231 819 -197
rect 853 -231 1011 -197
rect 1045 -231 1203 -197
rect 1237 -231 1395 -197
rect 1429 -231 1445 -197
rect 419 -247 1445 -231
rect 485 -278 515 -247
rect 581 -278 611 -247
rect 677 -278 707 -247
rect 773 -278 803 -247
rect 869 -278 899 -247
rect 965 -278 995 -247
rect 1061 -278 1091 -247
rect 1157 -278 1187 -247
rect 1253 -278 1283 -247
rect 1349 -278 1379 -247
rect 485 -408 515 -382
rect 581 -408 611 -382
rect 677 -408 707 -382
rect 773 -408 803 -382
rect 869 -408 899 -382
rect 965 -408 995 -382
rect 1061 -408 1091 -382
rect 1157 -408 1187 -382
rect 1253 -408 1283 -382
rect 1349 -408 1379 -382
rect 1661 -284 1691 -258
rect 1661 -406 1691 -384
rect 1940 -197 2966 -181
rect 1940 -231 1956 -197
rect 1990 -231 2148 -197
rect 2182 -231 2340 -197
rect 2374 -231 2532 -197
rect 2566 -231 2724 -197
rect 2758 -231 2916 -197
rect 2950 -231 2966 -197
rect 1940 -247 2966 -231
rect 2006 -278 2036 -247
rect 2102 -278 2132 -247
rect 2198 -278 2228 -247
rect 2294 -278 2324 -247
rect 2390 -278 2420 -247
rect 2486 -278 2516 -247
rect 2582 -278 2612 -247
rect 2678 -278 2708 -247
rect 2774 -278 2804 -247
rect 2870 -278 2900 -247
rect 1643 -422 1709 -406
rect 1643 -456 1659 -422
rect 1693 -456 1709 -422
rect 1643 -472 1709 -456
rect 2006 -408 2036 -382
rect 2102 -408 2132 -382
rect 2198 -408 2228 -382
rect 2294 -408 2324 -382
rect 2390 -408 2420 -382
rect 2486 -408 2516 -382
rect 2582 -408 2612 -382
rect 2678 -408 2708 -382
rect 2774 -408 2804 -382
rect 2870 -408 2900 -382
rect -2186 -688 -2156 -662
rect -2090 -688 -2060 -662
rect -1994 -688 -1964 -662
rect -1898 -688 -1868 -662
rect -1802 -688 -1772 -662
rect -1706 -688 -1676 -662
rect -1610 -688 -1580 -662
rect -1514 -688 -1484 -662
rect -1418 -688 -1388 -662
rect -1322 -688 -1292 -662
rect -2186 -992 -2156 -960
rect -2090 -992 -2060 -960
rect -1994 -992 -1964 -960
rect -1898 -992 -1868 -960
rect -1802 -992 -1772 -960
rect -1706 -992 -1676 -960
rect -1610 -992 -1580 -960
rect -1514 -992 -1484 -960
rect -1418 -992 -1388 -960
rect -1322 -992 -1292 -960
rect -2252 -1008 -1226 -992
rect -2252 -1042 -2236 -1008
rect -2202 -1042 -2044 -1008
rect -2010 -1042 -1852 -1008
rect -1818 -1042 -1660 -1008
rect -1626 -1042 -1468 -1008
rect -1434 -1042 -1276 -1008
rect -1242 -1042 -1226 -1008
rect -2252 -1058 -1226 -1042
rect -339 -699 -309 -673
rect -339 -851 -309 -829
rect -395 -867 -309 -851
rect -395 -901 -379 -867
rect -345 -901 -309 -867
rect -395 -917 -309 -901
rect -339 -949 -309 -917
rect 485 -688 515 -662
rect 581 -688 611 -662
rect 677 -688 707 -662
rect 773 -688 803 -662
rect 869 -688 899 -662
rect 965 -688 995 -662
rect 1061 -688 1091 -662
rect 1157 -688 1187 -662
rect 1253 -688 1283 -662
rect 1349 -688 1379 -662
rect 485 -992 515 -960
rect 581 -992 611 -960
rect 677 -992 707 -960
rect 773 -992 803 -960
rect 869 -992 899 -960
rect 965 -992 995 -960
rect 1061 -992 1091 -960
rect 1157 -992 1187 -960
rect 1253 -992 1283 -960
rect 1349 -992 1379 -960
rect 419 -1008 1445 -992
rect 419 -1042 435 -1008
rect 469 -1042 627 -1008
rect 661 -1042 819 -1008
rect 853 -1042 1011 -1008
rect 1045 -1042 1203 -1008
rect 1237 -1042 1395 -1008
rect 1429 -1042 1445 -1008
rect 419 -1058 1445 -1042
rect 2006 -688 2036 -662
rect 2102 -688 2132 -662
rect 2198 -688 2228 -662
rect 2294 -688 2324 -662
rect 2390 -688 2420 -662
rect 2486 -688 2516 -662
rect 2582 -688 2612 -662
rect 2678 -688 2708 -662
rect 2774 -688 2804 -662
rect 2870 -688 2900 -662
rect 2006 -992 2036 -960
rect 2102 -992 2132 -960
rect 2198 -992 2228 -960
rect 2294 -992 2324 -960
rect 2390 -992 2420 -960
rect 2486 -992 2516 -960
rect 2582 -992 2612 -960
rect 2678 -992 2708 -960
rect 2774 -992 2804 -960
rect 2870 -992 2900 -960
rect 1940 -1008 2966 -992
rect 1940 -1042 1956 -1008
rect 1990 -1042 2148 -1008
rect 2182 -1042 2340 -1008
rect 2374 -1042 2532 -1008
rect 2566 -1042 2724 -1008
rect 2758 -1042 2916 -1008
rect 2950 -1042 2966 -1008
rect 1940 -1058 2966 -1042
rect -339 -1175 -309 -1149
rect -339 -1243 -309 -1217
rect -2252 -1352 -1226 -1336
rect -2252 -1386 -2236 -1352
rect -2202 -1386 -2044 -1352
rect -2010 -1386 -1852 -1352
rect -1818 -1386 -1660 -1352
rect -1626 -1386 -1468 -1352
rect -1434 -1386 -1276 -1352
rect -1242 -1386 -1226 -1352
rect -2252 -1402 -1226 -1386
rect -2186 -1434 -2156 -1402
rect -2090 -1434 -2060 -1402
rect -1994 -1434 -1964 -1402
rect -1898 -1434 -1868 -1402
rect -1802 -1434 -1772 -1402
rect -1706 -1434 -1676 -1402
rect -1610 -1434 -1580 -1402
rect -1514 -1434 -1484 -1402
rect -1418 -1434 -1388 -1402
rect -1322 -1434 -1292 -1402
rect -2186 -1732 -2156 -1706
rect -2090 -1732 -2060 -1706
rect -1994 -1732 -1964 -1706
rect -1898 -1732 -1868 -1706
rect -1802 -1732 -1772 -1706
rect -1706 -1732 -1676 -1706
rect -1610 -1732 -1580 -1706
rect -1514 -1732 -1484 -1706
rect -1418 -1732 -1388 -1706
rect -1322 -1732 -1292 -1706
rect -339 -1475 -309 -1443
rect -395 -1491 -309 -1475
rect -395 -1525 -379 -1491
rect -345 -1525 -309 -1491
rect -395 -1541 -309 -1525
rect -339 -1563 -309 -1541
rect -339 -1719 -309 -1693
rect 419 -1531 1445 -1515
rect 419 -1565 435 -1531
rect 469 -1565 627 -1531
rect 661 -1565 819 -1531
rect 853 -1565 1011 -1531
rect 1045 -1565 1203 -1531
rect 1237 -1565 1395 -1531
rect 1429 -1565 1445 -1531
rect 419 -1581 1445 -1565
rect 485 -1612 515 -1581
rect 581 -1612 611 -1581
rect 677 -1612 707 -1581
rect 773 -1612 803 -1581
rect 869 -1612 899 -1581
rect 965 -1612 995 -1581
rect 1061 -1612 1091 -1581
rect 1157 -1612 1187 -1581
rect 1253 -1612 1283 -1581
rect 1349 -1612 1379 -1581
rect 485 -1742 515 -1716
rect 581 -1742 611 -1716
rect 677 -1742 707 -1716
rect 773 -1742 803 -1716
rect 869 -1742 899 -1716
rect 965 -1742 995 -1716
rect 1061 -1742 1091 -1716
rect 1157 -1742 1187 -1716
rect 1253 -1742 1283 -1716
rect 1349 -1742 1379 -1716
rect 1661 -1618 1691 -1592
rect 1661 -1740 1691 -1718
rect 1940 -1531 2966 -1515
rect 1940 -1565 1956 -1531
rect 1990 -1565 2148 -1531
rect 2182 -1565 2340 -1531
rect 2374 -1565 2532 -1531
rect 2566 -1565 2724 -1531
rect 2758 -1565 2916 -1531
rect 2950 -1565 2966 -1531
rect 1940 -1581 2966 -1565
rect 2006 -1612 2036 -1581
rect 2102 -1612 2132 -1581
rect 2198 -1612 2228 -1581
rect 2294 -1612 2324 -1581
rect 2390 -1612 2420 -1581
rect 2486 -1612 2516 -1581
rect 2582 -1612 2612 -1581
rect 2678 -1612 2708 -1581
rect 2774 -1612 2804 -1581
rect 2870 -1612 2900 -1581
rect 1643 -1756 1709 -1740
rect 1643 -1790 1659 -1756
rect 1693 -1790 1709 -1756
rect 1643 -1806 1709 -1790
rect 2006 -1742 2036 -1716
rect 2102 -1742 2132 -1716
rect 2198 -1742 2228 -1716
rect 2294 -1742 2324 -1716
rect 2390 -1742 2420 -1716
rect 2486 -1742 2516 -1716
rect 2582 -1742 2612 -1716
rect 2678 -1742 2708 -1716
rect 2774 -1742 2804 -1716
rect 2870 -1742 2900 -1716
rect -2186 -2012 -2156 -1986
rect -2090 -2012 -2060 -1986
rect -1994 -2012 -1964 -1986
rect -1898 -2012 -1868 -1986
rect -1802 -2012 -1772 -1986
rect -1706 -2012 -1676 -1986
rect -1610 -2012 -1580 -1986
rect -1514 -2012 -1484 -1986
rect -1418 -2012 -1388 -1986
rect -1322 -2012 -1292 -1986
rect -2186 -2147 -2156 -2116
rect -2090 -2147 -2060 -2116
rect -1994 -2147 -1964 -2116
rect -1898 -2147 -1868 -2116
rect -1802 -2147 -1772 -2116
rect -1706 -2147 -1676 -2116
rect -1610 -2147 -1580 -2116
rect -1514 -2147 -1484 -2116
rect -1418 -2147 -1388 -2116
rect -1322 -2147 -1292 -2116
rect -2252 -2163 -1226 -2147
rect -2252 -2197 -2236 -2163
rect -2202 -2197 -2044 -2163
rect -2010 -2197 -1852 -2163
rect -1818 -2197 -1660 -2163
rect -1626 -2197 -1468 -2163
rect -1434 -2197 -1276 -2163
rect -1242 -2197 -1226 -2163
rect -2252 -2213 -1226 -2197
rect 485 -2022 515 -1996
rect 581 -2022 611 -1996
rect 677 -2022 707 -1996
rect 773 -2022 803 -1996
rect 869 -2022 899 -1996
rect 965 -2022 995 -1996
rect 1061 -2022 1091 -1996
rect 1157 -2022 1187 -1996
rect 1253 -2022 1283 -1996
rect 1349 -2022 1379 -1996
rect 485 -2326 515 -2294
rect 581 -2326 611 -2294
rect 677 -2326 707 -2294
rect 773 -2326 803 -2294
rect 869 -2326 899 -2294
rect 965 -2326 995 -2294
rect 1061 -2326 1091 -2294
rect 1157 -2326 1187 -2294
rect 1253 -2326 1283 -2294
rect 1349 -2326 1379 -2294
rect 419 -2342 1445 -2326
rect 419 -2376 435 -2342
rect 469 -2376 627 -2342
rect 661 -2376 819 -2342
rect 853 -2376 1011 -2342
rect 1045 -2376 1203 -2342
rect 1237 -2376 1395 -2342
rect 1429 -2376 1445 -2342
rect 419 -2392 1445 -2376
rect 2006 -2022 2036 -1996
rect 2102 -2022 2132 -1996
rect 2198 -2022 2228 -1996
rect 2294 -2022 2324 -1996
rect 2390 -2022 2420 -1996
rect 2486 -2022 2516 -1996
rect 2582 -2022 2612 -1996
rect 2678 -2022 2708 -1996
rect 2774 -2022 2804 -1996
rect 2870 -2022 2900 -1996
rect 2006 -2326 2036 -2294
rect 2102 -2326 2132 -2294
rect 2198 -2326 2228 -2294
rect 2294 -2326 2324 -2294
rect 2390 -2326 2420 -2294
rect 2486 -2326 2516 -2294
rect 2582 -2326 2612 -2294
rect 2678 -2326 2708 -2294
rect 2774 -2326 2804 -2294
rect 2870 -2326 2900 -2294
rect 1940 -2342 2966 -2326
rect 1940 -2376 1956 -2342
rect 1990 -2376 2148 -2342
rect 2182 -2376 2340 -2342
rect 2374 -2376 2532 -2342
rect 2566 -2376 2724 -2342
rect 2758 -2376 2916 -2342
rect 2950 -2376 2966 -2342
rect 1940 -2392 2966 -2376
<< polycont >>
rect -2236 -231 -2202 -197
rect -2044 -231 -2010 -197
rect -1852 -231 -1818 -197
rect -1660 -231 -1626 -197
rect -1468 -231 -1434 -197
rect -1276 -231 -1242 -197
rect 435 -231 469 -197
rect 627 -231 661 -197
rect 819 -231 853 -197
rect 1011 -231 1045 -197
rect 1203 -231 1237 -197
rect 1395 -231 1429 -197
rect 1956 -231 1990 -197
rect 2148 -231 2182 -197
rect 2340 -231 2374 -197
rect 2532 -231 2566 -197
rect 2724 -231 2758 -197
rect 2916 -231 2950 -197
rect 1659 -456 1693 -422
rect -2236 -1042 -2202 -1008
rect -2044 -1042 -2010 -1008
rect -1852 -1042 -1818 -1008
rect -1660 -1042 -1626 -1008
rect -1468 -1042 -1434 -1008
rect -1276 -1042 -1242 -1008
rect -379 -901 -345 -867
rect 435 -1042 469 -1008
rect 627 -1042 661 -1008
rect 819 -1042 853 -1008
rect 1011 -1042 1045 -1008
rect 1203 -1042 1237 -1008
rect 1395 -1042 1429 -1008
rect 1956 -1042 1990 -1008
rect 2148 -1042 2182 -1008
rect 2340 -1042 2374 -1008
rect 2532 -1042 2566 -1008
rect 2724 -1042 2758 -1008
rect 2916 -1042 2950 -1008
rect -2236 -1386 -2202 -1352
rect -2044 -1386 -2010 -1352
rect -1852 -1386 -1818 -1352
rect -1660 -1386 -1626 -1352
rect -1468 -1386 -1434 -1352
rect -1276 -1386 -1242 -1352
rect -379 -1525 -345 -1491
rect 435 -1565 469 -1531
rect 627 -1565 661 -1531
rect 819 -1565 853 -1531
rect 1011 -1565 1045 -1531
rect 1203 -1565 1237 -1531
rect 1395 -1565 1429 -1531
rect 1956 -1565 1990 -1531
rect 2148 -1565 2182 -1531
rect 2340 -1565 2374 -1531
rect 2532 -1565 2566 -1531
rect 2724 -1565 2758 -1531
rect 2916 -1565 2950 -1531
rect 1659 -1790 1693 -1756
rect -2236 -2197 -2202 -2163
rect -2044 -2197 -2010 -2163
rect -1852 -2197 -1818 -2163
rect -1660 -2197 -1626 -2163
rect -1468 -2197 -1434 -2163
rect -1276 -2197 -1242 -2163
rect 435 -2376 469 -2342
rect 627 -2376 661 -2342
rect 819 -2376 853 -2342
rect 1011 -2376 1045 -2342
rect 1203 -2376 1237 -2342
rect 1395 -2376 1429 -2342
rect 1956 -2376 1990 -2342
rect 2148 -2376 2182 -2342
rect 2340 -2376 2374 -2342
rect 2532 -2376 2566 -2342
rect 2724 -2376 2758 -2342
rect 2916 -2376 2950 -2342
<< locali >>
rect -2626 115 3466 243
rect -2350 -138 -2254 -104
rect -1224 -138 -1128 -104
rect -2350 -200 -2316 -138
rect -2252 -197 -1226 -189
rect -2252 -231 -2236 -197
rect -2202 -231 -2044 -197
rect -2010 -231 -1852 -197
rect -1818 -231 -1660 -197
rect -1626 -231 -1468 -197
rect -1434 -231 -1276 -197
rect -1242 -231 -1226 -197
rect -2252 -239 -1226 -231
rect -1162 -200 -1128 -138
rect -2236 -290 -2202 -274
rect -2236 -386 -2202 -370
rect -2140 -290 -2106 -274
rect -2140 -386 -2106 -370
rect -2044 -290 -2010 -274
rect -2044 -386 -2010 -370
rect -1948 -290 -1914 -274
rect -1948 -386 -1914 -370
rect -1852 -290 -1818 -274
rect -1852 -386 -1818 -370
rect -1756 -290 -1722 -274
rect -1756 -386 -1722 -370
rect -1660 -290 -1626 -274
rect -1660 -386 -1626 -370
rect -1564 -290 -1530 -274
rect -1564 -386 -1530 -370
rect -1468 -290 -1434 -274
rect -1468 -386 -1434 -370
rect -1372 -290 -1338 -274
rect -1372 -386 -1338 -370
rect -1276 -290 -1242 -274
rect -1276 -386 -1242 -370
rect -2350 -429 -2316 -398
rect -2599 -460 -2316 -429
rect -1162 -460 -1128 -398
rect -2599 -493 -2254 -460
rect -2599 -2678 -2535 -493
rect -2350 -494 -2254 -493
rect -1224 -494 -1128 -460
rect -2350 -600 -2254 -566
rect -1224 -600 -1128 -566
rect -2350 -662 -2316 -600
rect -1162 -662 -1128 -600
rect -2236 -700 -2202 -684
rect -2236 -964 -2202 -948
rect -2140 -700 -2106 -684
rect -2140 -964 -2106 -948
rect -2044 -700 -2010 -684
rect -2044 -964 -2010 -948
rect -1948 -700 -1914 -684
rect -1948 -964 -1914 -948
rect -1852 -700 -1818 -684
rect -1852 -964 -1818 -948
rect -1756 -700 -1722 -684
rect -1756 -964 -1722 -948
rect -1660 -700 -1626 -684
rect -1660 -964 -1626 -948
rect -1564 -700 -1530 -684
rect -1564 -964 -1530 -948
rect -1468 -700 -1434 -684
rect -1468 -964 -1434 -948
rect -1372 -700 -1338 -684
rect -1372 -964 -1338 -948
rect -1276 -700 -1242 -684
rect -1276 -964 -1242 -948
rect -2350 -1110 -2316 -1048
rect -2252 -1008 -1226 -1000
rect -2252 -1042 -2236 -1008
rect -2202 -1042 -2044 -1008
rect -2010 -1042 -1852 -1008
rect -1818 -1042 -1660 -1008
rect -1626 -1042 -1468 -1008
rect -1434 -1042 -1276 -1008
rect -1242 -1042 -1226 -1008
rect -2252 -1050 -1226 -1042
rect -1162 -1110 -1128 -1048
rect -2350 -1144 -2254 -1110
rect -1224 -1123 -1128 -1110
rect -1224 -1144 -1122 -1123
rect -1186 -1162 -1122 -1144
rect -870 -1162 -806 115
rect -626 -635 -510 -620
rect -626 -669 -522 -635
rect -488 -669 -430 -635
rect -396 -669 -338 -635
rect -304 -669 -246 -635
rect -212 -669 -183 -635
rect -626 -684 -476 -669
rect -534 -763 -476 -684
rect -534 -797 -522 -763
rect -488 -797 -476 -763
rect -534 -814 -476 -797
rect -395 -715 -349 -669
rect -395 -749 -383 -715
rect -395 -783 -349 -749
rect -395 -817 -383 -783
rect -395 -833 -349 -817
rect -315 -715 -249 -703
rect -315 -749 -299 -715
rect -265 -749 -249 -715
rect -315 -778 -249 -749
rect -315 -783 -298 -778
rect -315 -817 -299 -783
rect -264 -812 -249 -778
rect -265 -817 -249 -812
rect -315 -829 -249 -817
rect -395 -873 -379 -867
rect -395 -907 -381 -873
rect -345 -901 -329 -867
rect -347 -907 -329 -901
rect -395 -915 -329 -907
rect -534 -981 -476 -946
rect -295 -949 -249 -829
rect -534 -1015 -522 -981
rect -488 -1015 -476 -981
rect -534 -1074 -476 -1015
rect -534 -1108 -522 -1074
rect -488 -1108 -476 -1074
rect -534 -1162 -476 -1108
rect -391 -967 -349 -951
rect -391 -1001 -383 -967
rect -391 -1035 -349 -1001
rect -391 -1069 -383 -1035
rect -391 -1103 -349 -1069
rect -391 -1137 -383 -1103
rect -391 -1162 -349 -1137
rect -315 -967 -249 -949
rect -315 -1001 -299 -967
rect -265 -1001 -249 -967
rect -315 -1035 -249 -1001
rect -315 -1069 -299 -1035
rect -265 -1069 -249 -1035
rect -315 -1103 -249 -1069
rect -315 -1137 -299 -1103
rect -265 -1137 -249 -1103
rect -315 -1145 -249 -1137
rect -74 -1077 -10 115
rect 1637 -51 3236 13
rect 1637 -102 1701 -51
rect 3172 -102 3236 -51
rect 1491 -104 1889 -102
rect 3038 -104 3236 -102
rect 321 -138 417 -104
rect 1447 -138 1938 -104
rect 2968 -138 3236 -104
rect 321 -200 355 -138
rect 1509 -170 1876 -138
rect 419 -197 1445 -189
rect 419 -231 435 -197
rect 469 -231 627 -197
rect 661 -231 819 -197
rect 853 -231 1011 -197
rect 1045 -231 1203 -197
rect 1237 -231 1395 -197
rect 1429 -231 1445 -197
rect 419 -239 1445 -231
rect 1509 -200 1543 -170
rect 435 -290 469 -274
rect 435 -386 469 -370
rect 531 -290 565 -274
rect 531 -386 565 -370
rect 627 -290 661 -274
rect 627 -386 661 -370
rect 723 -290 757 -274
rect 723 -386 757 -370
rect 819 -290 853 -274
rect 819 -386 853 -370
rect 915 -290 949 -274
rect 915 -386 949 -370
rect 1011 -290 1045 -274
rect 1011 -386 1045 -370
rect 1107 -290 1141 -274
rect 1107 -386 1141 -370
rect 1203 -290 1237 -274
rect 1203 -386 1237 -370
rect 1299 -290 1333 -274
rect 1299 -386 1333 -370
rect 1395 -290 1429 -274
rect 1395 -386 1429 -370
rect 1842 -200 1876 -170
rect 3030 -166 3236 -138
rect 321 -460 355 -398
rect 1615 -296 1649 -280
rect 1615 -388 1649 -372
rect 1703 -296 1737 -280
rect 1703 -388 1737 -372
rect 1509 -460 1543 -398
rect 1940 -197 2966 -189
rect 1940 -231 1956 -197
rect 1990 -231 2148 -197
rect 2182 -231 2340 -197
rect 2374 -231 2532 -197
rect 2566 -231 2724 -197
rect 2758 -231 2916 -197
rect 2950 -231 2966 -197
rect 1940 -239 2966 -231
rect 3030 -200 3064 -166
rect 1956 -290 1990 -274
rect 1956 -386 1990 -370
rect 2052 -290 2086 -274
rect 2052 -386 2086 -370
rect 2148 -290 2182 -274
rect 2148 -386 2182 -370
rect 2244 -290 2278 -274
rect 2244 -386 2278 -370
rect 2340 -290 2374 -274
rect 2340 -386 2374 -370
rect 2436 -290 2470 -274
rect 2436 -386 2470 -370
rect 2532 -290 2566 -274
rect 2532 -386 2566 -370
rect 2628 -290 2662 -274
rect 2628 -386 2662 -370
rect 2724 -290 2758 -274
rect 2724 -386 2758 -370
rect 2820 -290 2854 -274
rect 2820 -386 2854 -370
rect 2916 -290 2950 -274
rect 2916 -386 2950 -370
rect 1643 -456 1659 -422
rect 1693 -456 1709 -422
rect 321 -494 417 -460
rect 1447 -494 1543 -460
rect 1842 -460 1876 -398
rect 3030 -460 3064 -398
rect 1842 -494 1938 -460
rect 2968 -494 3064 -460
rect 321 -600 417 -566
rect 1447 -600 1543 -566
rect 321 -662 355 -600
rect 1509 -662 1543 -600
rect 435 -700 469 -684
rect 435 -964 469 -948
rect 531 -700 565 -684
rect 531 -964 565 -948
rect 627 -700 661 -684
rect 627 -964 661 -948
rect 723 -700 757 -684
rect 723 -964 757 -948
rect 819 -700 853 -684
rect 819 -964 853 -948
rect 915 -700 949 -684
rect 915 -964 949 -948
rect 1011 -700 1045 -684
rect 1011 -964 1045 -948
rect 1107 -700 1141 -684
rect 1107 -964 1141 -948
rect 1203 -700 1237 -684
rect 1203 -964 1237 -948
rect 1299 -700 1333 -684
rect 1299 -964 1333 -948
rect 1395 -700 1429 -684
rect 1395 -964 1429 -948
rect 321 -1077 355 -1048
rect 419 -1008 1445 -1000
rect 419 -1042 435 -1008
rect 469 -1042 627 -1008
rect 661 -1042 819 -1008
rect 853 -1042 1011 -1008
rect 1045 -1042 1203 -1008
rect 1237 -1042 1395 -1008
rect 1429 -1042 1445 -1008
rect 419 -1050 1445 -1042
rect -74 -1110 355 -1077
rect 1509 -1076 1543 -1048
rect 1842 -600 1938 -566
rect 2968 -600 3064 -566
rect 1842 -662 1876 -600
rect 3030 -662 3064 -600
rect 1956 -700 1990 -684
rect 1956 -964 1990 -948
rect 2052 -700 2086 -684
rect 2052 -964 2086 -948
rect 2148 -700 2182 -684
rect 2148 -964 2182 -948
rect 2244 -700 2278 -684
rect 2244 -964 2278 -948
rect 2340 -700 2374 -684
rect 2340 -964 2374 -948
rect 2436 -700 2470 -684
rect 2436 -964 2470 -948
rect 2532 -700 2566 -684
rect 2532 -964 2566 -948
rect 2628 -700 2662 -684
rect 2628 -964 2662 -948
rect 2724 -700 2758 -684
rect 2724 -964 2758 -948
rect 2820 -700 2854 -684
rect 2820 -964 2854 -948
rect 2916 -700 2950 -684
rect 2916 -964 2950 -948
rect 1647 -1076 1711 -1074
rect 1842 -1076 1876 -1048
rect 1940 -1008 2966 -1000
rect 1940 -1042 1956 -1008
rect 1990 -1042 2148 -1008
rect 2182 -1042 2340 -1008
rect 2374 -1042 2532 -1008
rect 2566 -1042 2724 -1008
rect 2758 -1042 2916 -1008
rect 2950 -1042 2966 -1008
rect 1940 -1050 2966 -1042
rect 1509 -1110 1882 -1076
rect 3030 -1110 3064 -1048
rect -74 -1141 417 -1110
rect -1186 -1179 -349 -1162
rect -1186 -1213 -522 -1179
rect -488 -1213 -430 -1179
rect -396 -1213 -338 -1179
rect -304 -1213 -246 -1179
rect -212 -1213 -183 -1179
rect -74 -1195 -10 -1141
rect 321 -1144 417 -1141
rect 1447 -1144 1938 -1110
rect 2968 -1144 3064 -1110
rect 1647 -1195 1711 -1144
rect -1186 -1226 -349 -1213
rect -1186 -1250 -1122 -1226
rect -2350 -1284 -2254 -1250
rect -1224 -1269 -1122 -1250
rect -1224 -1284 -1128 -1269
rect -2350 -1346 -2316 -1284
rect -2252 -1352 -1226 -1344
rect -2252 -1386 -2236 -1352
rect -2202 -1386 -2044 -1352
rect -2010 -1386 -1852 -1352
rect -1818 -1386 -1660 -1352
rect -1626 -1386 -1468 -1352
rect -1434 -1386 -1276 -1352
rect -1242 -1386 -1226 -1352
rect -2252 -1394 -1226 -1386
rect -1162 -1346 -1128 -1284
rect -2236 -1446 -2202 -1430
rect -2236 -1710 -2202 -1694
rect -2140 -1446 -2106 -1430
rect -2140 -1710 -2106 -1694
rect -2044 -1446 -2010 -1430
rect -2044 -1710 -2010 -1694
rect -1948 -1446 -1914 -1430
rect -1948 -1710 -1914 -1694
rect -1852 -1446 -1818 -1430
rect -1852 -1710 -1818 -1694
rect -1756 -1446 -1722 -1430
rect -1756 -1710 -1722 -1694
rect -1660 -1446 -1626 -1430
rect -1660 -1710 -1626 -1694
rect -1564 -1446 -1530 -1430
rect -1564 -1710 -1530 -1694
rect -1468 -1446 -1434 -1430
rect -1468 -1710 -1434 -1694
rect -1372 -1446 -1338 -1430
rect -1372 -1710 -1338 -1694
rect -1276 -1446 -1242 -1430
rect -1276 -1710 -1242 -1694
rect -2350 -1794 -2316 -1732
rect -534 -1284 -476 -1226
rect -534 -1318 -522 -1284
rect -488 -1318 -476 -1284
rect -534 -1377 -476 -1318
rect -534 -1411 -522 -1377
rect -488 -1411 -476 -1377
rect -534 -1446 -476 -1411
rect -391 -1255 -349 -1226
rect -391 -1289 -383 -1255
rect -391 -1323 -349 -1289
rect -391 -1357 -383 -1323
rect -391 -1391 -349 -1357
rect -391 -1425 -383 -1391
rect -391 -1441 -349 -1425
rect -315 -1255 -249 -1247
rect -315 -1289 -299 -1255
rect -265 -1289 -249 -1255
rect -315 -1323 -249 -1289
rect -315 -1382 -299 -1323
rect -265 -1382 -249 -1323
rect -315 -1391 -249 -1382
rect -315 -1425 -299 -1391
rect -265 -1425 -249 -1391
rect -315 -1443 -249 -1425
rect -395 -1486 -329 -1477
rect -395 -1520 -382 -1486
rect -348 -1491 -329 -1486
rect -395 -1525 -379 -1520
rect -345 -1525 -329 -1491
rect -395 -1575 -349 -1559
rect -295 -1563 -249 -1443
rect -534 -1595 -476 -1578
rect -534 -1629 -522 -1595
rect -488 -1629 -476 -1595
rect -534 -1710 -476 -1629
rect -1162 -1794 -1128 -1732
rect -697 -1718 -476 -1710
rect -697 -1779 -690 -1718
rect -626 -1723 -476 -1718
rect -395 -1609 -383 -1575
rect -395 -1643 -349 -1609
rect -395 -1677 -383 -1643
rect -395 -1723 -349 -1677
rect -315 -1575 -249 -1563
rect -315 -1609 -299 -1575
rect -265 -1609 -249 -1575
rect -315 -1643 -249 -1609
rect -315 -1677 -299 -1643
rect -265 -1677 -249 -1643
rect -315 -1689 -249 -1677
rect -74 -1259 1711 -1195
rect -626 -1757 -522 -1723
rect -488 -1757 -430 -1723
rect -396 -1757 -338 -1723
rect -304 -1757 -246 -1723
rect -212 -1757 -183 -1723
rect -626 -1779 -501 -1757
rect -626 -1782 -625 -1779
rect -2350 -1828 -2254 -1794
rect -1224 -1828 -1128 -1794
rect -2350 -1934 -2254 -1900
rect -1224 -1934 -1128 -1900
rect -2350 -1996 -2316 -1934
rect -1162 -1996 -1128 -1934
rect -2236 -2024 -2202 -2008
rect -2236 -2120 -2202 -2104
rect -2140 -2024 -2106 -2008
rect -2140 -2120 -2106 -2104
rect -2044 -2024 -2010 -2008
rect -2044 -2120 -2010 -2104
rect -1948 -2024 -1914 -2008
rect -1948 -2120 -1914 -2104
rect -1852 -2024 -1818 -2008
rect -1852 -2120 -1818 -2104
rect -1756 -2024 -1722 -2008
rect -1756 -2120 -1722 -2104
rect -1660 -2024 -1626 -2008
rect -1660 -2120 -1626 -2104
rect -1564 -2024 -1530 -2008
rect -1564 -2120 -1530 -2104
rect -1468 -2024 -1434 -2008
rect -1468 -2120 -1434 -2104
rect -1372 -2024 -1338 -2008
rect -1372 -2120 -1338 -2104
rect -1276 -2024 -1242 -2008
rect -1276 -2120 -1242 -2104
rect -2350 -2256 -2316 -2194
rect -2252 -2163 -1226 -2155
rect -2252 -2197 -2236 -2163
rect -2202 -2197 -2044 -2163
rect -2010 -2197 -1852 -2163
rect -1818 -2197 -1660 -2163
rect -1626 -2197 -1468 -2163
rect -1434 -2197 -1276 -2163
rect -1242 -2197 -1226 -2163
rect -2252 -2205 -1226 -2197
rect -1162 -2256 -1128 -2194
rect -2350 -2290 -2254 -2256
rect -1224 -2290 -1128 -2256
rect -1204 -2678 -1140 -2290
rect -689 -2678 -625 -1782
rect -74 -2410 -10 -1259
rect 3172 -1336 3236 -166
rect 1645 -1400 3236 -1336
rect 1645 -1436 1709 -1400
rect 1491 -1438 1889 -1436
rect 321 -1472 417 -1438
rect 1447 -1472 1938 -1438
rect 2968 -1442 3064 -1438
rect 3172 -1442 3236 -1400
rect 2968 -1472 3236 -1442
rect 321 -1534 355 -1472
rect 1509 -1504 1876 -1472
rect 419 -1531 1445 -1523
rect 419 -1565 435 -1531
rect 469 -1565 627 -1531
rect 661 -1565 819 -1531
rect 853 -1565 1011 -1531
rect 1045 -1565 1203 -1531
rect 1237 -1565 1395 -1531
rect 1429 -1565 1445 -1531
rect 419 -1573 1445 -1565
rect 1509 -1534 1543 -1504
rect 435 -1624 469 -1608
rect 435 -1720 469 -1704
rect 531 -1624 565 -1608
rect 531 -1720 565 -1704
rect 627 -1624 661 -1608
rect 627 -1720 661 -1704
rect 723 -1624 757 -1608
rect 723 -1720 757 -1704
rect 819 -1624 853 -1608
rect 819 -1720 853 -1704
rect 915 -1624 949 -1608
rect 915 -1720 949 -1704
rect 1011 -1624 1045 -1608
rect 1011 -1720 1045 -1704
rect 1107 -1624 1141 -1608
rect 1107 -1720 1141 -1704
rect 1203 -1624 1237 -1608
rect 1203 -1720 1237 -1704
rect 1299 -1624 1333 -1608
rect 1299 -1720 1333 -1704
rect 1395 -1624 1429 -1608
rect 1395 -1720 1429 -1704
rect 1842 -1534 1876 -1504
rect 3030 -1506 3236 -1472
rect 321 -1794 355 -1732
rect 1615 -1630 1649 -1614
rect 1615 -1722 1649 -1706
rect 1703 -1630 1737 -1614
rect 1703 -1722 1737 -1706
rect 1509 -1794 1543 -1732
rect 1940 -1531 2966 -1523
rect 1940 -1565 1956 -1531
rect 1990 -1565 2148 -1531
rect 2182 -1565 2340 -1531
rect 2374 -1565 2532 -1531
rect 2566 -1565 2724 -1531
rect 2758 -1565 2916 -1531
rect 2950 -1565 2966 -1531
rect 1940 -1573 2966 -1565
rect 3030 -1534 3064 -1506
rect 1956 -1624 1990 -1608
rect 1956 -1720 1990 -1704
rect 2052 -1624 2086 -1608
rect 2052 -1720 2086 -1704
rect 2148 -1624 2182 -1608
rect 2148 -1720 2182 -1704
rect 2244 -1624 2278 -1608
rect 2244 -1720 2278 -1704
rect 2340 -1624 2374 -1608
rect 2340 -1720 2374 -1704
rect 2436 -1624 2470 -1608
rect 2436 -1720 2470 -1704
rect 2532 -1624 2566 -1608
rect 2532 -1720 2566 -1704
rect 2628 -1624 2662 -1608
rect 2628 -1720 2662 -1704
rect 2724 -1624 2758 -1608
rect 2724 -1720 2758 -1704
rect 2820 -1624 2854 -1608
rect 2820 -1720 2854 -1704
rect 2916 -1624 2950 -1608
rect 2916 -1720 2950 -1704
rect 1643 -1790 1659 -1756
rect 1693 -1790 1709 -1756
rect 321 -1828 417 -1794
rect 1447 -1828 1543 -1794
rect 1842 -1794 1876 -1732
rect 3030 -1794 3064 -1732
rect 1842 -1828 1938 -1794
rect 2968 -1828 3064 -1794
rect 321 -1934 417 -1900
rect 1447 -1934 1543 -1900
rect 321 -1996 355 -1934
rect 1509 -1996 1543 -1934
rect 435 -2034 469 -2018
rect 435 -2298 469 -2282
rect 531 -2034 565 -2018
rect 531 -2298 565 -2282
rect 627 -2034 661 -2018
rect 627 -2298 661 -2282
rect 723 -2034 757 -2018
rect 723 -2298 757 -2282
rect 819 -2034 853 -2018
rect 819 -2298 853 -2282
rect 915 -2034 949 -2018
rect 915 -2298 949 -2282
rect 1011 -2034 1045 -2018
rect 1011 -2298 1045 -2282
rect 1107 -2034 1141 -2018
rect 1107 -2298 1141 -2282
rect 1203 -2034 1237 -2018
rect 1203 -2298 1237 -2282
rect 1299 -2034 1333 -2018
rect 1299 -2298 1333 -2282
rect 1395 -2034 1429 -2018
rect 1395 -2298 1429 -2282
rect 321 -2410 355 -2382
rect 419 -2342 1445 -2334
rect 419 -2376 435 -2342
rect 469 -2376 627 -2342
rect 661 -2376 819 -2342
rect 853 -2376 1011 -2342
rect 1045 -2376 1203 -2342
rect 1237 -2376 1395 -2342
rect 1429 -2376 1445 -2342
rect 419 -2384 1445 -2376
rect -74 -2444 355 -2410
rect 1509 -2410 1543 -2382
rect 1842 -1934 1938 -1900
rect 2968 -1934 3064 -1900
rect 1842 -1996 1876 -1934
rect 3030 -1996 3064 -1934
rect 1956 -2034 1990 -2018
rect 1956 -2298 1990 -2282
rect 2052 -2034 2086 -2018
rect 2052 -2298 2086 -2282
rect 2148 -2034 2182 -2018
rect 2148 -2298 2182 -2282
rect 2244 -2034 2278 -2018
rect 2244 -2298 2278 -2282
rect 2340 -2034 2374 -2018
rect 2340 -2298 2374 -2282
rect 2436 -2034 2470 -2018
rect 2436 -2298 2470 -2282
rect 2532 -2034 2566 -2018
rect 2532 -2298 2566 -2282
rect 2628 -2034 2662 -2018
rect 2628 -2298 2662 -2282
rect 2724 -2034 2758 -2018
rect 2724 -2298 2758 -2282
rect 2820 -2034 2854 -2018
rect 2820 -2298 2854 -2282
rect 2916 -2034 2950 -2018
rect 2916 -2298 2950 -2282
rect 1842 -2410 1876 -2382
rect 1940 -2342 2966 -2334
rect 1940 -2376 1956 -2342
rect 1990 -2376 2148 -2342
rect 2182 -2376 2340 -2342
rect 2374 -2376 2532 -2342
rect 2566 -2376 2724 -2342
rect 2758 -2376 2916 -2342
rect 2950 -2376 2966 -2342
rect 1940 -2384 2966 -2376
rect 1509 -2444 1882 -2410
rect 3030 -2444 3064 -2382
rect -74 -2474 417 -2444
rect -74 -2529 -10 -2474
rect 321 -2478 417 -2474
rect 1447 -2478 1938 -2444
rect 2968 -2478 3064 -2444
rect 1643 -2529 1707 -2478
rect -74 -2593 1707 -2529
rect 3172 -2678 3236 -1506
rect -2626 -2806 3466 -2678
<< viali >>
rect -1276 -231 -1242 -197
rect -2236 -370 -2202 -290
rect -2140 -370 -2106 -290
rect -2044 -370 -2010 -290
rect -1948 -370 -1914 -290
rect -1852 -370 -1818 -290
rect -1756 -370 -1722 -290
rect -1660 -370 -1626 -290
rect -1564 -370 -1530 -290
rect -1468 -370 -1434 -290
rect -1372 -370 -1338 -290
rect -1276 -370 -1242 -290
rect -2236 -948 -2202 -700
rect -2140 -948 -2106 -700
rect -2044 -948 -2010 -700
rect -1948 -948 -1914 -700
rect -1852 -948 -1818 -700
rect -1756 -948 -1722 -700
rect -1660 -948 -1626 -700
rect -1564 -948 -1530 -700
rect -1468 -948 -1434 -700
rect -1372 -948 -1338 -700
rect -1276 -948 -1242 -700
rect -1276 -1042 -1242 -1008
rect -690 -684 -626 -620
rect -522 -669 -488 -635
rect -430 -669 -396 -635
rect -338 -669 -304 -635
rect -246 -669 -212 -635
rect -298 -783 -264 -778
rect -298 -812 -265 -783
rect -265 -812 -264 -783
rect -381 -901 -379 -873
rect -379 -901 -347 -873
rect -381 -907 -347 -901
rect 435 -231 469 -197
rect 1395 -231 1429 -197
rect 435 -370 469 -290
rect 531 -370 565 -290
rect 627 -370 661 -290
rect 723 -370 757 -290
rect 819 -370 853 -290
rect 915 -370 949 -290
rect 1011 -370 1045 -290
rect 1107 -370 1141 -290
rect 1203 -370 1237 -290
rect 1299 -370 1333 -290
rect 1395 -370 1429 -290
rect 1509 -385 1543 -285
rect 1615 -372 1649 -296
rect 1703 -372 1737 -296
rect 1956 -231 1990 -197
rect 2916 -231 2950 -197
rect 1956 -370 1990 -290
rect 2052 -370 2086 -290
rect 2148 -370 2182 -290
rect 2244 -370 2278 -290
rect 2340 -370 2374 -290
rect 2436 -370 2470 -290
rect 2532 -370 2566 -290
rect 2628 -370 2662 -290
rect 2724 -370 2758 -290
rect 2820 -370 2854 -290
rect 2916 -370 2950 -290
rect 1659 -456 1693 -422
rect 435 -948 469 -700
rect 531 -948 565 -700
rect 627 -948 661 -700
rect 723 -948 757 -700
rect 819 -948 853 -700
rect 915 -948 949 -700
rect 1011 -948 1045 -700
rect 1107 -948 1141 -700
rect 1203 -948 1237 -700
rect 1299 -948 1333 -700
rect 1395 -948 1429 -700
rect 435 -1042 469 -1008
rect 1395 -1042 1429 -1008
rect 1956 -948 1990 -700
rect 2052 -948 2086 -700
rect 2148 -948 2182 -700
rect 2244 -948 2278 -700
rect 2340 -948 2374 -700
rect 2436 -948 2470 -700
rect 2532 -948 2566 -700
rect 2628 -948 2662 -700
rect 2724 -948 2758 -700
rect 2820 -948 2854 -700
rect 2916 -948 2950 -700
rect 1956 -1042 1990 -1008
rect 2916 -1042 2950 -1008
rect -522 -1213 -488 -1179
rect -430 -1213 -396 -1179
rect -338 -1213 -304 -1179
rect -246 -1213 -212 -1179
rect -1276 -1386 -1242 -1352
rect -2236 -1694 -2202 -1446
rect -2140 -1694 -2106 -1446
rect -2044 -1694 -2010 -1446
rect -1948 -1694 -1914 -1446
rect -1852 -1694 -1818 -1446
rect -1756 -1694 -1722 -1446
rect -1660 -1694 -1626 -1446
rect -1564 -1694 -1530 -1446
rect -1468 -1694 -1434 -1446
rect -1372 -1694 -1338 -1446
rect -1276 -1694 -1242 -1446
rect -299 -1357 -265 -1348
rect -299 -1382 -265 -1357
rect -382 -1491 -348 -1486
rect -382 -1520 -379 -1491
rect -379 -1520 -348 -1491
rect -690 -1782 -626 -1718
rect -522 -1757 -488 -1723
rect -430 -1757 -396 -1723
rect -338 -1757 -304 -1723
rect -246 -1757 -212 -1723
rect -2236 -2104 -2202 -2024
rect -2140 -2104 -2106 -2024
rect -2044 -2104 -2010 -2024
rect -1948 -2104 -1914 -2024
rect -1852 -2104 -1818 -2024
rect -1756 -2104 -1722 -2024
rect -1660 -2104 -1626 -2024
rect -1564 -2104 -1530 -2024
rect -1468 -2104 -1434 -2024
rect -1372 -2104 -1338 -2024
rect -1276 -2104 -1242 -2024
rect -1276 -2197 -1242 -2163
rect 435 -1565 469 -1531
rect 1395 -1565 1429 -1531
rect 435 -1704 469 -1624
rect 531 -1704 565 -1624
rect 627 -1704 661 -1624
rect 723 -1704 757 -1624
rect 819 -1704 853 -1624
rect 915 -1704 949 -1624
rect 1011 -1704 1045 -1624
rect 1107 -1704 1141 -1624
rect 1203 -1704 1237 -1624
rect 1299 -1704 1333 -1624
rect 1395 -1704 1429 -1624
rect 1509 -1719 1543 -1619
rect 1615 -1706 1649 -1630
rect 1703 -1706 1737 -1630
rect 1956 -1565 1990 -1531
rect 2916 -1565 2950 -1531
rect 1956 -1704 1990 -1624
rect 2052 -1704 2086 -1624
rect 2148 -1704 2182 -1624
rect 2244 -1704 2278 -1624
rect 2340 -1704 2374 -1624
rect 2436 -1704 2470 -1624
rect 2532 -1704 2566 -1624
rect 2628 -1704 2662 -1624
rect 2724 -1704 2758 -1624
rect 2820 -1704 2854 -1624
rect 2916 -1704 2950 -1624
rect 1659 -1790 1693 -1756
rect 435 -2282 469 -2034
rect 531 -2282 565 -2034
rect 627 -2282 661 -2034
rect 723 -2282 757 -2034
rect 819 -2282 853 -2034
rect 915 -2282 949 -2034
rect 1011 -2282 1045 -2034
rect 1107 -2282 1141 -2034
rect 1203 -2282 1237 -2034
rect 1299 -2282 1333 -2034
rect 1395 -2282 1429 -2034
rect 435 -2376 469 -2342
rect 1395 -2376 1429 -2342
rect 1956 -2282 1990 -2034
rect 2052 -2282 2086 -2034
rect 2148 -2282 2182 -2034
rect 2244 -2282 2278 -2034
rect 2340 -2282 2374 -2034
rect 2436 -2282 2470 -2034
rect 2532 -2282 2566 -2034
rect 2628 -2282 2662 -2034
rect 2724 -2282 2758 -2034
rect 2820 -2282 2854 -2034
rect 2916 -2282 2950 -2034
rect 1956 -2376 1990 -2342
rect 2916 -2376 2950 -2342
<< metal1 >>
rect -2386 -136 -1338 -102
rect -2386 -513 -2352 -136
rect -2140 -278 -2106 -136
rect -1948 -278 -1914 -136
rect -1756 -278 -1722 -136
rect -1564 -278 -1530 -136
rect -1372 -278 -1338 -136
rect 285 -136 1333 -102
rect -1297 -240 -1287 -188
rect -1235 -240 -1225 -188
rect -2242 -290 -2196 -278
rect -2242 -370 -2236 -290
rect -2202 -370 -2196 -290
rect -2242 -382 -2196 -370
rect -2146 -290 -2100 -278
rect -2146 -370 -2140 -290
rect -2106 -370 -2100 -290
rect -2146 -382 -2100 -370
rect -2050 -290 -2004 -278
rect -2050 -370 -2044 -290
rect -2010 -370 -2004 -290
rect -2050 -382 -2004 -370
rect -1954 -290 -1908 -278
rect -1954 -370 -1948 -290
rect -1914 -370 -1908 -290
rect -1954 -382 -1908 -370
rect -1858 -290 -1812 -278
rect -1858 -370 -1852 -290
rect -1818 -370 -1812 -290
rect -1858 -382 -1812 -370
rect -1762 -290 -1716 -278
rect -1762 -370 -1756 -290
rect -1722 -370 -1716 -290
rect -1762 -382 -1716 -370
rect -1666 -290 -1620 -278
rect -1666 -370 -1660 -290
rect -1626 -370 -1620 -290
rect -1666 -382 -1620 -370
rect -1570 -290 -1524 -278
rect -1570 -370 -1564 -290
rect -1530 -370 -1524 -290
rect -1570 -382 -1524 -370
rect -1474 -290 -1428 -278
rect -1474 -370 -1468 -290
rect -1434 -370 -1428 -290
rect -1474 -382 -1428 -370
rect -1378 -290 -1332 -278
rect -1378 -370 -1372 -290
rect -1338 -370 -1332 -290
rect -1378 -382 -1332 -370
rect -1282 -290 -1236 -278
rect -1282 -370 -1276 -290
rect -1242 -370 -1236 -290
rect -1282 -382 -1236 -370
rect -2638 -547 -2352 -513
rect -2386 -1110 -2352 -547
rect -2236 -513 -2202 -382
rect -2044 -513 -2010 -382
rect -1852 -513 -1818 -382
rect -1660 -513 -1626 -382
rect -1468 -513 -1434 -382
rect -1276 -513 -1242 -382
rect -1046 -479 104 -445
rect -1046 -513 -1012 -479
rect -2236 -547 -1012 -513
rect 70 -503 104 -479
rect 285 -503 319 -136
rect 415 -238 425 -186
rect 477 -238 487 -186
rect 531 -278 565 -136
rect 723 -278 757 -136
rect 915 -278 949 -136
rect 1107 -278 1141 -136
rect 1299 -278 1333 -136
rect 1806 -136 2854 -102
rect 1377 -240 1387 -188
rect 1439 -240 1449 -188
rect 429 -290 475 -278
rect 429 -370 435 -290
rect 469 -370 475 -290
rect 429 -382 475 -370
rect 525 -290 571 -278
rect 525 -370 531 -290
rect 565 -370 571 -290
rect 525 -382 571 -370
rect 621 -290 667 -278
rect 621 -370 627 -290
rect 661 -370 667 -290
rect 621 -382 667 -370
rect 717 -290 763 -278
rect 717 -370 723 -290
rect 757 -370 763 -290
rect 717 -382 763 -370
rect 813 -290 859 -278
rect 813 -370 819 -290
rect 853 -370 859 -290
rect 813 -382 859 -370
rect 909 -290 955 -278
rect 909 -370 915 -290
rect 949 -370 955 -290
rect 909 -382 955 -370
rect 1005 -290 1051 -278
rect 1005 -370 1011 -290
rect 1045 -370 1051 -290
rect 1005 -382 1051 -370
rect 1101 -290 1147 -278
rect 1101 -370 1107 -290
rect 1141 -370 1147 -290
rect 1101 -382 1147 -370
rect 1197 -290 1243 -278
rect 1197 -370 1203 -290
rect 1237 -370 1243 -290
rect 1197 -382 1243 -370
rect 1293 -290 1339 -278
rect 1293 -370 1299 -290
rect 1333 -370 1339 -290
rect 1293 -382 1339 -370
rect 1389 -290 1435 -278
rect 1389 -370 1395 -290
rect 1429 -370 1435 -290
rect 1389 -382 1435 -370
rect 1503 -285 1549 -273
rect 1609 -285 1655 -284
rect 70 -547 319 -503
rect -2236 -688 -2202 -547
rect -2044 -688 -2010 -547
rect -1852 -688 -1818 -547
rect -1660 -688 -1626 -547
rect -1468 -688 -1434 -547
rect -1276 -688 -1242 -547
rect 71 -555 319 -547
rect -702 -620 -614 -614
rect -702 -684 -690 -620
rect -626 -684 -614 -620
rect -2242 -700 -2196 -688
rect -2242 -948 -2236 -700
rect -2202 -948 -2196 -700
rect -2242 -960 -2196 -948
rect -2146 -700 -2100 -688
rect -2146 -948 -2140 -700
rect -2106 -948 -2100 -700
rect -2146 -960 -2100 -948
rect -2050 -700 -2004 -688
rect -2050 -948 -2044 -700
rect -2010 -948 -2004 -700
rect -2050 -960 -2004 -948
rect -1954 -700 -1908 -688
rect -1954 -948 -1948 -700
rect -1914 -948 -1908 -700
rect -1954 -960 -1908 -948
rect -1858 -700 -1812 -688
rect -1858 -948 -1852 -700
rect -1818 -948 -1812 -700
rect -1858 -960 -1812 -948
rect -1762 -700 -1716 -688
rect -1762 -948 -1756 -700
rect -1722 -948 -1716 -700
rect -1762 -960 -1716 -948
rect -1666 -700 -1620 -688
rect -1666 -948 -1660 -700
rect -1626 -948 -1620 -700
rect -1666 -960 -1620 -948
rect -1570 -700 -1524 -688
rect -1570 -948 -1564 -700
rect -1530 -948 -1524 -700
rect -1570 -960 -1524 -948
rect -1474 -700 -1428 -688
rect -1474 -948 -1468 -700
rect -1434 -948 -1428 -700
rect -1474 -960 -1428 -948
rect -1378 -700 -1332 -688
rect -1378 -948 -1372 -700
rect -1338 -948 -1332 -700
rect -1378 -960 -1332 -948
rect -1282 -700 -1236 -688
rect -702 -690 -614 -684
rect -551 -635 -183 -604
rect -551 -669 -522 -635
rect -488 -669 -430 -635
rect -396 -669 -338 -635
rect -304 -669 -246 -635
rect -212 -669 -183 -635
rect -551 -700 -183 -669
rect -1282 -948 -1276 -700
rect -1242 -948 -1236 -700
rect -43 -772 -33 -769
rect -310 -778 -33 -772
rect -310 -812 -298 -778
rect -264 -812 -33 -778
rect -310 -818 -33 -812
rect -43 -821 -33 -818
rect 19 -821 29 -769
rect -401 -917 -391 -865
rect -339 -917 -329 -865
rect -1282 -960 -1236 -948
rect -2140 -1110 -2106 -960
rect -1948 -1110 -1914 -960
rect -1756 -1110 -1722 -960
rect -1564 -1110 -1530 -960
rect -1372 -1110 -1338 -960
rect 139 -1000 149 -997
rect -1298 -1052 -1288 -1000
rect -1236 -1052 -1226 -1000
rect -176 -1052 -166 -1000
rect -114 -1049 149 -1000
rect 201 -1049 211 -997
rect -114 -1052 198 -1049
rect -2386 -1144 -1338 -1110
rect 285 -1110 319 -555
rect 435 -513 469 -382
rect 627 -513 661 -382
rect 819 -513 853 -382
rect 1011 -513 1045 -382
rect 1203 -513 1237 -382
rect 1395 -513 1429 -382
rect 1503 -385 1509 -285
rect 1543 -296 1655 -285
rect 1543 -372 1615 -296
rect 1649 -372 1655 -296
rect 1543 -384 1655 -372
rect 1697 -285 1743 -284
rect 1806 -285 1840 -136
rect 1938 -240 1948 -188
rect 2000 -240 2010 -188
rect 2052 -278 2086 -136
rect 2244 -278 2278 -136
rect 2436 -278 2470 -136
rect 2628 -278 2662 -136
rect 2820 -278 2854 -136
rect 2898 -240 2908 -188
rect 2960 -240 2970 -188
rect 1697 -296 1840 -285
rect 1697 -372 1703 -296
rect 1737 -372 1840 -296
rect 1697 -384 1840 -372
rect 1950 -290 1996 -278
rect 1950 -370 1956 -290
rect 1990 -370 1996 -290
rect 1950 -382 1996 -370
rect 2046 -290 2092 -278
rect 2046 -370 2052 -290
rect 2086 -370 2092 -290
rect 2046 -382 2092 -370
rect 2142 -290 2188 -278
rect 2142 -370 2148 -290
rect 2182 -370 2188 -290
rect 2142 -382 2188 -370
rect 2238 -290 2284 -278
rect 2238 -370 2244 -290
rect 2278 -370 2284 -290
rect 2238 -382 2284 -370
rect 2334 -290 2380 -278
rect 2334 -370 2340 -290
rect 2374 -370 2380 -290
rect 2334 -382 2380 -370
rect 2430 -290 2476 -278
rect 2430 -370 2436 -290
rect 2470 -370 2476 -290
rect 2430 -382 2476 -370
rect 2526 -290 2572 -278
rect 2526 -370 2532 -290
rect 2566 -370 2572 -290
rect 2526 -382 2572 -370
rect 2622 -290 2668 -278
rect 2622 -370 2628 -290
rect 2662 -370 2668 -290
rect 2622 -382 2668 -370
rect 2718 -290 2764 -278
rect 2718 -370 2724 -290
rect 2758 -370 2764 -290
rect 2718 -382 2764 -370
rect 2814 -290 2860 -278
rect 2814 -370 2820 -290
rect 2854 -370 2860 -290
rect 2814 -382 2860 -370
rect 2910 -290 2956 -278
rect 2910 -370 2916 -290
rect 2950 -370 2956 -290
rect 2910 -382 2956 -370
rect 1543 -385 1649 -384
rect 1703 -385 1840 -384
rect 1503 -397 1549 -385
rect 1647 -422 1705 -416
rect 1647 -423 1659 -422
rect 1693 -423 1705 -422
rect 1640 -475 1650 -423
rect 1702 -475 1712 -423
rect 1806 -513 1840 -385
rect 435 -547 1840 -513
rect 435 -688 469 -547
rect 627 -688 661 -547
rect 819 -688 853 -547
rect 1011 -688 1045 -547
rect 1203 -688 1237 -547
rect 1395 -688 1429 -547
rect 429 -700 475 -688
rect 429 -948 435 -700
rect 469 -948 475 -700
rect 429 -960 475 -948
rect 525 -700 571 -688
rect 525 -948 531 -700
rect 565 -948 571 -700
rect 525 -960 571 -948
rect 621 -700 667 -688
rect 621 -948 627 -700
rect 661 -948 667 -700
rect 621 -960 667 -948
rect 717 -700 763 -688
rect 717 -948 723 -700
rect 757 -948 763 -700
rect 717 -960 763 -948
rect 813 -700 859 -688
rect 813 -948 819 -700
rect 853 -948 859 -700
rect 813 -960 859 -948
rect 909 -700 955 -688
rect 909 -948 915 -700
rect 949 -948 955 -700
rect 909 -960 955 -948
rect 1005 -700 1051 -688
rect 1005 -948 1011 -700
rect 1045 -948 1051 -700
rect 1005 -960 1051 -948
rect 1101 -700 1147 -688
rect 1101 -948 1107 -700
rect 1141 -948 1147 -700
rect 1101 -960 1147 -948
rect 1197 -700 1243 -688
rect 1197 -948 1203 -700
rect 1237 -948 1243 -700
rect 1197 -960 1243 -948
rect 1293 -700 1339 -688
rect 1293 -948 1299 -700
rect 1333 -948 1339 -700
rect 1293 -960 1339 -948
rect 1389 -700 1435 -688
rect 1389 -948 1395 -700
rect 1429 -948 1435 -700
rect 1389 -960 1435 -948
rect 416 -1051 426 -999
rect 478 -1051 488 -999
rect 531 -1110 565 -960
rect 723 -1110 757 -960
rect 915 -1110 949 -960
rect 1107 -1110 1141 -960
rect 1299 -1110 1333 -960
rect 1375 -1052 1385 -1000
rect 1437 -1052 1447 -1000
rect 285 -1144 1333 -1110
rect 1806 -1110 1840 -547
rect 1956 -513 1990 -382
rect 2148 -513 2182 -382
rect 2340 -513 2374 -382
rect 2532 -513 2566 -382
rect 2724 -513 2758 -382
rect 2916 -513 2950 -382
rect 1956 -547 3258 -513
rect 1956 -688 1990 -547
rect 2148 -688 2182 -547
rect 2340 -688 2374 -547
rect 2532 -688 2566 -547
rect 2724 -688 2758 -547
rect 2916 -688 2950 -547
rect 1950 -700 1996 -688
rect 1950 -948 1956 -700
rect 1990 -948 1996 -700
rect 1950 -960 1996 -948
rect 2046 -700 2092 -688
rect 2046 -948 2052 -700
rect 2086 -948 2092 -700
rect 2046 -960 2092 -948
rect 2142 -700 2188 -688
rect 2142 -948 2148 -700
rect 2182 -948 2188 -700
rect 2142 -960 2188 -948
rect 2238 -700 2284 -688
rect 2238 -948 2244 -700
rect 2278 -948 2284 -700
rect 2238 -960 2284 -948
rect 2334 -700 2380 -688
rect 2334 -948 2340 -700
rect 2374 -948 2380 -700
rect 2334 -960 2380 -948
rect 2430 -700 2476 -688
rect 2430 -948 2436 -700
rect 2470 -948 2476 -700
rect 2430 -960 2476 -948
rect 2526 -700 2572 -688
rect 2526 -948 2532 -700
rect 2566 -948 2572 -700
rect 2526 -960 2572 -948
rect 2622 -700 2668 -688
rect 2622 -948 2628 -700
rect 2662 -948 2668 -700
rect 2622 -960 2668 -948
rect 2718 -700 2764 -688
rect 2718 -948 2724 -700
rect 2758 -948 2764 -700
rect 2718 -960 2764 -948
rect 2814 -700 2860 -688
rect 2814 -948 2820 -700
rect 2854 -948 2860 -700
rect 2814 -960 2860 -948
rect 2910 -700 2956 -688
rect 2910 -948 2916 -700
rect 2950 -948 2956 -700
rect 2910 -960 2956 -948
rect 1936 -1052 1946 -1000
rect 1998 -1052 2008 -1000
rect 2052 -1110 2086 -960
rect 2244 -1110 2278 -960
rect 2436 -1110 2470 -960
rect 2628 -1110 2662 -960
rect 2820 -1110 2854 -960
rect 2896 -1052 2906 -1000
rect 2958 -1052 2968 -1000
rect 1806 -1144 2854 -1110
rect -551 -1179 -183 -1148
rect -551 -1213 -522 -1179
rect -488 -1213 -430 -1179
rect -396 -1213 -338 -1179
rect -304 -1213 -246 -1179
rect -212 -1213 -183 -1179
rect -551 -1244 -183 -1213
rect -2386 -1284 -1338 -1250
rect -2386 -1847 -2352 -1284
rect -2140 -1434 -2106 -1284
rect -1948 -1434 -1914 -1284
rect -1756 -1434 -1722 -1284
rect -1564 -1434 -1530 -1284
rect -1372 -1434 -1338 -1284
rect 3224 -1270 3258 -547
rect 3224 -1304 3429 -1270
rect -1295 -1395 -1285 -1343
rect -1233 -1395 -1223 -1343
rect -1025 -1394 -1015 -1342
rect -963 -1348 -253 -1342
rect -963 -1382 -299 -1348
rect -265 -1382 -253 -1348
rect -963 -1388 -253 -1382
rect -963 -1394 -953 -1388
rect -2242 -1446 -2196 -1434
rect -2242 -1694 -2236 -1446
rect -2202 -1694 -2196 -1446
rect -2242 -1706 -2196 -1694
rect -2146 -1446 -2100 -1434
rect -2146 -1694 -2140 -1446
rect -2106 -1694 -2100 -1446
rect -2146 -1706 -2100 -1694
rect -2050 -1446 -2004 -1434
rect -2050 -1694 -2044 -1446
rect -2010 -1694 -2004 -1446
rect -2050 -1706 -2004 -1694
rect -1954 -1446 -1908 -1434
rect -1954 -1694 -1948 -1446
rect -1914 -1694 -1908 -1446
rect -1954 -1706 -1908 -1694
rect -1858 -1446 -1812 -1434
rect -1858 -1694 -1852 -1446
rect -1818 -1694 -1812 -1446
rect -1858 -1706 -1812 -1694
rect -1762 -1446 -1716 -1434
rect -1762 -1694 -1756 -1446
rect -1722 -1694 -1716 -1446
rect -1762 -1706 -1716 -1694
rect -1666 -1446 -1620 -1434
rect -1666 -1694 -1660 -1446
rect -1626 -1694 -1620 -1446
rect -1666 -1706 -1620 -1694
rect -1570 -1446 -1524 -1434
rect -1570 -1694 -1564 -1446
rect -1530 -1694 -1524 -1446
rect -1570 -1706 -1524 -1694
rect -1474 -1446 -1428 -1434
rect -1474 -1694 -1468 -1446
rect -1434 -1694 -1428 -1446
rect -1474 -1706 -1428 -1694
rect -1378 -1446 -1332 -1434
rect -1378 -1694 -1372 -1446
rect -1338 -1694 -1332 -1446
rect -1378 -1706 -1332 -1694
rect -1282 -1446 -1236 -1434
rect -1282 -1694 -1276 -1446
rect -1242 -1694 -1236 -1446
rect 285 -1470 1333 -1436
rect -401 -1530 -391 -1478
rect -339 -1530 -329 -1478
rect -1282 -1706 -1236 -1694
rect -2638 -1881 -2352 -1847
rect -2386 -2258 -2352 -1881
rect -2236 -1847 -2202 -1706
rect -2044 -1847 -2010 -1706
rect -1852 -1847 -1818 -1706
rect -1660 -1847 -1626 -1706
rect -1468 -1847 -1434 -1706
rect -1276 -1847 -1242 -1706
rect -702 -1718 -614 -1712
rect -702 -1782 -690 -1718
rect -626 -1782 -614 -1718
rect -702 -1788 -614 -1782
rect -551 -1723 -183 -1692
rect -551 -1757 -522 -1723
rect -488 -1757 -430 -1723
rect -396 -1757 -338 -1723
rect -304 -1757 -246 -1723
rect -212 -1757 -183 -1723
rect -551 -1788 -183 -1757
rect 285 -1837 319 -1470
rect 415 -1572 425 -1520
rect 477 -1572 487 -1520
rect 531 -1612 565 -1470
rect 723 -1612 757 -1470
rect 915 -1612 949 -1470
rect 1107 -1612 1141 -1470
rect 1299 -1612 1333 -1470
rect 1806 -1470 2854 -1436
rect 1377 -1574 1387 -1522
rect 1439 -1574 1449 -1522
rect 429 -1624 475 -1612
rect 429 -1704 435 -1624
rect 469 -1704 475 -1624
rect 429 -1716 475 -1704
rect 525 -1624 571 -1612
rect 525 -1704 531 -1624
rect 565 -1704 571 -1624
rect 525 -1716 571 -1704
rect 621 -1624 667 -1612
rect 621 -1704 627 -1624
rect 661 -1704 667 -1624
rect 621 -1716 667 -1704
rect 717 -1624 763 -1612
rect 717 -1704 723 -1624
rect 757 -1704 763 -1624
rect 717 -1716 763 -1704
rect 813 -1624 859 -1612
rect 813 -1704 819 -1624
rect 853 -1704 859 -1624
rect 813 -1716 859 -1704
rect 909 -1624 955 -1612
rect 909 -1704 915 -1624
rect 949 -1704 955 -1624
rect 909 -1716 955 -1704
rect 1005 -1624 1051 -1612
rect 1005 -1704 1011 -1624
rect 1045 -1704 1051 -1624
rect 1005 -1716 1051 -1704
rect 1101 -1624 1147 -1612
rect 1101 -1704 1107 -1624
rect 1141 -1704 1147 -1624
rect 1101 -1716 1147 -1704
rect 1197 -1624 1243 -1612
rect 1197 -1704 1203 -1624
rect 1237 -1704 1243 -1624
rect 1197 -1716 1243 -1704
rect 1293 -1624 1339 -1612
rect 1293 -1704 1299 -1624
rect 1333 -1704 1339 -1624
rect 1293 -1716 1339 -1704
rect 1389 -1624 1435 -1612
rect 1389 -1704 1395 -1624
rect 1429 -1704 1435 -1624
rect 1389 -1716 1435 -1704
rect 1503 -1619 1549 -1607
rect 1609 -1619 1655 -1618
rect -2236 -1881 -989 -1847
rect -2236 -2012 -2202 -1881
rect -2044 -2012 -2010 -1881
rect -1852 -2012 -1818 -1881
rect -1660 -2012 -1626 -1881
rect -1468 -2012 -1434 -1881
rect -1276 -2012 -1242 -1881
rect -1023 -2007 -989 -1881
rect -875 -1910 -865 -1858
rect -813 -1910 -390 -1858
rect -338 -1910 -328 -1858
rect 69 -1889 319 -1837
rect 69 -2007 103 -1889
rect -2242 -2024 -2196 -2012
rect -2242 -2104 -2236 -2024
rect -2202 -2104 -2196 -2024
rect -2242 -2116 -2196 -2104
rect -2146 -2024 -2100 -2012
rect -2146 -2104 -2140 -2024
rect -2106 -2104 -2100 -2024
rect -2146 -2116 -2100 -2104
rect -2050 -2024 -2004 -2012
rect -2050 -2104 -2044 -2024
rect -2010 -2104 -2004 -2024
rect -2050 -2116 -2004 -2104
rect -1954 -2024 -1908 -2012
rect -1954 -2104 -1948 -2024
rect -1914 -2104 -1908 -2024
rect -1954 -2116 -1908 -2104
rect -1858 -2024 -1812 -2012
rect -1858 -2104 -1852 -2024
rect -1818 -2104 -1812 -2024
rect -1858 -2116 -1812 -2104
rect -1762 -2024 -1716 -2012
rect -1762 -2104 -1756 -2024
rect -1722 -2104 -1716 -2024
rect -1762 -2116 -1716 -2104
rect -1666 -2024 -1620 -2012
rect -1666 -2104 -1660 -2024
rect -1626 -2104 -1620 -2024
rect -1666 -2116 -1620 -2104
rect -1570 -2024 -1524 -2012
rect -1570 -2104 -1564 -2024
rect -1530 -2104 -1524 -2024
rect -1570 -2116 -1524 -2104
rect -1474 -2024 -1428 -2012
rect -1474 -2104 -1468 -2024
rect -1434 -2104 -1428 -2024
rect -1474 -2116 -1428 -2104
rect -1378 -2024 -1332 -2012
rect -1378 -2104 -1372 -2024
rect -1338 -2104 -1332 -2024
rect -1378 -2116 -1332 -2104
rect -1282 -2024 -1236 -2012
rect -1282 -2104 -1276 -2024
rect -1242 -2104 -1236 -2024
rect -1023 -2041 103 -2007
rect -1282 -2116 -1236 -2104
rect -2140 -2258 -2106 -2116
rect -1948 -2258 -1914 -2116
rect -1756 -2258 -1722 -2116
rect -1564 -2258 -1530 -2116
rect -1372 -2258 -1338 -2116
rect -1296 -2206 -1286 -2154
rect -1234 -2206 -1224 -2154
rect -2386 -2292 -1338 -2258
rect 285 -2444 319 -1889
rect 435 -1847 469 -1716
rect 627 -1847 661 -1716
rect 819 -1847 853 -1716
rect 1011 -1847 1045 -1716
rect 1203 -1847 1237 -1716
rect 1395 -1847 1429 -1716
rect 1503 -1719 1509 -1619
rect 1543 -1630 1655 -1619
rect 1543 -1706 1615 -1630
rect 1649 -1706 1655 -1630
rect 1543 -1718 1655 -1706
rect 1697 -1619 1743 -1618
rect 1806 -1619 1840 -1470
rect 1938 -1574 1948 -1522
rect 2000 -1574 2010 -1522
rect 2052 -1612 2086 -1470
rect 2244 -1612 2278 -1470
rect 2436 -1612 2470 -1470
rect 2628 -1612 2662 -1470
rect 2820 -1612 2854 -1470
rect 2898 -1574 2908 -1522
rect 2960 -1574 2970 -1522
rect 1697 -1630 1840 -1619
rect 1697 -1706 1703 -1630
rect 1737 -1706 1840 -1630
rect 1697 -1718 1840 -1706
rect 1950 -1624 1996 -1612
rect 1950 -1704 1956 -1624
rect 1990 -1704 1996 -1624
rect 1950 -1716 1996 -1704
rect 2046 -1624 2092 -1612
rect 2046 -1704 2052 -1624
rect 2086 -1704 2092 -1624
rect 2046 -1716 2092 -1704
rect 2142 -1624 2188 -1612
rect 2142 -1704 2148 -1624
rect 2182 -1704 2188 -1624
rect 2142 -1716 2188 -1704
rect 2238 -1624 2284 -1612
rect 2238 -1704 2244 -1624
rect 2278 -1704 2284 -1624
rect 2238 -1716 2284 -1704
rect 2334 -1624 2380 -1612
rect 2334 -1704 2340 -1624
rect 2374 -1704 2380 -1624
rect 2334 -1716 2380 -1704
rect 2430 -1624 2476 -1612
rect 2430 -1704 2436 -1624
rect 2470 -1704 2476 -1624
rect 2430 -1716 2476 -1704
rect 2526 -1624 2572 -1612
rect 2526 -1704 2532 -1624
rect 2566 -1704 2572 -1624
rect 2526 -1716 2572 -1704
rect 2622 -1624 2668 -1612
rect 2622 -1704 2628 -1624
rect 2662 -1704 2668 -1624
rect 2622 -1716 2668 -1704
rect 2718 -1624 2764 -1612
rect 2718 -1704 2724 -1624
rect 2758 -1704 2764 -1624
rect 2718 -1716 2764 -1704
rect 2814 -1624 2860 -1612
rect 2814 -1704 2820 -1624
rect 2854 -1704 2860 -1624
rect 2814 -1716 2860 -1704
rect 2910 -1624 2956 -1612
rect 2910 -1704 2916 -1624
rect 2950 -1704 2956 -1624
rect 2910 -1716 2956 -1704
rect 1543 -1719 1649 -1718
rect 1703 -1719 1840 -1718
rect 1503 -1731 1549 -1719
rect 1647 -1756 1705 -1750
rect 1647 -1757 1659 -1756
rect 1693 -1757 1705 -1756
rect 1640 -1809 1650 -1757
rect 1702 -1809 1712 -1757
rect 1806 -1847 1840 -1719
rect 435 -1881 1840 -1847
rect 435 -2022 469 -1881
rect 627 -2022 661 -1881
rect 819 -2022 853 -1881
rect 1011 -2022 1045 -1881
rect 1203 -2022 1237 -1881
rect 1395 -2022 1429 -1881
rect 429 -2034 475 -2022
rect 429 -2282 435 -2034
rect 469 -2282 475 -2034
rect 429 -2294 475 -2282
rect 525 -2034 571 -2022
rect 525 -2282 531 -2034
rect 565 -2282 571 -2034
rect 525 -2294 571 -2282
rect 621 -2034 667 -2022
rect 621 -2282 627 -2034
rect 661 -2282 667 -2034
rect 621 -2294 667 -2282
rect 717 -2034 763 -2022
rect 717 -2282 723 -2034
rect 757 -2282 763 -2034
rect 717 -2294 763 -2282
rect 813 -2034 859 -2022
rect 813 -2282 819 -2034
rect 853 -2282 859 -2034
rect 813 -2294 859 -2282
rect 909 -2034 955 -2022
rect 909 -2282 915 -2034
rect 949 -2282 955 -2034
rect 909 -2294 955 -2282
rect 1005 -2034 1051 -2022
rect 1005 -2282 1011 -2034
rect 1045 -2282 1051 -2034
rect 1005 -2294 1051 -2282
rect 1101 -2034 1147 -2022
rect 1101 -2282 1107 -2034
rect 1141 -2282 1147 -2034
rect 1101 -2294 1147 -2282
rect 1197 -2034 1243 -2022
rect 1197 -2282 1203 -2034
rect 1237 -2282 1243 -2034
rect 1197 -2294 1243 -2282
rect 1293 -2034 1339 -2022
rect 1293 -2282 1299 -2034
rect 1333 -2282 1339 -2034
rect 1293 -2294 1339 -2282
rect 1389 -2034 1435 -2022
rect 1389 -2282 1395 -2034
rect 1429 -2282 1435 -2034
rect 1389 -2294 1435 -2282
rect 416 -2385 426 -2333
rect 478 -2385 488 -2333
rect 531 -2444 565 -2294
rect 723 -2444 757 -2294
rect 915 -2444 949 -2294
rect 1107 -2444 1141 -2294
rect 1299 -2444 1333 -2294
rect 1375 -2386 1385 -2334
rect 1437 -2386 1447 -2334
rect 285 -2478 1333 -2444
rect 1806 -2444 1840 -1881
rect 1956 -1847 1990 -1716
rect 2148 -1847 2182 -1716
rect 2340 -1847 2374 -1716
rect 2532 -1847 2566 -1716
rect 2724 -1847 2758 -1716
rect 2916 -1847 2950 -1716
rect 3224 -1847 3258 -1304
rect 1956 -1881 3258 -1847
rect 1956 -2022 1990 -1881
rect 2148 -2022 2182 -1881
rect 2340 -2022 2374 -1881
rect 2532 -2022 2566 -1881
rect 2724 -2022 2758 -1881
rect 2916 -2022 2950 -1881
rect 1950 -2034 1996 -2022
rect 1950 -2282 1956 -2034
rect 1990 -2282 1996 -2034
rect 1950 -2294 1996 -2282
rect 2046 -2034 2092 -2022
rect 2046 -2282 2052 -2034
rect 2086 -2282 2092 -2034
rect 2046 -2294 2092 -2282
rect 2142 -2034 2188 -2022
rect 2142 -2282 2148 -2034
rect 2182 -2282 2188 -2034
rect 2142 -2294 2188 -2282
rect 2238 -2034 2284 -2022
rect 2238 -2282 2244 -2034
rect 2278 -2282 2284 -2034
rect 2238 -2294 2284 -2282
rect 2334 -2034 2380 -2022
rect 2334 -2282 2340 -2034
rect 2374 -2282 2380 -2034
rect 2334 -2294 2380 -2282
rect 2430 -2034 2476 -2022
rect 2430 -2282 2436 -2034
rect 2470 -2282 2476 -2034
rect 2430 -2294 2476 -2282
rect 2526 -2034 2572 -2022
rect 2526 -2282 2532 -2034
rect 2566 -2282 2572 -2034
rect 2526 -2294 2572 -2282
rect 2622 -2034 2668 -2022
rect 2622 -2282 2628 -2034
rect 2662 -2282 2668 -2034
rect 2622 -2294 2668 -2282
rect 2718 -2034 2764 -2022
rect 2718 -2282 2724 -2034
rect 2758 -2282 2764 -2034
rect 2718 -2294 2764 -2282
rect 2814 -2034 2860 -2022
rect 2814 -2282 2820 -2034
rect 2854 -2282 2860 -2034
rect 2814 -2294 2860 -2282
rect 2910 -2034 2956 -2022
rect 2910 -2282 2916 -2034
rect 2950 -2282 2956 -2034
rect 2910 -2294 2956 -2282
rect 1936 -2386 1946 -2334
rect 1998 -2386 2008 -2334
rect 2052 -2444 2086 -2294
rect 2244 -2444 2278 -2294
rect 2436 -2444 2470 -2294
rect 2628 -2444 2662 -2294
rect 2820 -2444 2854 -2294
rect 2896 -2386 2906 -2334
rect 2958 -2386 2968 -2334
rect 1806 -2478 2854 -2444
<< via1 >>
rect -1287 -197 -1235 -188
rect -1287 -231 -1276 -197
rect -1276 -231 -1242 -197
rect -1242 -231 -1235 -197
rect -1287 -240 -1235 -231
rect 425 -197 477 -186
rect 425 -231 435 -197
rect 435 -231 469 -197
rect 469 -231 477 -197
rect 425 -238 477 -231
rect 1387 -197 1439 -188
rect 1387 -231 1395 -197
rect 1395 -231 1429 -197
rect 1429 -231 1439 -197
rect 1387 -240 1439 -231
rect -690 -684 -626 -620
rect -33 -821 19 -769
rect -391 -873 -339 -865
rect -391 -907 -381 -873
rect -381 -907 -347 -873
rect -347 -907 -339 -873
rect -391 -917 -339 -907
rect -1288 -1008 -1236 -1000
rect -1288 -1042 -1276 -1008
rect -1276 -1042 -1242 -1008
rect -1242 -1042 -1236 -1008
rect -1288 -1052 -1236 -1042
rect -166 -1052 -114 -1000
rect 149 -1049 201 -997
rect 1948 -197 2000 -188
rect 1948 -231 1956 -197
rect 1956 -231 1990 -197
rect 1990 -231 2000 -197
rect 1948 -240 2000 -231
rect 2908 -197 2960 -188
rect 2908 -231 2916 -197
rect 2916 -231 2950 -197
rect 2950 -231 2960 -197
rect 2908 -240 2960 -231
rect 1650 -456 1659 -423
rect 1659 -456 1693 -423
rect 1693 -456 1702 -423
rect 1650 -475 1702 -456
rect 426 -1008 478 -999
rect 426 -1042 435 -1008
rect 435 -1042 469 -1008
rect 469 -1042 478 -1008
rect 426 -1051 478 -1042
rect 1385 -1008 1437 -1000
rect 1385 -1042 1395 -1008
rect 1395 -1042 1429 -1008
rect 1429 -1042 1437 -1008
rect 1385 -1052 1437 -1042
rect 1946 -1008 1998 -1000
rect 1946 -1042 1956 -1008
rect 1956 -1042 1990 -1008
rect 1990 -1042 1998 -1008
rect 1946 -1052 1998 -1042
rect 2906 -1008 2958 -1000
rect 2906 -1042 2916 -1008
rect 2916 -1042 2950 -1008
rect 2950 -1042 2958 -1008
rect 2906 -1052 2958 -1042
rect -1285 -1352 -1233 -1343
rect -1285 -1386 -1276 -1352
rect -1276 -1386 -1242 -1352
rect -1242 -1386 -1233 -1352
rect -1285 -1395 -1233 -1386
rect -1015 -1394 -963 -1342
rect -391 -1486 -339 -1478
rect -391 -1520 -382 -1486
rect -382 -1520 -348 -1486
rect -348 -1520 -339 -1486
rect -391 -1530 -339 -1520
rect -690 -1782 -626 -1718
rect 425 -1531 477 -1520
rect 425 -1565 435 -1531
rect 435 -1565 469 -1531
rect 469 -1565 477 -1531
rect 425 -1572 477 -1565
rect 1387 -1531 1439 -1522
rect 1387 -1565 1395 -1531
rect 1395 -1565 1429 -1531
rect 1429 -1565 1439 -1531
rect 1387 -1574 1439 -1565
rect -865 -1910 -813 -1858
rect -390 -1910 -338 -1858
rect -1286 -2163 -1234 -2154
rect -1286 -2197 -1276 -2163
rect -1276 -2197 -1242 -2163
rect -1242 -2197 -1234 -2163
rect -1286 -2206 -1234 -2197
rect 1948 -1531 2000 -1522
rect 1948 -1565 1956 -1531
rect 1956 -1565 1990 -1531
rect 1990 -1565 2000 -1531
rect 1948 -1574 2000 -1565
rect 2908 -1531 2960 -1522
rect 2908 -1565 2916 -1531
rect 2916 -1565 2950 -1531
rect 2950 -1565 2960 -1531
rect 2908 -1574 2960 -1565
rect 1650 -1790 1659 -1757
rect 1659 -1790 1693 -1757
rect 1693 -1790 1702 -1757
rect 1650 -1809 1702 -1790
rect 426 -2342 478 -2333
rect 426 -2376 435 -2342
rect 435 -2376 469 -2342
rect 469 -2376 478 -2342
rect 426 -2385 478 -2376
rect 1385 -2342 1437 -2334
rect 1385 -2376 1395 -2342
rect 1395 -2376 1429 -2342
rect 1429 -2376 1437 -2342
rect 1385 -2386 1437 -2376
rect 1946 -2342 1998 -2334
rect 1946 -2376 1956 -2342
rect 1956 -2376 1990 -2342
rect 1990 -2376 1998 -2342
rect 1946 -2386 1998 -2376
rect 2906 -2342 2958 -2334
rect 2906 -2376 2916 -2342
rect 2916 -2376 2950 -2342
rect 2950 -2376 2958 -2342
rect 2906 -2386 2958 -2376
<< metal2 >>
rect -1287 -188 -1235 -178
rect -1306 -240 -1287 -192
rect -1235 -240 -813 -192
rect -1306 -244 -813 -240
rect -1287 -250 -1235 -244
rect -1288 -1000 -1236 -990
rect -1312 -1052 -1288 -1000
rect -1236 -1052 -963 -1000
rect -1288 -1062 -1236 -1052
rect -1285 -1342 -1233 -1333
rect -1015 -1342 -963 -1052
rect -1285 -1343 -1015 -1342
rect -1233 -1394 -1015 -1343
rect -1285 -1405 -1233 -1395
rect -1015 -1404 -963 -1394
rect -865 -1858 -813 -244
rect -690 -620 -626 -610
rect -690 -1718 -626 -684
rect -391 -865 -339 115
rect 425 -186 477 -176
rect -391 -1000 -339 -917
rect -33 -238 425 -193
rect 517 -193 583 -181
rect 1387 -188 1439 -178
rect 477 -238 1387 -193
rect -33 -240 1387 -238
rect 1948 -188 2000 -178
rect 1439 -240 1948 -193
rect 2908 -188 2960 -178
rect 2000 -240 2908 -193
rect -33 -245 2960 -240
rect -33 -769 19 -245
rect 425 -248 477 -245
rect 517 -247 583 -245
rect 1387 -250 1439 -245
rect 1948 -250 2000 -245
rect 2908 -250 2960 -245
rect -166 -1000 -114 -990
rect -391 -1052 -166 -1000
rect -166 -1062 -114 -1052
rect -690 -1792 -626 -1782
rect -391 -1478 -339 -1468
rect -1286 -2149 -1234 -2144
rect -865 -2149 -813 -1910
rect -1297 -2154 -813 -2149
rect -1297 -2201 -1286 -2154
rect -1234 -2201 -813 -2154
rect -391 -1848 -339 -1530
rect -391 -1858 -338 -1848
rect -391 -1910 -390 -1858
rect -391 -1920 -338 -1910
rect -1286 -2216 -1234 -2206
rect -391 -2457 -339 -1920
rect -33 -2334 19 -821
rect 1650 -423 1702 -413
rect 149 -997 201 -987
rect 426 -999 478 -989
rect 201 -1049 426 -1000
rect 149 -1051 426 -1049
rect 1385 -1000 1437 -990
rect 1650 -1000 1702 -475
rect 1946 -1000 1998 -990
rect 2906 -1000 2958 -990
rect 478 -1051 1385 -1000
rect 149 -1052 1385 -1051
rect 1437 -1052 1946 -1000
rect 1998 -1052 2906 -1000
rect 2958 -1052 2972 -1000
rect 149 -1527 201 -1052
rect 426 -1061 478 -1052
rect 1385 -1062 1437 -1052
rect 1946 -1062 1998 -1052
rect 2906 -1062 2958 -1052
rect 425 -1520 477 -1510
rect 149 -1572 425 -1527
rect 517 -1527 583 -1515
rect 1387 -1522 1439 -1512
rect 477 -1572 1387 -1527
rect 149 -1574 1387 -1572
rect 1948 -1522 2000 -1512
rect 1439 -1574 1948 -1527
rect 2908 -1522 2960 -1512
rect 2000 -1574 2908 -1527
rect 149 -1579 2960 -1574
rect 149 -1589 201 -1579
rect 425 -1582 477 -1579
rect 517 -1581 583 -1579
rect 1387 -1584 1439 -1579
rect 1948 -1584 2000 -1579
rect 2908 -1584 2960 -1579
rect 1650 -1757 1702 -1747
rect 426 -2333 478 -2323
rect -33 -2385 426 -2334
rect 1385 -2334 1437 -2324
rect 1650 -2334 1702 -1809
rect 1946 -2334 1998 -2324
rect 2906 -2334 2958 -2324
rect 478 -2385 1385 -2334
rect -33 -2386 1385 -2385
rect 1437 -2386 1946 -2334
rect 1998 -2386 2906 -2334
rect 2958 -2386 2972 -2334
rect 426 -2395 478 -2386
rect 1385 -2396 1437 -2386
rect 1946 -2396 1998 -2386
rect 2906 -2396 2958 -2386
<< labels >>
flabel metal1 -2635 -530 -2635 -530 3 FreeSans 400 0 0 0 in0
port 3 e
flabel metal1 -2634 -1864 -2634 -1864 3 FreeSans 400 0 0 0 in1
port 4 e
flabel metal2 -365 -2445 -365 -2445 1 FreeSans 400 0 0 0 en
port 1 n
flabel metal1 3423 -1288 3423 -1288 1 FreeSans 400 0 0 0 out
port 5 n
flabel metal2 -366 110 -366 110 5 FreeSans 400 0 0 0 s0
port 2 s
flabel locali -2575 182 -2575 182 1 FreeSans 400 0 0 0 VDD
port 6 n power bidirectional
flabel locali -2569 -2738 -2569 -2738 1 FreeSans 400 0 0 0 VSS
port 7 n power bidirectional
<< end >>
