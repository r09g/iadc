magic
tech sky130A
magscale 1 2
timestamp 1654752884
<< locali >>
rect 15025 21777 15117 21811
rect 15410 21777 15611 21811
rect 18538 21777 18906 21811
rect 15025 21743 15059 21777
rect 15577 21675 15611 21777
rect 18613 21675 18647 21777
rect 15577 21641 15686 21675
rect 13202 21233 13495 21267
rect 16606 21233 16974 21267
rect 13461 21199 13495 21233
rect 17693 21199 17727 21369
rect 13461 21165 13647 21199
rect 17693 21165 17802 21199
rect 21206 21165 21281 21199
rect 22954 21097 23155 21131
rect 14323 20825 14398 20859
rect 14289 20689 14398 20723
rect 14289 20655 14323 20689
rect 15393 20655 15427 20825
rect 15333 20621 15427 20655
rect 23121 20587 23155 21097
rect 8861 19635 8895 19737
rect 8861 19601 8970 19635
rect 17325 19601 17618 19635
rect 9338 19533 9447 19567
rect 8234 19465 8343 19499
rect 8309 19431 8343 19465
rect 9413 19431 9447 19533
rect 17325 19499 17359 19601
rect 15853 19465 15962 19499
rect 15853 19431 15887 19465
rect 6469 19057 6578 19091
rect 6469 18887 6503 19057
rect 11546 18989 11621 19023
rect 21833 18479 21867 18649
rect 21833 18445 21942 18479
rect 7849 18071 7883 18105
rect 7774 18037 7883 18071
rect 16313 18003 16347 18105
rect 5917 17969 6394 18003
rect 16313 17969 16422 18003
rect 5917 17935 5951 17969
rect 5641 17901 5951 17935
rect 21315 17901 21390 17935
rect 5641 17459 5675 17901
rect 5641 17425 6026 17459
rect 19933 17425 20119 17459
rect 20085 17255 20119 17425
rect 13645 16813 13754 16847
rect 20453 16813 20562 16847
rect 13645 16779 13679 16813
rect 15778 16745 15853 16779
rect 20453 16711 20487 16813
rect 21114 16677 21189 16711
rect 17250 16473 17325 16507
rect 12098 16337 12207 16371
rect 6578 16269 6670 16303
rect 12173 16235 12207 16337
rect 13185 16303 13219 16473
rect 16514 16405 16589 16439
rect 22477 16303 22511 16473
rect 13110 16269 13219 16303
rect 22402 16269 22511 16303
rect 19441 15759 19475 15793
rect 8694 15725 8803 15759
rect 10902 15725 10977 15759
rect 11011 15725 11270 15759
rect 18739 15725 18799 15759
rect 19366 15725 19475 15759
rect 8769 15623 8803 15725
rect 19659 15657 19734 15691
rect 11454 15589 11730 15623
rect 17509 15283 17543 15385
rect 7147 15249 7207 15283
rect 14766 15249 14950 15283
rect 17509 15249 17618 15283
rect 22017 15215 22051 15385
rect 22017 15181 22126 15215
rect 20853 14841 20913 14875
rect 8769 14671 8803 14841
rect 8341 14637 8401 14671
rect 8769 14637 8878 14671
rect 10919 14637 11063 14671
rect 19015 14297 19070 14331
rect 14766 14161 14841 14195
rect 20119 13957 20194 13991
rect 23121 13855 23155 14025
rect 23121 13821 23247 13855
rect 6193 13719 6227 13753
rect 6193 13685 6302 13719
rect 7222 13617 7314 13651
rect 12817 13583 12851 13685
rect 12742 13549 12851 13583
rect 6285 12087 6319 12121
rect 6285 12053 6394 12087
rect 16345 12053 16405 12087
rect 16054 11373 16255 11407
rect 16221 11271 16255 11373
rect 20395 11305 20470 11339
rect 23213 11067 23247 13821
rect 23489 11815 23523 18853
rect 23121 11033 23247 11067
rect 23397 11781 23523 11815
rect 23121 10863 23155 11033
rect 6561 10761 6670 10795
rect 6561 10727 6595 10761
rect 23397 10659 23431 11781
rect 23673 11679 23707 11849
rect 23627 11645 23707 11679
rect 23627 10659 23661 11645
rect 23305 10625 23431 10659
rect 23581 10625 23661 10659
rect 6561 10319 6595 10421
rect 18337 10319 18371 10489
rect 20913 10319 20947 10353
rect 6486 10285 6595 10319
rect 18262 10285 18371 10319
rect 20853 10285 20947 10319
rect 11753 10217 11805 10251
rect 6193 9843 6227 9945
rect 6745 9843 6779 9945
rect 6118 9809 6227 9843
rect 6285 9809 6394 9843
rect 6670 9809 6779 9843
rect 6285 9707 6319 9809
rect 19366 9741 19475 9775
rect 6118 9673 6319 9707
rect 19441 9639 19475 9741
rect 23305 9639 23339 10625
rect 23581 9775 23615 10625
rect 23765 9911 23799 19669
rect 23857 11203 23891 11373
rect 23857 11169 23937 11203
rect 23903 10523 23937 11169
rect 24041 10727 24075 10897
rect 24041 10693 24259 10727
rect 23903 10489 23983 10523
rect 23949 9775 23983 10489
rect 23581 9741 23707 9775
rect 23305 9605 23431 9639
rect 18262 9197 18371 9231
rect 20853 9197 20947 9231
rect 18337 9095 18371 9197
rect 20913 9095 20947 9197
rect 6854 8721 6929 8755
rect 7021 8721 7207 8755
rect 12098 8721 12391 8755
rect 7021 8551 7055 8721
rect 12357 8687 12391 8721
rect 12357 8653 12635 8687
rect 17509 8551 17543 8857
rect 6285 8279 6319 8313
rect 6285 8245 6394 8279
rect 20913 8143 20947 8313
rect 13294 8109 13647 8143
rect 20838 8109 20947 8143
rect 13461 8007 13495 8109
rect 23397 7939 23431 9605
rect 23397 7905 23523 7939
rect 5641 7769 5842 7803
rect 6854 7769 6929 7803
rect 5549 6579 5583 7021
rect 5641 6919 5675 7769
rect 23489 7735 23523 7905
rect 5733 7633 5842 7667
rect 6026 7633 6135 7667
rect 5733 7463 5767 7633
rect 6101 7463 6135 7633
rect 19826 7565 19935 7599
rect 19901 7531 19935 7565
rect 23673 7531 23707 9741
rect 12098 7497 12207 7531
rect 23581 7497 23707 7531
rect 23857 9741 23983 9775
rect 12173 7463 12207 7497
rect 18262 7089 18371 7123
rect 15594 6953 15761 6987
rect 18337 6919 18371 7089
rect 21114 7021 21189 7055
rect 23581 6919 23615 7497
rect 23857 7055 23891 9741
rect 24225 9639 24259 10693
rect 24133 9605 24259 9639
rect 24133 6919 24167 9605
rect 23581 6885 23707 6919
rect 23673 6715 23707 6885
rect 24041 6885 24167 6919
rect 7481 6579 7515 6613
rect 5549 6545 6026 6579
rect 6302 6545 6411 6579
rect 7481 6545 7573 6579
rect 6377 6511 6411 6545
rect 24041 6443 24075 6885
rect 18001 6137 18061 6171
rect 7757 6103 7791 6137
rect 7757 6069 7866 6103
rect 10425 5967 10459 6137
rect 13645 6069 13754 6103
rect 13645 5967 13679 6069
rect 17509 6001 17618 6035
rect 17509 5967 17543 6001
rect 10425 5933 10534 5967
rect 13478 5933 13679 5967
rect 17250 5933 17543 5967
<< viali >>
rect 18429 21913 18463 21947
rect 15209 21845 15243 21879
rect 18981 21845 19015 21879
rect 19165 21845 19199 21879
rect 15117 21777 15151 21811
rect 15669 21777 15703 21811
rect 15853 21777 15887 21811
rect 18337 21777 18371 21811
rect 20269 21777 20303 21811
rect 20545 21777 20579 21811
rect 21005 21777 21039 21811
rect 22661 21777 22695 21811
rect 22845 21777 22879 21811
rect 10333 21709 10367 21743
rect 15025 21709 15059 21743
rect 19717 21709 19751 21743
rect 20453 21709 20487 21743
rect 20913 21709 20947 21743
rect 21741 21709 21775 21743
rect 22017 21709 22051 21743
rect 10149 21641 10183 21675
rect 18613 21641 18647 21675
rect 19533 21641 19567 21675
rect 20085 21641 20119 21675
rect 22753 21641 22787 21675
rect 10517 21573 10551 21607
rect 15393 21573 15427 21607
rect 15669 21573 15703 21607
rect 19165 21573 19199 21607
rect 19901 21573 19935 21607
rect 20729 21573 20763 21607
rect 21557 21573 21591 21607
rect 22385 21573 22419 21607
rect 10149 21369 10183 21403
rect 15945 21369 15979 21403
rect 17325 21369 17359 21403
rect 17693 21369 17727 21403
rect 18153 21369 18187 21403
rect 21465 21369 21499 21403
rect 14013 21233 14047 21267
rect 16405 21233 16439 21267
rect 17417 21233 17451 21267
rect 19257 21301 19291 21335
rect 19717 21301 19751 21335
rect 22492 21301 22526 21335
rect 19073 21233 19107 21267
rect 19533 21233 19567 21267
rect 13001 21165 13035 21199
rect 13829 21165 13863 21199
rect 14105 21165 14139 21199
rect 15761 21165 15795 21199
rect 17141 21165 17175 21199
rect 17969 21165 18003 21199
rect 19809 21165 19843 21199
rect 21281 21165 21315 21199
rect 15500 21097 15534 21131
rect 17877 21097 17911 21131
rect 20065 21088 20099 21122
rect 10057 21029 10091 21063
rect 12817 21029 12851 21063
rect 14381 21029 14415 21063
rect 15853 21029 15887 21063
rect 16221 21029 16255 21063
rect 18061 21029 18095 21063
rect 18889 21029 18923 21063
rect 19349 21029 19383 21063
rect 14289 20825 14323 20859
rect 15393 20825 15427 20859
rect 21465 20825 21499 20859
rect 10900 20767 10934 20801
rect 12618 20767 12652 20801
rect 7558 20689 7592 20723
rect 11161 20689 11195 20723
rect 12357 20689 12391 20723
rect 14565 20689 14599 20723
rect 15117 20689 15151 20723
rect 16206 20757 16240 20791
rect 18904 20757 18938 20791
rect 20346 20757 20380 20791
rect 21925 20689 21959 20723
rect 7297 20621 7331 20655
rect 14289 20621 14323 20655
rect 15945 20621 15979 20655
rect 19165 20621 19199 20655
rect 20085 20621 20119 20655
rect 21741 20621 21775 20655
rect 21557 20553 21591 20587
rect 23121 20553 23155 20587
rect 8677 20485 8711 20519
rect 9781 20485 9815 20519
rect 13737 20485 13771 20519
rect 14933 20485 14967 20519
rect 17325 20485 17359 20519
rect 17785 20485 17819 20519
rect 11069 20281 11103 20315
rect 6837 20145 6871 20179
rect 10517 20145 10551 20179
rect 22937 20145 22971 20179
rect 12449 20077 12483 20111
rect 15577 20077 15611 20111
rect 16221 20077 16255 20111
rect 20177 20077 20211 20111
rect 7098 20009 7132 20043
rect 10256 20009 10290 20043
rect 12188 20009 12222 20043
rect 15316 20009 15350 20043
rect 16482 20009 16516 20043
rect 19916 20009 19950 20043
rect 22676 20009 22710 20043
rect 8217 19941 8251 19975
rect 9137 19941 9171 19975
rect 14197 19941 14231 19975
rect 17601 19941 17635 19975
rect 18797 19941 18831 19975
rect 21557 19941 21591 19975
rect 7849 19737 7883 19771
rect 8861 19737 8895 19771
rect 9137 19737 9171 19771
rect 10333 19737 10367 19771
rect 15485 19737 15519 19771
rect 16313 19737 16347 19771
rect 16773 19737 16807 19771
rect 21097 19737 21131 19771
rect 9045 19669 9079 19703
rect 12725 19669 12759 19703
rect 13078 19669 13112 19703
rect 22216 19669 22250 19703
rect 23765 19669 23799 19703
rect 8033 19601 8067 19635
rect 10517 19601 10551 19635
rect 11989 19601 12023 19635
rect 12541 19601 12575 19635
rect 12817 19601 12851 19635
rect 15301 19601 15335 19635
rect 16129 19601 16163 19635
rect 16589 19601 16623 19635
rect 9045 19465 9079 19499
rect 8309 19397 8343 19431
rect 22477 19533 22511 19567
rect 10701 19465 10735 19499
rect 12357 19465 12391 19499
rect 15117 19465 15151 19499
rect 16405 19465 16439 19499
rect 17325 19465 17359 19499
rect 18038 19465 18072 19499
rect 9413 19397 9447 19431
rect 11897 19397 11931 19431
rect 14197 19397 14231 19431
rect 15853 19397 15887 19431
rect 19073 19397 19107 19431
rect 6929 19193 6963 19227
rect 10333 19193 10367 19227
rect 15945 19193 15979 19227
rect 21097 19193 21131 19227
rect 10517 19125 10551 19159
rect 11253 19125 11287 19159
rect 12334 19125 12368 19159
rect 13369 19125 13403 19159
rect 14910 19125 14944 19159
rect 20062 19125 20096 19159
rect 9689 19057 9723 19091
rect 9965 19057 9999 19091
rect 11713 19057 11747 19091
rect 11989 19057 12023 19091
rect 14565 19057 14599 19091
rect 6745 18989 6779 19023
rect 10701 18989 10735 19023
rect 11253 18989 11287 19023
rect 11621 18989 11655 19023
rect 11805 18989 11839 19023
rect 17233 18989 17267 19023
rect 17494 18989 17528 19023
rect 22845 18989 22879 19023
rect 11437 18921 11471 18955
rect 22584 18921 22618 18955
rect 6469 18853 6503 18887
rect 9505 18853 9539 18887
rect 10885 18853 10919 18887
rect 18613 18853 18647 18887
rect 19717 18853 19751 18887
rect 21465 18853 21499 18887
rect 23489 18853 23523 18887
rect 6101 18649 6135 18683
rect 8309 18649 8343 18683
rect 12081 18649 12115 18683
rect 12541 18649 12575 18683
rect 19809 18649 19843 18683
rect 21833 18649 21867 18683
rect 22293 18649 22327 18683
rect 14013 18581 14047 18615
rect 17064 18581 17098 18615
rect 17693 18581 17727 18615
rect 17785 18581 17819 18615
rect 20346 18581 20380 18615
rect 6745 18513 6779 18547
rect 7665 18513 7699 18547
rect 10962 18513 10996 18547
rect 17509 18513 17543 18547
rect 17877 18513 17911 18547
rect 19349 18513 19383 18547
rect 22109 18513 22143 18547
rect 6653 18445 6687 18479
rect 7941 18445 7975 18479
rect 8769 18445 8803 18479
rect 9045 18445 9079 18479
rect 10701 18445 10735 18479
rect 17325 18445 17359 18479
rect 19625 18445 19659 18479
rect 20085 18445 20119 18479
rect 7481 18377 7515 18411
rect 8585 18377 8619 18411
rect 12886 18377 12920 18411
rect 6929 18309 6963 18343
rect 9413 18309 9447 18343
rect 15945 18309 15979 18343
rect 18061 18309 18095 18343
rect 18981 18309 19015 18343
rect 21465 18309 21499 18343
rect 7849 18105 7883 18139
rect 9689 18105 9723 18139
rect 16313 18105 16347 18139
rect 21189 18105 21223 18139
rect 6745 18037 6779 18071
rect 13024 18037 13058 18071
rect 16037 18037 16071 18071
rect 17693 18037 17727 18071
rect 9965 17969 9999 18003
rect 11805 17969 11839 18003
rect 11897 17969 11931 18003
rect 16589 17969 16623 18003
rect 22753 17969 22787 18003
rect 6561 17901 6595 17935
rect 7573 17901 7607 17935
rect 9873 17901 9907 17935
rect 11621 17901 11655 17935
rect 14013 17901 14047 17935
rect 15485 17901 15519 17935
rect 15761 17901 15795 17935
rect 15853 17901 15887 17935
rect 19809 17901 19843 17935
rect 20070 17901 20104 17935
rect 21281 17901 21315 17935
rect 22492 17901 22526 17935
rect 14274 17833 14308 17867
rect 15669 17833 15703 17867
rect 7389 17765 7423 17799
rect 10517 17765 10551 17799
rect 11437 17765 11471 17799
rect 13369 17765 13403 17799
rect 15393 17765 15427 17799
rect 21189 17765 21223 17799
rect 12173 17561 12207 17595
rect 14749 17561 14783 17595
rect 9413 17493 9447 17527
rect 13630 17493 13664 17527
rect 15393 17493 15427 17527
rect 19717 17493 19751 17527
rect 7205 17425 7239 17459
rect 7466 17425 7500 17459
rect 9137 17425 9171 17459
rect 9229 17425 9263 17459
rect 10425 17425 10459 17459
rect 10793 17425 10827 17459
rect 11054 17425 11088 17459
rect 12909 17425 12943 17459
rect 13093 17425 13127 17459
rect 13369 17425 13403 17459
rect 15301 17425 15335 17459
rect 15485 17425 15519 17459
rect 15669 17425 15703 17459
rect 17877 17425 17911 17459
rect 18138 17425 18172 17459
rect 19533 17425 19567 17459
rect 19625 17425 19659 17459
rect 22216 17425 22250 17459
rect 22477 17425 22511 17459
rect 6561 17357 6595 17391
rect 6653 17357 6687 17391
rect 10241 17357 10275 17391
rect 13277 17289 13311 17323
rect 19257 17289 19291 17323
rect 21097 17289 21131 17323
rect 6837 17221 6871 17255
rect 8585 17221 8619 17255
rect 9137 17221 9171 17255
rect 10609 17221 10643 17255
rect 15117 17221 15151 17255
rect 19349 17221 19383 17255
rect 20085 17221 20119 17255
rect 9505 17017 9539 17051
rect 11345 17017 11379 17051
rect 11989 17017 12023 17051
rect 14289 17017 14323 17051
rect 16773 17017 16807 17051
rect 20177 17017 20211 17051
rect 13016 16949 13050 16983
rect 10885 16881 10919 16915
rect 11713 16881 11747 16915
rect 18153 16881 18187 16915
rect 18797 16881 18831 16915
rect 10624 16813 10658 16847
rect 11529 16813 11563 16847
rect 11805 16813 11839 16847
rect 13921 16813 13955 16847
rect 14013 16813 14047 16847
rect 14105 16813 14139 16847
rect 14381 16813 14415 16847
rect 14642 16813 14676 16847
rect 19058 16813 19092 16847
rect 20913 16813 20947 16847
rect 13645 16745 13679 16779
rect 15853 16745 15887 16779
rect 17892 16745 17926 16779
rect 20729 16745 20763 16779
rect 20821 16745 20855 16779
rect 13369 16677 13403 16711
rect 20453 16677 20487 16711
rect 21189 16677 21223 16711
rect 8769 16473 8803 16507
rect 11805 16473 11839 16507
rect 13185 16473 13219 16507
rect 13369 16473 13403 16507
rect 17325 16473 17359 16507
rect 19901 16473 19935 16507
rect 21465 16473 21499 16507
rect 22017 16473 22051 16507
rect 22477 16473 22511 16507
rect 7021 16405 7055 16439
rect 7650 16405 7684 16439
rect 10600 16415 10634 16449
rect 6193 16337 6227 16371
rect 6837 16337 6871 16371
rect 7389 16337 7423 16371
rect 9045 16337 9079 16371
rect 9137 16337 9171 16371
rect 10333 16337 10367 16371
rect 11805 16337 11839 16371
rect 11897 16337 11931 16371
rect 12909 16337 12943 16371
rect 6285 16269 6319 16303
rect 8861 16269 8895 16303
rect 9413 16269 9447 16303
rect 9965 16269 9999 16303
rect 14488 16405 14522 16439
rect 15378 16405 15412 16439
rect 16589 16405 16623 16439
rect 16865 16405 16899 16439
rect 16957 16405 16991 16439
rect 18782 16405 18816 16439
rect 20346 16405 20380 16439
rect 14749 16337 14783 16371
rect 15117 16337 15151 16371
rect 16681 16337 16715 16371
rect 17049 16337 17083 16371
rect 20085 16337 20119 16371
rect 18521 16269 18555 16303
rect 22201 16269 22235 16303
rect 9229 16201 9263 16235
rect 9781 16201 9815 16235
rect 11713 16201 11747 16235
rect 12173 16201 12207 16235
rect 8769 16133 8803 16167
rect 9137 16133 9171 16167
rect 9597 16133 9631 16167
rect 10149 16133 10183 16167
rect 12725 16133 12759 16167
rect 21465 16133 21499 16167
rect 8585 15929 8619 15963
rect 9413 15929 9447 15963
rect 11805 15929 11839 15963
rect 13461 15929 13495 15963
rect 9045 15861 9079 15895
rect 16681 15793 16715 15827
rect 19441 15793 19475 15827
rect 22753 15793 22787 15827
rect 6929 15725 6963 15759
rect 8493 15725 8527 15759
rect 9229 15725 9263 15759
rect 9505 15725 9539 15759
rect 9766 15725 9800 15759
rect 10977 15725 11011 15759
rect 11437 15725 11471 15759
rect 12081 15725 12115 15759
rect 14381 15725 14415 15759
rect 16497 15725 16531 15759
rect 18705 15725 18739 15759
rect 18981 15725 19015 15759
rect 19073 15725 19107 15759
rect 20836 15725 20870 15759
rect 21097 15725 21131 15759
rect 7196 15648 7230 15682
rect 12342 15648 12376 15682
rect 14642 15657 14676 15691
rect 19165 15657 19199 15691
rect 19625 15657 19659 15691
rect 22492 15657 22526 15691
rect 8309 15589 8343 15623
rect 8769 15589 8803 15623
rect 11345 15589 11379 15623
rect 15761 15589 15795 15623
rect 17785 15589 17819 15623
rect 21373 15589 21407 15623
rect 6101 15385 6135 15419
rect 9965 15385 9999 15419
rect 16313 15385 16347 15419
rect 17509 15385 17543 15419
rect 8324 15317 8358 15351
rect 9045 15317 9079 15351
rect 12173 15317 12207 15351
rect 15194 15317 15228 15351
rect 16681 15317 16715 15351
rect 22017 15385 22051 15419
rect 21204 15317 21238 15351
rect 6561 15249 6595 15283
rect 7113 15249 7147 15283
rect 8585 15249 8619 15283
rect 8861 15249 8895 15283
rect 10149 15249 10183 15283
rect 10333 15249 10367 15283
rect 16405 15249 16439 15283
rect 16589 15249 16623 15283
rect 16773 15249 16807 15283
rect 18782 15249 18816 15283
rect 6285 15181 6319 15215
rect 10425 15181 10459 15215
rect 10701 15181 10735 15215
rect 13185 15181 13219 15215
rect 18521 15181 18555 15215
rect 21465 15181 21499 15215
rect 22293 15181 22327 15215
rect 6929 15113 6963 15147
rect 8677 15113 8711 15147
rect 11054 15113 11088 15147
rect 13369 15113 13403 15147
rect 14473 15113 14507 15147
rect 20085 15113 20119 15147
rect 16957 15045 16991 15079
rect 19901 15045 19935 15079
rect 22477 15045 22511 15079
rect 8769 14841 8803 14875
rect 10333 14841 10367 14875
rect 17601 14841 17635 14875
rect 20913 14841 20947 14875
rect 6929 14705 6963 14739
rect 9298 14773 9332 14807
rect 13645 14773 13679 14807
rect 21373 14773 21407 14807
rect 18797 14705 18831 14739
rect 22753 14705 22787 14739
rect 7190 14637 7224 14671
rect 8401 14637 8435 14671
rect 10885 14637 10919 14671
rect 12188 14637 12222 14671
rect 12449 14637 12483 14671
rect 13829 14637 13863 14671
rect 14473 14637 14507 14671
rect 16221 14637 16255 14671
rect 16482 14637 16516 14671
rect 18245 14637 18279 14671
rect 18521 14637 18555 14671
rect 20257 14637 20291 14671
rect 20545 14637 20579 14671
rect 20637 14620 20671 14654
rect 22492 14637 22526 14671
rect 14734 14569 14768 14603
rect 19053 14569 19087 14603
rect 20453 14569 20487 14603
rect 8309 14501 8343 14535
rect 14013 14501 14047 14535
rect 15853 14501 15887 14535
rect 20177 14501 20211 14535
rect 10793 14297 10827 14331
rect 14105 14297 14139 14331
rect 17509 14297 17543 14331
rect 18981 14297 19015 14331
rect 22017 14297 22051 14331
rect 12986 14229 13020 14263
rect 14473 14229 14507 14263
rect 6561 14161 6595 14195
rect 7849 14161 7883 14195
rect 8110 14161 8144 14195
rect 11912 14161 11946 14195
rect 14197 14161 14231 14195
rect 14381 14161 14415 14195
rect 14565 14161 14599 14195
rect 14841 14161 14875 14195
rect 16773 14161 16807 14195
rect 18628 14161 18662 14195
rect 18889 14161 18923 14195
rect 19257 14161 19291 14195
rect 19349 14161 19383 14195
rect 19441 14161 19475 14195
rect 19625 14161 19659 14195
rect 21296 14161 21330 14195
rect 21557 14161 21591 14195
rect 22201 14161 22235 14195
rect 6653 14093 6687 14127
rect 12173 14093 12207 14127
rect 12725 14093 12759 14127
rect 16589 14093 16623 14127
rect 15485 14025 15519 14059
rect 22385 14025 22419 14059
rect 23121 14025 23155 14059
rect 6285 13957 6319 13991
rect 9229 13957 9263 13991
rect 10793 13957 10827 13991
rect 20085 13957 20119 13991
rect 6193 13753 6227 13787
rect 6653 13753 6687 13787
rect 7665 13753 7699 13787
rect 9321 13753 9355 13787
rect 11253 13753 11287 13787
rect 16221 13753 16255 13787
rect 18337 13753 18371 13787
rect 20177 13753 20211 13787
rect 10356 13685 10390 13719
rect 12288 13685 12322 13719
rect 12817 13685 12851 13719
rect 13829 13685 13863 13719
rect 20269 13685 20303 13719
rect 21373 13685 21407 13719
rect 6745 13617 6779 13651
rect 12909 13617 12943 13651
rect 17601 13617 17635 13651
rect 18797 13617 18831 13651
rect 22753 13617 22787 13651
rect 6469 13549 6503 13583
rect 6837 13549 6871 13583
rect 7021 13549 7055 13583
rect 7481 13549 7515 13583
rect 13093 13549 13127 13583
rect 14013 13549 14047 13583
rect 18153 13549 18187 13583
rect 20453 13549 20487 13583
rect 20821 13549 20855 13583
rect 22492 13549 22526 13583
rect 17340 13481 17374 13515
rect 19058 13481 19092 13515
rect 20545 13481 20579 13515
rect 20637 13481 20671 13515
rect 10701 13413 10735 13447
rect 13277 13413 13311 13447
rect 14197 13413 14231 13447
rect 6653 13209 6687 13243
rect 8677 13209 8711 13243
rect 14197 13209 14231 13243
rect 15945 13209 15979 13243
rect 20085 13209 20119 13243
rect 10609 13141 10643 13175
rect 12173 13141 12207 13175
rect 13078 13141 13112 13175
rect 15393 13141 15427 13175
rect 15485 13141 15519 13175
rect 18628 13141 18662 13175
rect 21212 13141 21246 13175
rect 21925 13141 21959 13175
rect 6561 13073 6595 13107
rect 6745 13073 6779 13107
rect 7558 13073 7592 13107
rect 10057 13073 10091 13107
rect 15301 13073 15335 13107
rect 15669 13073 15703 13107
rect 17064 13073 17098 13107
rect 17325 13073 17359 13107
rect 18889 13073 18923 13107
rect 21741 13073 21775 13107
rect 21833 13073 21867 13107
rect 22109 13073 22143 13107
rect 7297 13005 7331 13039
rect 10241 13005 10275 13039
rect 10425 13005 10459 13039
rect 12817 13005 12851 13039
rect 14749 13005 14783 13039
rect 21465 13005 21499 13039
rect 11736 12937 11770 12971
rect 15117 12869 15151 12903
rect 17509 12869 17543 12903
rect 21557 12869 21591 12903
rect 8769 12665 8803 12699
rect 11897 12665 11931 12699
rect 17141 12665 17175 12699
rect 22753 12665 22787 12699
rect 9804 12597 9838 12631
rect 13277 12529 13311 12563
rect 18613 12529 18647 12563
rect 6377 12461 6411 12495
rect 6561 12461 6595 12495
rect 7113 12461 7147 12495
rect 13016 12461 13050 12495
rect 13645 12461 13679 12495
rect 13906 12461 13940 12495
rect 16589 12461 16623 12495
rect 16773 12461 16807 12495
rect 16865 12461 16899 12495
rect 16957 12461 16991 12495
rect 20177 12461 20211 12495
rect 21097 12461 21131 12495
rect 21373 12461 21407 12495
rect 6929 12393 6963 12427
rect 18352 12393 18386 12427
rect 21634 12393 21668 12427
rect 6469 12325 6503 12359
rect 10149 12325 10183 12359
rect 15025 12325 15059 12359
rect 17233 12325 17267 12359
rect 6285 12121 6319 12155
rect 6561 12121 6595 12155
rect 8861 12121 8895 12155
rect 14749 12121 14783 12155
rect 21557 12121 21591 12155
rect 10609 12053 10643 12087
rect 13630 12053 13664 12087
rect 15194 12053 15228 12087
rect 16405 12053 16439 12087
rect 16957 12053 16991 12087
rect 17049 12053 17083 12087
rect 17877 12053 17911 12087
rect 17969 12053 18003 12087
rect 18782 12053 18816 12087
rect 6653 11985 6687 12019
rect 7742 11985 7776 12019
rect 9873 11985 9907 12019
rect 13369 11985 13403 12019
rect 14933 11985 14967 12019
rect 16773 11985 16807 12019
rect 17141 11985 17175 12019
rect 17785 11985 17819 12019
rect 18153 11985 18187 12019
rect 21204 11985 21238 12019
rect 7481 11917 7515 11951
rect 10057 11917 10091 11951
rect 10241 11917 10275 11951
rect 12081 11917 12115 11951
rect 18521 11917 18555 11951
rect 21465 11917 21499 11951
rect 21741 11917 21775 11951
rect 11736 11849 11770 11883
rect 17325 11849 17359 11883
rect 21925 11849 21959 11883
rect 6377 11781 6411 11815
rect 17601 11781 17635 11815
rect 19901 11781 19935 11815
rect 20085 11781 20119 11815
rect 8309 11577 8343 11611
rect 10609 11577 10643 11611
rect 13461 11577 13495 11611
rect 6469 11509 6503 11543
rect 9574 11509 9608 11543
rect 11437 11509 11471 11543
rect 20177 11509 20211 11543
rect 14013 11441 14047 11475
rect 22753 11441 22787 11475
rect 6653 11373 6687 11407
rect 6929 11373 6963 11407
rect 11621 11373 11655 11407
rect 12081 11373 12115 11407
rect 14274 11373 14308 11407
rect 15485 11373 15519 11407
rect 15853 11373 15887 11407
rect 16865 11373 16899 11407
rect 17126 11373 17160 11407
rect 18797 11373 18831 11407
rect 20637 11373 20671 11407
rect 21005 11373 21039 11407
rect 22492 11373 22526 11407
rect 6837 11305 6871 11339
rect 7185 11296 7219 11330
rect 11805 11305 11839 11339
rect 12337 11296 12371 11330
rect 15669 11305 15703 11339
rect 15761 11305 15795 11339
rect 19058 11305 19092 11339
rect 20361 11305 20395 11339
rect 20729 11305 20763 11339
rect 20821 11305 20855 11339
rect 9229 11237 9263 11271
rect 15393 11237 15427 11271
rect 16221 11237 16255 11271
rect 18245 11237 18279 11271
rect 21373 11237 21407 11271
rect 11897 11033 11931 11067
rect 14749 11033 14783 11067
rect 19717 11033 19751 11067
rect 23673 11849 23707 11883
rect 10425 10965 10459 10999
rect 13630 10965 13664 10999
rect 21212 10965 21246 10999
rect 6837 10897 6871 10931
rect 7021 10897 7055 10931
rect 7558 10897 7592 10931
rect 9137 10897 9171 10931
rect 13369 10897 13403 10931
rect 16328 10897 16362 10931
rect 18337 10897 18371 10931
rect 18598 10897 18632 10931
rect 22109 10897 22143 10931
rect 7297 10829 7331 10863
rect 8953 10829 8987 10863
rect 16589 10829 16623 10863
rect 21465 10829 21499 10863
rect 22017 10829 22051 10863
rect 22477 10829 22511 10863
rect 23121 10829 23155 10863
rect 11552 10761 11586 10795
rect 15209 10761 15243 10795
rect 6561 10693 6595 10727
rect 8677 10693 8711 10727
rect 9321 10693 9355 10727
rect 20085 10693 20119 10727
rect 6653 10489 6687 10523
rect 10609 10489 10643 10523
rect 13461 10489 13495 10523
rect 14013 10489 14047 10523
rect 16221 10489 16255 10523
rect 18337 10489 18371 10523
rect 20269 10489 20303 10523
rect 6561 10421 6595 10455
rect 7021 10421 7055 10455
rect 11345 10421 11379 10455
rect 17693 10421 17727 10455
rect 11529 10353 11563 10387
rect 18797 10353 18831 10387
rect 20913 10353 20947 10387
rect 6285 10285 6319 10319
rect 6837 10285 6871 10319
rect 7113 10285 7147 10319
rect 9229 10285 9263 10319
rect 12081 10285 12115 10319
rect 14197 10285 14231 10319
rect 14381 10285 14415 10319
rect 14565 10285 14599 10319
rect 16037 10285 16071 10319
rect 17601 10285 17635 10319
rect 17877 10285 17911 10319
rect 18061 10285 18095 10319
rect 20453 10285 20487 10319
rect 20637 10285 20671 10319
rect 21373 10285 21407 10319
rect 6377 10217 6411 10251
rect 9490 10217 9524 10251
rect 11805 10217 11839 10251
rect 12337 10208 12371 10242
rect 14289 10217 14323 10251
rect 15776 10217 15810 10251
rect 17340 10217 17374 10251
rect 17969 10217 18003 10251
rect 19058 10217 19092 10251
rect 20545 10217 20579 10251
rect 21634 10217 21668 10251
rect 14657 10149 14691 10183
rect 20177 10149 20211 10183
rect 22753 10149 22787 10183
rect 6009 9945 6043 9979
rect 6193 9945 6227 9979
rect 6745 9945 6779 9979
rect 17325 9945 17359 9979
rect 18061 9945 18095 9979
rect 21465 9945 21499 9979
rect 22477 9945 22511 9979
rect 6837 9877 6871 9911
rect 9321 9877 9355 9911
rect 15485 9877 15519 9911
rect 16206 9877 16240 9911
rect 22017 9877 22051 9911
rect 5917 9809 5951 9843
rect 6561 9809 6595 9843
rect 7021 9809 7055 9843
rect 12618 9809 12652 9843
rect 15301 9809 15335 9843
rect 15577 9809 15611 9843
rect 15669 9809 15703 9843
rect 15945 9809 15979 9843
rect 20085 9809 20119 9843
rect 20346 9809 20380 9843
rect 21833 9809 21867 9843
rect 22293 9809 22327 9843
rect 7849 9741 7883 9775
rect 10149 9741 10183 9775
rect 12357 9741 12391 9775
rect 8194 9673 8228 9707
rect 9965 9673 9999 9707
rect 10701 9673 10735 9707
rect 11736 9673 11770 9707
rect 15853 9673 15887 9707
rect 19165 9673 19199 9707
rect 21649 9673 21683 9707
rect 22109 9673 22143 9707
rect 6377 9605 6411 9639
rect 10333 9605 10367 9639
rect 12058 9605 12092 9639
rect 13737 9605 13771 9639
rect 19441 9605 19475 9639
rect 23857 11373 23891 11407
rect 24041 10897 24075 10931
rect 23765 9877 23799 9911
rect 8309 9401 8343 9435
rect 10701 9401 10735 9435
rect 11529 9401 11563 9435
rect 15025 9401 15059 9435
rect 16221 9401 16255 9435
rect 20269 9401 20303 9435
rect 21557 9401 21591 9435
rect 6469 9333 6503 9367
rect 13001 9333 13035 9367
rect 6653 9265 6687 9299
rect 9321 9265 9355 9299
rect 13185 9265 13219 9299
rect 13645 9265 13679 9299
rect 22017 9265 22051 9299
rect 22201 9265 22235 9299
rect 6929 9197 6963 9231
rect 9582 9197 9616 9231
rect 12909 9197 12943 9231
rect 16405 9197 16439 9231
rect 16773 9197 16807 9231
rect 17984 9197 18018 9231
rect 18797 9197 18831 9231
rect 20453 9197 20487 9231
rect 20637 9197 20671 9231
rect 6837 9129 6871 9163
rect 7190 9120 7224 9154
rect 12648 9129 12682 9163
rect 13369 9129 13403 9163
rect 13906 9129 13940 9163
rect 16497 9129 16531 9163
rect 16589 9129 16623 9163
rect 19058 9129 19092 9163
rect 20545 9129 20579 9163
rect 11529 9061 11563 9095
rect 16865 9061 16899 9095
rect 18337 9061 18371 9095
rect 20177 9061 20211 9095
rect 20913 9061 20947 9095
rect 22385 9061 22419 9095
rect 8125 8857 8159 8891
rect 13001 8857 13035 8891
rect 13185 8857 13219 8891
rect 14749 8857 14783 8891
rect 16865 8857 16899 8891
rect 17509 8857 17543 8891
rect 21557 8857 21591 8891
rect 7297 8789 7331 8823
rect 10517 8789 10551 8823
rect 13630 8789 13664 8823
rect 6561 8721 6595 8755
rect 6929 8721 6963 8755
rect 7389 8721 7423 8755
rect 13277 8721 13311 8755
rect 13369 8721 13403 8755
rect 15485 8721 15519 8755
rect 15746 8721 15780 8755
rect 12817 8653 12851 8687
rect 8478 8585 8512 8619
rect 11644 8585 11678 8619
rect 20085 8789 20119 8823
rect 19809 8721 19843 8755
rect 18521 8585 18555 8619
rect 19625 8585 19659 8619
rect 21212 8585 21246 8619
rect 6377 8517 6411 8551
rect 6745 8517 6779 8551
rect 7021 8517 7055 8551
rect 9505 8517 9539 8551
rect 17509 8517 17543 8551
rect 6285 8313 6319 8347
rect 8309 8313 8343 8347
rect 10701 8313 10735 8347
rect 13185 8313 13219 8347
rect 17233 8313 17267 8347
rect 20269 8313 20303 8347
rect 20913 8313 20947 8347
rect 22753 8313 22787 8347
rect 12449 8245 12483 8279
rect 11069 8177 11103 8211
rect 13737 8177 13771 8211
rect 18613 8177 18647 8211
rect 6561 8109 6595 8143
rect 6929 8109 6963 8143
rect 9321 8109 9355 8143
rect 13093 8109 13127 8143
rect 14289 8109 14323 8143
rect 15117 8109 15151 8143
rect 15301 8109 15335 8143
rect 18352 8109 18386 8143
rect 18797 8109 18831 8143
rect 19058 8109 19092 8143
rect 20453 8109 20487 8143
rect 20545 8109 20579 8143
rect 21373 8109 21407 8143
rect 6745 8041 6779 8075
rect 7185 8032 7219 8066
rect 9582 8041 9616 8075
rect 11330 8041 11364 8075
rect 14933 8041 14967 8075
rect 20637 8041 20671 8075
rect 21634 8041 21668 8075
rect 12449 7973 12483 8007
rect 13461 7973 13495 8007
rect 15117 7973 15151 8007
rect 20177 7973 20211 8007
rect 6929 7769 6963 7803
rect 9229 7769 9263 7803
rect 11253 7769 11287 7803
rect 13737 7769 13771 7803
rect 16037 7769 16071 7803
rect 21557 7769 21591 7803
rect 5549 7021 5583 7055
rect 7466 7701 7500 7735
rect 11713 7701 11747 7735
rect 12618 7701 12652 7735
rect 20085 7701 20119 7735
rect 22293 7701 22327 7735
rect 23489 7701 23523 7735
rect 6653 7633 6687 7667
rect 7205 7633 7239 7667
rect 10900 7633 10934 7667
rect 11437 7633 11471 7667
rect 11897 7633 11931 7667
rect 14105 7633 14139 7667
rect 14197 7633 14231 7667
rect 18889 7633 18923 7667
rect 5733 7429 5767 7463
rect 8861 7565 8895 7599
rect 9045 7565 9079 7599
rect 11161 7565 11195 7599
rect 12357 7565 12391 7599
rect 14381 7565 14415 7599
rect 17141 7565 17175 7599
rect 17325 7565 17359 7599
rect 22109 7565 22143 7599
rect 6469 7497 6503 7531
rect 9781 7497 9815 7531
rect 11621 7497 11655 7531
rect 14289 7497 14323 7531
rect 19901 7497 19935 7531
rect 21212 7497 21246 7531
rect 21925 7497 21959 7531
rect 6101 7429 6135 7463
rect 8585 7429 8619 7463
rect 12173 7429 12207 7463
rect 13737 7429 13771 7463
rect 6009 7225 6043 7259
rect 6377 7225 6411 7259
rect 15025 7225 15059 7259
rect 17601 7225 17635 7259
rect 17877 7225 17911 7259
rect 20637 7225 20671 7259
rect 12196 7157 12230 7191
rect 15209 7157 15243 7191
rect 18797 7157 18831 7191
rect 5917 7089 5951 7123
rect 6929 7089 6963 7123
rect 12541 7089 12575 7123
rect 16221 7089 16255 7123
rect 19257 7089 19291 7123
rect 20729 7089 20763 7123
rect 20913 7089 20947 7123
rect 21373 7089 21407 7123
rect 6193 7021 6227 7055
rect 9321 7021 9355 7055
rect 13645 7021 13679 7055
rect 15393 7021 15427 7055
rect 18061 7021 18095 7055
rect 7190 6953 7224 6987
rect 10241 6953 10275 6987
rect 11069 6953 11103 6987
rect 13906 6953 13940 6987
rect 15761 6953 15795 6987
rect 16482 6953 16516 6987
rect 18981 7021 19015 7055
rect 21189 7021 21223 7055
rect 19165 6953 19199 6987
rect 19518 6953 19552 6987
rect 21634 6953 21668 6987
rect 23857 7021 23891 7055
rect 5641 6885 5675 6919
rect 6469 6885 6503 6919
rect 6561 6885 6595 6919
rect 8309 6885 8343 6919
rect 18337 6885 18371 6919
rect 22753 6885 22787 6919
rect 6193 6681 6227 6715
rect 12081 6681 12115 6715
rect 13737 6681 13771 6715
rect 20177 6681 20211 6715
rect 22293 6681 22327 6715
rect 23673 6681 23707 6715
rect 6101 6613 6135 6647
rect 7481 6613 7515 6647
rect 7665 6613 7699 6647
rect 7849 6613 7883 6647
rect 10609 6613 10643 6647
rect 15194 6613 15228 6647
rect 6745 6545 6779 6579
rect 7021 6545 7055 6579
rect 7573 6545 7607 6579
rect 7941 6545 7975 6579
rect 8125 6553 8159 6587
rect 8478 6545 8512 6579
rect 12357 6545 12391 6579
rect 12618 6545 12652 6579
rect 14933 6545 14967 6579
rect 18337 6545 18371 6579
rect 20821 6545 20855 6579
rect 21649 6545 21683 6579
rect 21925 6545 21959 6579
rect 6377 6477 6411 6511
rect 6929 6477 6963 6511
rect 8033 6477 8067 6511
rect 8217 6477 8251 6511
rect 18613 6477 18647 6511
rect 20545 6477 20579 6511
rect 9597 6409 9631 6443
rect 11736 6409 11770 6443
rect 21005 6409 21039 6443
rect 24041 6409 24075 6443
rect 6561 6341 6595 6375
rect 7849 6341 7883 6375
rect 16313 6341 16347 6375
rect 21465 6341 21499 6375
rect 6929 6137 6963 6171
rect 7757 6137 7791 6171
rect 8217 6137 8251 6171
rect 10425 6137 10459 6171
rect 12357 6137 12391 6171
rect 13185 6137 13219 6171
rect 18061 6137 18095 6171
rect 18981 6137 19015 6171
rect 19809 6137 19843 6171
rect 21097 6137 21131 6171
rect 22385 6137 22419 6171
rect 6561 6001 6595 6035
rect 16405 6069 16439 6103
rect 20269 6069 20303 6103
rect 21557 6069 21591 6103
rect 12541 6001 12575 6035
rect 12725 6001 12759 6035
rect 12817 6001 12851 6035
rect 13369 6001 13403 6035
rect 14289 6001 14323 6035
rect 16589 6001 16623 6035
rect 19533 6001 19567 6035
rect 20453 6001 20487 6035
rect 20729 6001 20763 6035
rect 21741 6001 21775 6035
rect 21833 6001 21867 6035
rect 6745 5933 6779 5967
rect 8033 5933 8067 5967
rect 10609 5933 10643 5967
rect 13001 5933 13035 5967
rect 13277 5933 13311 5967
rect 13737 5933 13771 5967
rect 13921 5933 13955 5967
rect 14105 5933 14139 5967
rect 16865 5933 16899 5967
rect 17785 5933 17819 5967
rect 19625 5933 19659 5967
<< metal1 >>
rect 5796 21984 23000 22080
rect 18417 21947 18475 21953
rect 18417 21913 18429 21947
rect 18463 21944 18475 21947
rect 18463 21916 19104 21944
rect 18463 21913 18475 21916
rect 18417 21907 18475 21913
rect 15197 21879 15255 21885
rect 15197 21845 15209 21879
rect 15243 21876 15255 21879
rect 18969 21879 19027 21885
rect 18969 21876 18981 21879
rect 15243 21848 15792 21876
rect 15243 21845 15255 21848
rect 15197 21839 15255 21845
rect 15105 21811 15163 21817
rect 15105 21777 15117 21811
rect 15151 21808 15163 21811
rect 15657 21811 15715 21817
rect 15657 21808 15669 21811
rect 15151 21780 15669 21808
rect 15151 21777 15163 21780
rect 15105 21771 15163 21777
rect 15657 21777 15669 21780
rect 15703 21777 15715 21811
rect 15764 21808 15792 21848
rect 18432 21848 18981 21876
rect 15841 21811 15899 21817
rect 15841 21808 15853 21811
rect 15764 21780 15853 21808
rect 15657 21771 15715 21777
rect 15841 21777 15853 21780
rect 15887 21808 15899 21811
rect 15930 21808 15936 21820
rect 15887 21780 15936 21808
rect 15887 21777 15899 21780
rect 15841 21771 15899 21777
rect 15930 21768 15936 21780
rect 15988 21768 15994 21820
rect 16684 21780 17540 21808
rect 10318 21740 10324 21752
rect 10263 21712 10324 21740
rect 10318 21700 10324 21712
rect 10376 21700 10382 21752
rect 14274 21700 14280 21752
rect 14332 21740 14338 21752
rect 15013 21743 15071 21749
rect 15013 21740 15025 21743
rect 14332 21712 15025 21740
rect 14332 21700 14338 21712
rect 15013 21709 15025 21712
rect 15059 21709 15071 21743
rect 15013 21703 15071 21709
rect 16482 21700 16488 21752
rect 16540 21740 16546 21752
rect 16684 21740 16712 21780
rect 16540 21712 16712 21740
rect 17512 21740 17540 21780
rect 18230 21768 18236 21820
rect 18288 21808 18294 21820
rect 18325 21811 18383 21817
rect 18325 21808 18337 21811
rect 18288 21780 18337 21808
rect 18288 21768 18294 21780
rect 18325 21777 18337 21780
rect 18371 21808 18383 21811
rect 18432 21808 18460 21848
rect 18969 21845 18981 21848
rect 19015 21845 19027 21879
rect 19076 21876 19104 21916
rect 19153 21879 19211 21885
rect 19153 21876 19165 21879
rect 19076 21848 19165 21876
rect 18969 21839 19027 21845
rect 19153 21845 19165 21848
rect 19199 21876 19211 21879
rect 20732 21882 21404 21910
rect 20732 21876 20760 21882
rect 19199 21848 20760 21876
rect 21376 21876 21404 21882
rect 21376 21848 21864 21876
rect 19199 21845 19211 21848
rect 19153 21839 19211 21845
rect 20548 21817 20576 21848
rect 18371 21780 18460 21808
rect 20257 21811 20315 21817
rect 18371 21777 18383 21780
rect 18325 21771 18383 21777
rect 20257 21777 20269 21811
rect 20303 21777 20315 21811
rect 20257 21771 20315 21777
rect 20533 21811 20591 21817
rect 20533 21777 20545 21811
rect 20579 21777 20591 21811
rect 20533 21771 20591 21777
rect 20993 21811 21051 21817
rect 20993 21777 21005 21811
rect 21039 21808 21051 21811
rect 21266 21808 21272 21820
rect 21039 21780 21272 21808
rect 21039 21777 21051 21780
rect 20993 21771 21051 21777
rect 19610 21740 19616 21752
rect 17512 21712 19616 21740
rect 16540 21700 16546 21712
rect 19610 21700 19616 21712
rect 19668 21740 19674 21752
rect 19705 21743 19763 21749
rect 19705 21740 19717 21743
rect 19668 21712 19717 21740
rect 19668 21700 19674 21712
rect 19705 21709 19717 21712
rect 19751 21709 19763 21743
rect 19705 21703 19763 21709
rect 10134 21672 10140 21684
rect 10079 21644 10140 21672
rect 10134 21632 10140 21644
rect 10192 21632 10198 21684
rect 15856 21644 16344 21672
rect 10502 21604 10508 21616
rect 10447 21576 10508 21604
rect 10502 21564 10508 21576
rect 10560 21564 10566 21616
rect 15381 21607 15439 21613
rect 15381 21573 15393 21607
rect 15427 21604 15439 21607
rect 15470 21604 15476 21616
rect 15427 21576 15476 21604
rect 15427 21573 15439 21576
rect 15381 21567 15439 21573
rect 15470 21564 15476 21576
rect 15528 21564 15534 21616
rect 15657 21607 15715 21613
rect 15657 21573 15669 21607
rect 15703 21604 15715 21607
rect 15856 21604 15884 21644
rect 16316 21638 16344 21644
rect 16316 21610 17264 21638
rect 18414 21632 18420 21684
rect 18472 21672 18478 21684
rect 18601 21675 18659 21681
rect 18601 21672 18613 21675
rect 18472 21644 18613 21672
rect 18472 21632 18478 21644
rect 18601 21641 18613 21644
rect 18647 21641 18659 21675
rect 18601 21635 18659 21641
rect 19521 21675 19579 21681
rect 19521 21641 19533 21675
rect 19567 21672 19579 21675
rect 20073 21675 20131 21681
rect 20073 21672 20085 21675
rect 19567 21644 20085 21672
rect 19567 21641 19579 21644
rect 19521 21635 19579 21641
rect 20073 21641 20085 21644
rect 20119 21641 20131 21675
rect 20272 21672 20300 21771
rect 21266 21768 21272 21780
rect 21324 21768 21330 21820
rect 21836 21808 21864 21848
rect 22649 21811 22707 21817
rect 22649 21808 22661 21811
rect 21836 21780 22661 21808
rect 22649 21777 22661 21780
rect 22695 21777 22707 21811
rect 22649 21771 22707 21777
rect 22738 21768 22744 21820
rect 22796 21808 22802 21820
rect 22833 21811 22891 21817
rect 22833 21808 22845 21811
rect 22796 21780 22845 21808
rect 22796 21768 22802 21780
rect 22833 21777 22845 21780
rect 22879 21777 22891 21811
rect 22833 21771 22891 21777
rect 20346 21700 20352 21752
rect 20404 21740 20410 21752
rect 20441 21743 20499 21749
rect 20441 21740 20453 21743
rect 20404 21712 20453 21740
rect 20404 21700 20410 21712
rect 20441 21709 20453 21712
rect 20487 21709 20499 21743
rect 20901 21743 20959 21749
rect 20901 21740 20913 21743
rect 20441 21703 20499 21709
rect 20548 21712 20913 21740
rect 20548 21672 20576 21712
rect 20901 21709 20913 21712
rect 20947 21709 20959 21743
rect 20901 21703 20959 21709
rect 20272 21644 20576 21672
rect 20916 21672 20944 21703
rect 21082 21700 21088 21752
rect 21140 21740 21146 21752
rect 21729 21743 21787 21749
rect 21729 21740 21741 21743
rect 21140 21712 21741 21740
rect 21140 21700 21146 21712
rect 21729 21709 21741 21712
rect 21775 21709 21787 21743
rect 22002 21740 22008 21752
rect 21947 21712 22008 21740
rect 21729 21703 21787 21709
rect 22002 21700 22008 21712
rect 22060 21700 22066 21752
rect 22741 21675 22799 21681
rect 22741 21672 22753 21675
rect 20916 21644 22753 21672
rect 20073 21635 20131 21641
rect 22741 21641 22753 21644
rect 22787 21641 22799 21675
rect 22741 21635 22799 21641
rect 15703 21576 15884 21604
rect 17236 21604 17264 21610
rect 17402 21604 17408 21616
rect 17236 21576 17408 21604
rect 15703 21573 15715 21576
rect 15657 21567 15715 21573
rect 17402 21564 17408 21576
rect 17460 21564 17466 21616
rect 19150 21604 19156 21616
rect 19095 21576 19156 21604
rect 19150 21564 19156 21576
rect 19208 21564 19214 21616
rect 19886 21604 19892 21616
rect 19831 21576 19892 21604
rect 19886 21564 19892 21576
rect 19944 21564 19950 21616
rect 19978 21564 19984 21616
rect 20036 21604 20042 21616
rect 20717 21607 20775 21613
rect 20717 21604 20729 21607
rect 20036 21576 20729 21604
rect 20036 21564 20042 21576
rect 20717 21573 20729 21576
rect 20763 21573 20775 21607
rect 20717 21567 20775 21573
rect 21545 21607 21603 21613
rect 21545 21573 21557 21607
rect 21591 21604 21603 21607
rect 21634 21604 21640 21616
rect 21591 21576 21640 21604
rect 21591 21573 21603 21576
rect 21545 21567 21603 21573
rect 21634 21564 21640 21576
rect 21692 21564 21698 21616
rect 22370 21604 22376 21616
rect 22315 21576 22376 21604
rect 22370 21564 22376 21576
rect 22428 21564 22434 21616
rect 5796 21440 23000 21536
rect 10134 21400 10140 21412
rect 10079 21372 10140 21400
rect 10134 21360 10140 21372
rect 10192 21360 10198 21412
rect 15930 21400 15936 21412
rect 15875 21372 15936 21400
rect 15930 21360 15936 21372
rect 15988 21360 15994 21412
rect 17313 21403 17371 21409
rect 17313 21400 17325 21403
rect 17144 21372 17325 21400
rect 17144 21344 17172 21372
rect 17313 21369 17325 21372
rect 17359 21400 17371 21403
rect 17681 21403 17739 21409
rect 17681 21400 17693 21403
rect 17359 21372 17693 21400
rect 17359 21369 17371 21372
rect 17313 21363 17371 21369
rect 17681 21369 17693 21372
rect 17727 21369 17739 21403
rect 17681 21363 17739 21369
rect 18141 21403 18199 21409
rect 18141 21369 18153 21403
rect 18187 21400 18199 21403
rect 18230 21400 18236 21412
rect 18187 21372 18236 21400
rect 18187 21369 18199 21372
rect 18141 21363 18199 21369
rect 18230 21360 18236 21372
rect 18288 21360 18294 21412
rect 19978 21400 19984 21412
rect 19812 21372 19984 21400
rect 17126 21292 17132 21344
rect 17184 21292 17190 21344
rect 19150 21292 19156 21344
rect 19208 21332 19214 21344
rect 19245 21335 19303 21341
rect 19245 21332 19257 21335
rect 19208 21304 19257 21332
rect 19208 21292 19214 21304
rect 19245 21301 19257 21304
rect 19291 21301 19303 21335
rect 19245 21295 19303 21301
rect 19705 21335 19763 21341
rect 19705 21301 19717 21335
rect 19751 21332 19763 21335
rect 19812 21332 19840 21372
rect 19978 21360 19984 21372
rect 20036 21360 20042 21412
rect 21453 21403 21511 21409
rect 21453 21369 21465 21403
rect 21499 21400 21511 21403
rect 22002 21400 22008 21412
rect 21499 21372 22008 21400
rect 21499 21369 21511 21372
rect 21453 21363 21511 21369
rect 22002 21360 22008 21372
rect 22060 21360 22066 21412
rect 19751 21304 19840 21332
rect 19751 21301 19763 21304
rect 19705 21295 19763 21301
rect 22186 21292 22192 21344
rect 22244 21332 22250 21344
rect 22480 21335 22538 21341
rect 22480 21332 22492 21335
rect 22244 21304 22492 21332
rect 22244 21292 22250 21304
rect 22480 21301 22492 21304
rect 22526 21301 22538 21335
rect 22480 21295 22538 21301
rect 14001 21267 14059 21273
rect 14001 21264 14013 21267
rect 13372 21236 14013 21264
rect 13372 21208 13400 21236
rect 14001 21233 14013 21236
rect 14047 21233 14059 21267
rect 16393 21267 16451 21273
rect 16393 21264 16405 21267
rect 14001 21227 14059 21233
rect 15672 21236 16405 21264
rect 10962 21156 10968 21208
rect 11020 21196 11026 21208
rect 12989 21199 13047 21205
rect 12989 21196 13001 21199
rect 11020 21168 13001 21196
rect 11020 21156 11026 21168
rect 12989 21165 13001 21168
rect 13035 21196 13047 21199
rect 13078 21196 13084 21208
rect 13035 21168 13084 21196
rect 13035 21165 13047 21168
rect 12989 21159 13047 21165
rect 13078 21156 13084 21168
rect 13136 21156 13142 21208
rect 13354 21156 13360 21208
rect 13412 21156 13418 21208
rect 13817 21199 13875 21205
rect 13817 21165 13829 21199
rect 13863 21165 13875 21199
rect 13817 21159 13875 21165
rect 14093 21199 14151 21205
rect 14093 21165 14105 21199
rect 14139 21196 14151 21199
rect 14458 21196 14464 21208
rect 14139 21168 14464 21196
rect 14139 21165 14151 21168
rect 14093 21159 14151 21165
rect 13832 21128 13860 21159
rect 14458 21156 14464 21168
rect 14516 21156 14522 21208
rect 15102 21156 15108 21208
rect 15160 21196 15166 21208
rect 15672 21196 15700 21236
rect 16393 21233 16405 21236
rect 16439 21264 16451 21267
rect 16482 21264 16488 21276
rect 16439 21236 16488 21264
rect 16439 21233 16451 21236
rect 16393 21227 16451 21233
rect 16482 21224 16488 21236
rect 16540 21224 16546 21276
rect 17402 21264 17408 21276
rect 17347 21236 17408 21264
rect 17402 21224 17408 21236
rect 17460 21264 17466 21276
rect 19061 21267 19119 21273
rect 17460 21236 18000 21264
rect 17460 21224 17466 21236
rect 15160 21168 15700 21196
rect 15749 21199 15807 21205
rect 15160 21156 15166 21168
rect 15749 21165 15761 21199
rect 15795 21196 15807 21199
rect 15930 21196 15936 21208
rect 15795 21168 15936 21196
rect 15795 21165 15807 21168
rect 15749 21159 15807 21165
rect 15930 21156 15936 21168
rect 15988 21156 15994 21208
rect 17972 21205 18000 21236
rect 19061 21233 19073 21267
rect 19107 21264 19119 21267
rect 19521 21267 19579 21273
rect 19521 21264 19533 21267
rect 19107 21236 19533 21264
rect 19107 21233 19119 21236
rect 19061 21227 19119 21233
rect 19521 21233 19533 21236
rect 19567 21264 19579 21267
rect 19610 21264 19616 21276
rect 19567 21236 19616 21264
rect 19567 21233 19579 21236
rect 19521 21227 19579 21233
rect 19610 21224 19616 21236
rect 19668 21224 19674 21276
rect 21450 21224 21456 21276
rect 21508 21264 21514 21276
rect 21508 21236 21758 21264
rect 21508 21224 21514 21236
rect 17129 21199 17187 21205
rect 17129 21165 17141 21199
rect 17175 21196 17187 21199
rect 17957 21199 18015 21205
rect 17175 21168 17356 21196
rect 17175 21165 17187 21168
rect 17129 21159 17187 21165
rect 14274 21128 14280 21140
rect 13832 21100 14280 21128
rect 14274 21088 14280 21100
rect 14332 21088 14338 21140
rect 15488 21131 15546 21137
rect 15488 21097 15500 21131
rect 15534 21128 15546 21131
rect 16114 21128 16120 21140
rect 15534 21100 16120 21128
rect 15534 21097 15546 21100
rect 15488 21091 15546 21097
rect 16114 21088 16120 21100
rect 16172 21088 16178 21140
rect 17328 21128 17356 21168
rect 17957 21165 17969 21199
rect 18003 21165 18015 21199
rect 17957 21159 18015 21165
rect 19797 21199 19855 21205
rect 19797 21165 19809 21199
rect 19843 21196 19855 21199
rect 20070 21196 20076 21208
rect 19843 21168 20076 21196
rect 19843 21165 19855 21168
rect 19797 21159 19855 21165
rect 20070 21156 20076 21168
rect 20128 21156 20134 21208
rect 21266 21156 21272 21208
rect 21324 21196 21330 21208
rect 21324 21168 21666 21196
rect 21324 21156 21330 21168
rect 17865 21131 17923 21137
rect 17865 21128 17877 21131
rect 17328 21100 17877 21128
rect 17865 21097 17877 21100
rect 17911 21128 17923 21131
rect 18414 21128 18420 21140
rect 17911 21100 18420 21128
rect 17911 21097 17923 21100
rect 17865 21091 17923 21097
rect 18414 21088 18420 21100
rect 18472 21088 18478 21140
rect 19996 21122 20111 21128
rect 19996 21100 20065 21122
rect 9950 21020 9956 21072
rect 10008 21060 10014 21072
rect 10045 21063 10103 21069
rect 10045 21060 10057 21063
rect 10008 21032 10057 21060
rect 10008 21020 10014 21032
rect 10045 21029 10057 21032
rect 10091 21029 10103 21063
rect 10045 21023 10103 21029
rect 12618 21020 12624 21072
rect 12676 21060 12682 21072
rect 12805 21063 12863 21069
rect 12805 21060 12817 21063
rect 12676 21032 12817 21060
rect 12676 21020 12682 21032
rect 12805 21029 12817 21032
rect 12851 21029 12863 21063
rect 14366 21060 14372 21072
rect 14311 21032 14372 21060
rect 12805 21023 12863 21029
rect 14366 21020 14372 21032
rect 14424 21020 14430 21072
rect 14734 21020 14740 21072
rect 14792 21060 14798 21072
rect 15841 21063 15899 21069
rect 15841 21060 15853 21063
rect 14792 21032 15853 21060
rect 14792 21020 14798 21032
rect 15841 21029 15853 21032
rect 15887 21029 15899 21063
rect 16206 21060 16212 21072
rect 16151 21032 16212 21060
rect 15841 21023 15899 21029
rect 16206 21020 16212 21032
rect 16264 21020 16270 21072
rect 17678 21020 17684 21072
rect 17736 21060 17742 21072
rect 18049 21063 18107 21069
rect 18049 21060 18061 21063
rect 17736 21032 18061 21060
rect 17736 21020 17742 21032
rect 18049 21029 18061 21032
rect 18095 21029 18107 21063
rect 18874 21060 18880 21072
rect 18819 21032 18880 21060
rect 18049 21023 18107 21029
rect 18874 21020 18880 21032
rect 18932 21020 18938 21072
rect 19337 21063 19395 21069
rect 19337 21029 19349 21063
rect 19383 21060 19395 21063
rect 19996 21060 20024 21100
rect 20053 21088 20065 21100
rect 20099 21088 20111 21122
rect 20053 21082 20111 21088
rect 19383 21032 20024 21060
rect 19383 21029 19395 21032
rect 19337 21023 19395 21029
rect 5796 20896 23000 20992
rect 10885 20816 10891 20868
rect 10943 20816 10949 20868
rect 10885 20801 10949 20816
rect 10885 20767 10900 20801
rect 10934 20767 10949 20801
rect 10885 20761 10949 20767
rect 12603 20816 12609 20868
rect 12661 20816 12667 20868
rect 14274 20856 14280 20868
rect 14219 20828 14280 20856
rect 14274 20816 14280 20828
rect 14332 20816 14338 20868
rect 15381 20859 15439 20865
rect 15381 20825 15393 20859
rect 15427 20856 15439 20859
rect 15470 20856 15476 20868
rect 15427 20828 15476 20856
rect 15427 20825 15439 20828
rect 15381 20819 15439 20825
rect 15470 20816 15476 20828
rect 15528 20816 15534 20868
rect 20438 20816 20444 20868
rect 20496 20856 20502 20868
rect 21453 20859 21511 20865
rect 21453 20856 21465 20859
rect 20496 20828 20668 20856
rect 20496 20816 20502 20828
rect 12603 20801 12667 20816
rect 12603 20767 12618 20801
rect 12652 20767 12667 20801
rect 12603 20761 12667 20767
rect 13078 20748 13084 20800
rect 13136 20788 13142 20800
rect 16206 20797 16212 20800
rect 16194 20791 16212 20797
rect 16194 20788 16206 20791
rect 13136 20760 14688 20788
rect 16151 20760 16206 20788
rect 13136 20748 13142 20760
rect 7558 20729 7564 20732
rect 7546 20723 7564 20729
rect 7546 20720 7558 20723
rect 7503 20692 7558 20720
rect 7546 20689 7558 20692
rect 7546 20683 7564 20689
rect 7558 20680 7564 20683
rect 7616 20680 7622 20732
rect 10870 20680 10876 20732
rect 10928 20720 10934 20732
rect 11149 20723 11207 20729
rect 11149 20720 11161 20723
rect 10928 20692 11161 20720
rect 10928 20680 10934 20692
rect 11149 20689 11161 20692
rect 11195 20689 11207 20723
rect 11149 20683 11207 20689
rect 12345 20723 12403 20729
rect 12345 20689 12357 20723
rect 12391 20720 12403 20723
rect 12618 20720 12624 20732
rect 12391 20692 12624 20720
rect 12391 20689 12403 20692
rect 12345 20683 12403 20689
rect 12618 20680 12624 20692
rect 12676 20680 12682 20732
rect 14553 20723 14611 20729
rect 14553 20689 14565 20723
rect 14599 20689 14611 20723
rect 14660 20720 14688 20760
rect 16194 20757 16206 20760
rect 16194 20751 16212 20757
rect 16206 20748 16212 20751
rect 16264 20748 16270 20800
rect 18874 20788 18880 20800
rect 18932 20797 18938 20800
rect 18932 20791 18950 20797
rect 18831 20760 18880 20788
rect 18874 20748 18880 20760
rect 18938 20757 18950 20791
rect 18932 20751 18950 20757
rect 18932 20748 18938 20751
rect 19886 20748 19892 20800
rect 19944 20788 19950 20800
rect 20334 20791 20392 20797
rect 20334 20788 20346 20791
rect 19944 20760 20346 20788
rect 19944 20748 19950 20760
rect 20334 20757 20346 20760
rect 20380 20757 20392 20791
rect 20640 20788 20668 20828
rect 21284 20828 21465 20856
rect 21284 20788 21312 20828
rect 21453 20825 21465 20828
rect 21499 20825 21511 20859
rect 21453 20819 21511 20825
rect 20640 20760 21312 20788
rect 20334 20751 20392 20757
rect 15102 20720 15108 20732
rect 14660 20692 15108 20720
rect 14553 20683 14611 20689
rect 7282 20652 7288 20664
rect 7227 20624 7288 20652
rect 7282 20612 7288 20624
rect 7340 20612 7346 20664
rect 14277 20655 14335 20661
rect 14277 20652 14289 20655
rect 13372 20624 14289 20652
rect 11514 20544 11520 20596
rect 11572 20584 11578 20596
rect 13372 20584 13400 20624
rect 14277 20621 14289 20624
rect 14323 20652 14335 20655
rect 14458 20652 14464 20664
rect 14323 20624 14464 20652
rect 14323 20621 14335 20624
rect 14277 20615 14335 20621
rect 14458 20612 14464 20624
rect 14516 20612 14522 20664
rect 11572 20556 12020 20584
rect 11572 20544 11578 20556
rect 8665 20519 8723 20525
rect 8665 20485 8677 20519
rect 8711 20516 8723 20519
rect 9122 20516 9128 20528
rect 8711 20488 9128 20516
rect 8711 20485 8723 20488
rect 8665 20479 8723 20485
rect 9122 20476 9128 20488
rect 9180 20476 9186 20528
rect 9769 20519 9827 20525
rect 9769 20485 9781 20519
rect 9815 20516 9827 20519
rect 9950 20516 9956 20528
rect 9815 20488 9956 20516
rect 9815 20485 9827 20488
rect 9769 20479 9827 20485
rect 9950 20476 9956 20488
rect 10008 20476 10014 20528
rect 11992 20516 12020 20556
rect 13280 20556 13400 20584
rect 13280 20516 13308 20556
rect 11992 20488 13308 20516
rect 13354 20476 13360 20528
rect 13412 20516 13418 20528
rect 13725 20519 13783 20525
rect 13725 20516 13737 20519
rect 13412 20488 13737 20516
rect 13412 20476 13418 20488
rect 13725 20485 13737 20488
rect 13771 20516 13783 20519
rect 14568 20516 14596 20683
rect 15102 20680 15108 20692
rect 15160 20680 15166 20732
rect 21913 20723 21971 20729
rect 21913 20689 21925 20723
rect 21959 20720 21971 20723
rect 22554 20720 22560 20732
rect 21959 20692 22560 20720
rect 21959 20689 21971 20692
rect 21913 20683 21971 20689
rect 22554 20680 22560 20692
rect 22612 20680 22618 20732
rect 15930 20652 15936 20664
rect 15875 20624 15936 20652
rect 15930 20612 15936 20624
rect 15988 20612 15994 20664
rect 19150 20652 19156 20664
rect 19095 20624 19156 20652
rect 19150 20612 19156 20624
rect 19208 20612 19214 20664
rect 20070 20652 20076 20664
rect 20015 20624 20076 20652
rect 20070 20612 20076 20624
rect 20128 20612 20134 20664
rect 21729 20655 21787 20661
rect 21729 20621 21741 20655
rect 21775 20652 21787 20655
rect 22002 20652 22008 20664
rect 21775 20624 22008 20652
rect 21775 20621 21787 20624
rect 21729 20615 21787 20621
rect 22002 20612 22008 20624
rect 22060 20612 22066 20664
rect 21545 20587 21603 20593
rect 21545 20553 21557 20587
rect 21591 20584 21603 20587
rect 23109 20587 23167 20593
rect 23109 20584 23121 20587
rect 21591 20556 23121 20584
rect 21591 20553 21603 20556
rect 21545 20547 21603 20553
rect 23109 20553 23121 20556
rect 23155 20553 23167 20587
rect 23109 20547 23167 20553
rect 13771 20488 14596 20516
rect 14921 20519 14979 20525
rect 13771 20485 13783 20488
rect 13725 20479 13783 20485
rect 14921 20485 14933 20519
rect 14967 20516 14979 20519
rect 15470 20516 15476 20528
rect 14967 20488 15476 20516
rect 14967 20485 14979 20488
rect 14921 20479 14979 20485
rect 15470 20476 15476 20488
rect 15528 20476 15534 20528
rect 17126 20476 17132 20528
rect 17184 20516 17190 20528
rect 17313 20519 17371 20525
rect 17313 20516 17325 20519
rect 17184 20488 17325 20516
rect 17184 20476 17190 20488
rect 17313 20485 17325 20488
rect 17359 20485 17371 20519
rect 17313 20479 17371 20485
rect 17678 20476 17684 20528
rect 17736 20516 17742 20528
rect 17773 20519 17831 20525
rect 17773 20516 17785 20519
rect 17736 20488 17785 20516
rect 17736 20476 17742 20488
rect 17773 20485 17785 20488
rect 17819 20485 17831 20519
rect 17773 20479 17831 20485
rect 5796 20352 23000 20448
rect 10318 20272 10324 20324
rect 10376 20312 10382 20324
rect 11057 20315 11115 20321
rect 11057 20312 11069 20315
rect 10376 20284 11069 20312
rect 10376 20272 10382 20284
rect 11057 20281 11069 20284
rect 11103 20281 11115 20315
rect 11057 20275 11115 20281
rect 6822 20176 6828 20188
rect 6767 20148 6828 20176
rect 6822 20136 6828 20148
rect 6880 20136 6886 20188
rect 10505 20179 10563 20185
rect 10505 20145 10517 20179
rect 10551 20176 10563 20179
rect 10686 20176 10692 20188
rect 10551 20148 10692 20176
rect 10551 20145 10563 20148
rect 10505 20139 10563 20145
rect 10686 20136 10692 20148
rect 10744 20136 10750 20188
rect 22922 20176 22928 20188
rect 22867 20148 22928 20176
rect 22922 20136 22928 20148
rect 22980 20136 22986 20188
rect 12437 20111 12495 20117
rect 12437 20077 12449 20111
rect 12483 20108 12495 20111
rect 12618 20108 12624 20120
rect 12483 20080 12624 20108
rect 12483 20077 12495 20080
rect 12437 20071 12495 20077
rect 12618 20068 12624 20080
rect 12676 20108 12682 20120
rect 15565 20111 15623 20117
rect 15565 20108 15577 20111
rect 12676 20080 15577 20108
rect 12676 20068 12682 20080
rect 15565 20077 15577 20080
rect 15611 20108 15623 20111
rect 15930 20108 15936 20120
rect 15611 20080 15936 20108
rect 15611 20077 15623 20080
rect 15565 20071 15623 20077
rect 15930 20068 15936 20080
rect 15988 20108 15994 20120
rect 16209 20111 16267 20117
rect 16209 20108 16221 20111
rect 15988 20080 16221 20108
rect 15988 20068 15994 20080
rect 16209 20077 16221 20080
rect 16255 20077 16267 20111
rect 16209 20071 16267 20077
rect 20070 20068 20076 20120
rect 20128 20108 20134 20120
rect 20165 20111 20223 20117
rect 20165 20108 20177 20111
rect 20128 20080 20177 20108
rect 20128 20068 20134 20080
rect 20165 20077 20177 20080
rect 20211 20077 20223 20111
rect 20165 20071 20223 20077
rect 20364 20080 21404 20108
rect 6914 20000 6920 20052
rect 6972 20040 6978 20052
rect 7086 20043 7144 20049
rect 7086 20040 7098 20043
rect 6972 20012 7098 20040
rect 6972 20000 6978 20012
rect 7086 20009 7098 20012
rect 7132 20009 7144 20043
rect 10226 20040 10232 20052
rect 10284 20049 10290 20052
rect 10284 20043 10302 20049
rect 7086 20003 7144 20009
rect 7300 20012 8064 20040
rect 10183 20012 10232 20040
rect 6730 19932 6736 19984
rect 6788 19972 6794 19984
rect 7300 19972 7328 20012
rect 6788 19944 7328 19972
rect 8036 19972 8064 20012
rect 10226 20000 10232 20012
rect 10290 20009 10302 20043
rect 10284 20003 10302 20009
rect 12176 20043 12234 20049
rect 12176 20009 12188 20043
rect 12222 20040 12234 20043
rect 12342 20040 12348 20052
rect 12222 20012 12348 20040
rect 12222 20009 12234 20012
rect 12176 20003 12234 20009
rect 10284 20000 10290 20003
rect 12342 20000 12348 20012
rect 12400 20000 12406 20052
rect 15304 20043 15362 20049
rect 15304 20009 15316 20043
rect 15350 20040 15362 20043
rect 15470 20040 15476 20052
rect 15350 20012 15476 20040
rect 15350 20009 15362 20012
rect 15304 20003 15362 20009
rect 15470 20000 15476 20012
rect 15528 20000 15534 20052
rect 16298 20000 16304 20052
rect 16356 20040 16362 20052
rect 16470 20043 16528 20049
rect 16470 20040 16482 20043
rect 16356 20012 16482 20040
rect 16356 20000 16362 20012
rect 16470 20009 16482 20012
rect 16516 20009 16528 20043
rect 16470 20003 16528 20009
rect 16684 20012 17448 20040
rect 8205 19975 8263 19981
rect 8205 19972 8217 19975
rect 8036 19944 8217 19972
rect 6788 19932 6794 19944
rect 8205 19941 8217 19944
rect 8251 19972 8263 19975
rect 8754 19972 8760 19984
rect 8251 19944 8760 19972
rect 8251 19941 8263 19944
rect 8205 19935 8263 19941
rect 8754 19932 8760 19944
rect 8812 19932 8818 19984
rect 8938 19932 8944 19984
rect 8996 19972 9002 19984
rect 9125 19975 9183 19981
rect 9125 19972 9137 19975
rect 8996 19944 9137 19972
rect 8996 19932 9002 19944
rect 9125 19941 9137 19944
rect 9171 19941 9183 19975
rect 9125 19935 9183 19941
rect 13446 19932 13452 19984
rect 13504 19972 13510 19984
rect 14185 19975 14243 19981
rect 14185 19972 14197 19975
rect 13504 19944 14197 19972
rect 13504 19932 13510 19944
rect 14185 19941 14197 19944
rect 14231 19972 14243 19975
rect 14734 19972 14740 19984
rect 14231 19944 14740 19972
rect 14231 19941 14243 19944
rect 14185 19935 14243 19941
rect 14734 19932 14740 19944
rect 14792 19932 14798 19984
rect 16022 19932 16028 19984
rect 16080 19972 16086 19984
rect 16684 19972 16712 20012
rect 16080 19944 16712 19972
rect 17420 19972 17448 20012
rect 18064 20012 18644 20040
rect 17589 19975 17647 19981
rect 17589 19972 17601 19975
rect 17420 19944 17601 19972
rect 16080 19932 16086 19944
rect 17589 19941 17601 19944
rect 17635 19941 17647 19975
rect 17589 19935 17647 19941
rect 17862 19932 17868 19984
rect 17920 19972 17926 19984
rect 18064 19972 18092 20012
rect 17920 19944 18092 19972
rect 18616 19972 18644 20012
rect 18874 20000 18880 20052
rect 18932 20040 18938 20052
rect 19904 20043 19962 20049
rect 19904 20040 19916 20043
rect 18932 20012 19916 20040
rect 18932 20000 18938 20012
rect 19904 20009 19916 20012
rect 19950 20009 19962 20043
rect 19904 20003 19962 20009
rect 18785 19975 18843 19981
rect 18785 19972 18797 19975
rect 18616 19944 18797 19972
rect 17920 19932 17926 19944
rect 18785 19941 18797 19944
rect 18831 19941 18843 19975
rect 18785 19935 18843 19941
rect 20162 19932 20168 19984
rect 20220 19972 20226 19984
rect 20364 19972 20392 20080
rect 20220 19944 20392 19972
rect 21376 19972 21404 20080
rect 22664 20043 22722 20049
rect 22664 20009 22676 20043
rect 22710 20040 22722 20043
rect 22922 20040 22928 20052
rect 22710 20012 22928 20040
rect 22710 20009 22722 20012
rect 22664 20003 22722 20009
rect 22922 20000 22928 20012
rect 22980 20000 22986 20052
rect 21545 19975 21603 19981
rect 21545 19972 21557 19975
rect 21376 19944 21557 19972
rect 20220 19932 20226 19944
rect 21545 19941 21557 19944
rect 21591 19941 21603 19975
rect 21545 19935 21603 19941
rect 5796 19808 23000 19904
rect 7558 19728 7564 19780
rect 7616 19768 7622 19780
rect 7837 19771 7895 19777
rect 7837 19768 7849 19771
rect 7616 19740 7849 19768
rect 7616 19728 7622 19740
rect 7837 19737 7849 19740
rect 7883 19737 7895 19771
rect 7837 19731 7895 19737
rect 8849 19771 8907 19777
rect 8849 19737 8861 19771
rect 8895 19768 8907 19771
rect 8938 19768 8944 19780
rect 8895 19740 8944 19768
rect 8895 19737 8907 19740
rect 8849 19731 8907 19737
rect 8938 19728 8944 19740
rect 8996 19728 9002 19780
rect 9122 19768 9128 19780
rect 9067 19740 9128 19768
rect 9122 19728 9128 19740
rect 9180 19728 9186 19780
rect 10226 19728 10232 19780
rect 10284 19768 10290 19780
rect 10321 19771 10379 19777
rect 10321 19768 10333 19771
rect 10284 19740 10333 19768
rect 10284 19728 10290 19740
rect 10321 19737 10333 19740
rect 10367 19737 10379 19771
rect 10321 19731 10379 19737
rect 15473 19771 15531 19777
rect 15473 19737 15485 19771
rect 15519 19768 15531 19771
rect 16114 19768 16120 19780
rect 15519 19740 16120 19768
rect 15519 19737 15531 19740
rect 15473 19731 15531 19737
rect 16114 19728 16120 19740
rect 16172 19728 16178 19780
rect 16298 19768 16304 19780
rect 16243 19740 16304 19768
rect 16298 19728 16304 19740
rect 16356 19728 16362 19780
rect 16761 19771 16819 19777
rect 16761 19737 16773 19771
rect 16807 19768 16819 19771
rect 18874 19768 18880 19780
rect 16807 19740 16988 19768
rect 16807 19737 16819 19740
rect 16761 19731 16819 19737
rect 16960 19734 16988 19740
rect 17880 19740 18880 19768
rect 17880 19734 17908 19740
rect 8754 19660 8760 19712
rect 8812 19700 8818 19712
rect 9033 19703 9091 19709
rect 9033 19700 9045 19703
rect 8812 19672 9045 19700
rect 8812 19660 8818 19672
rect 9033 19669 9045 19672
rect 9079 19669 9091 19703
rect 9033 19663 9091 19669
rect 12713 19703 12771 19709
rect 12713 19669 12725 19703
rect 12759 19700 12771 19703
rect 13066 19703 13124 19709
rect 16960 19706 17908 19734
rect 18874 19728 18880 19740
rect 18932 19728 18938 19780
rect 21085 19771 21143 19777
rect 21085 19737 21097 19771
rect 21131 19768 21143 19771
rect 22002 19768 22008 19780
rect 21131 19740 21312 19768
rect 21131 19737 21143 19740
rect 21085 19731 21143 19737
rect 13066 19700 13078 19703
rect 12759 19672 13078 19700
rect 12759 19669 12771 19672
rect 12713 19663 12771 19669
rect 13066 19669 13078 19672
rect 13112 19669 13124 19703
rect 21284 19700 21312 19740
rect 21836 19740 22008 19768
rect 21836 19700 21864 19740
rect 22002 19728 22008 19740
rect 22060 19728 22066 19780
rect 13066 19663 13124 19669
rect 13280 19672 15056 19700
rect 21284 19672 21864 19700
rect 22204 19703 22262 19709
rect 7006 19592 7012 19644
rect 7064 19632 7070 19644
rect 8021 19635 8079 19641
rect 8021 19632 8033 19635
rect 7064 19604 8033 19632
rect 7064 19592 7070 19604
rect 8021 19601 8033 19604
rect 8067 19632 8079 19635
rect 10502 19632 10508 19644
rect 8067 19604 10508 19632
rect 8067 19601 8079 19604
rect 8021 19595 8079 19601
rect 10502 19592 10508 19604
rect 10560 19592 10566 19644
rect 11977 19635 12035 19641
rect 11977 19601 11989 19635
rect 12023 19632 12035 19635
rect 12158 19632 12164 19644
rect 12023 19604 12164 19632
rect 12023 19601 12035 19604
rect 11977 19595 12035 19601
rect 12158 19592 12164 19604
rect 12216 19592 12222 19644
rect 12342 19592 12348 19644
rect 12400 19632 12406 19644
rect 12529 19635 12587 19641
rect 12529 19632 12541 19635
rect 12400 19604 12541 19632
rect 12400 19592 12406 19604
rect 12529 19601 12541 19604
rect 12575 19601 12587 19635
rect 12529 19595 12587 19601
rect 12544 19564 12572 19595
rect 12618 19592 12624 19644
rect 12676 19632 12682 19644
rect 12805 19635 12863 19641
rect 12805 19632 12817 19635
rect 12676 19604 12817 19632
rect 12676 19592 12682 19604
rect 12805 19601 12817 19604
rect 12851 19601 12863 19635
rect 13280 19632 13308 19672
rect 12805 19595 12863 19601
rect 12912 19604 13308 19632
rect 15028 19632 15056 19672
rect 22204 19669 22216 19703
rect 22250 19700 22262 19703
rect 23753 19703 23811 19709
rect 23753 19700 23765 19703
rect 22250 19672 23765 19700
rect 22250 19669 22262 19672
rect 22204 19663 22262 19669
rect 23753 19669 23765 19672
rect 23799 19669 23811 19703
rect 23753 19663 23811 19669
rect 15289 19635 15347 19641
rect 15289 19632 15301 19635
rect 15028 19604 15301 19632
rect 12710 19564 12716 19576
rect 12544 19536 12716 19564
rect 7926 19456 7932 19508
rect 7984 19496 7990 19508
rect 8128 19502 8892 19530
rect 12710 19524 12716 19536
rect 12768 19564 12774 19576
rect 12912 19564 12940 19604
rect 15289 19601 15301 19604
rect 15335 19632 15347 19635
rect 16117 19635 16175 19641
rect 16117 19632 16129 19635
rect 15335 19604 16129 19632
rect 15335 19601 15347 19604
rect 15289 19595 15347 19601
rect 16117 19601 16129 19604
rect 16163 19632 16175 19635
rect 16577 19635 16635 19641
rect 16577 19632 16589 19635
rect 16163 19604 16589 19632
rect 16163 19601 16175 19604
rect 16117 19595 16175 19601
rect 16577 19601 16589 19604
rect 16623 19632 16635 19635
rect 16850 19632 16856 19644
rect 16623 19604 16856 19632
rect 16623 19601 16635 19604
rect 16577 19595 16635 19601
rect 16850 19592 16856 19604
rect 16908 19592 16914 19644
rect 17678 19592 17684 19644
rect 17736 19632 17742 19644
rect 17736 19604 17986 19632
rect 17736 19592 17742 19604
rect 12768 19536 12940 19564
rect 12768 19524 12774 19536
rect 8128 19496 8156 19502
rect 7984 19468 8156 19496
rect 8864 19496 8892 19502
rect 9033 19499 9091 19505
rect 9033 19496 9045 19499
rect 8864 19468 9045 19496
rect 7984 19456 7990 19468
rect 9033 19465 9045 19468
rect 9079 19465 9091 19499
rect 9033 19459 9091 19465
rect 10318 19456 10324 19508
rect 10376 19496 10382 19508
rect 10689 19499 10747 19505
rect 10689 19496 10701 19499
rect 10376 19468 10701 19496
rect 10376 19456 10382 19468
rect 10689 19465 10701 19468
rect 10735 19465 10747 19499
rect 10689 19459 10747 19465
rect 11974 19456 11980 19508
rect 12032 19496 12038 19508
rect 12345 19499 12403 19505
rect 12345 19496 12357 19499
rect 12032 19468 12357 19496
rect 12032 19456 12038 19468
rect 12345 19465 12357 19468
rect 12391 19465 12403 19499
rect 13924 19502 14964 19530
rect 17862 19524 17868 19576
rect 17920 19524 17926 19576
rect 22465 19567 22523 19573
rect 22465 19533 22477 19567
rect 22511 19564 22523 19567
rect 22738 19564 22744 19576
rect 22511 19536 22744 19564
rect 22511 19533 22523 19536
rect 22465 19527 22523 19533
rect 22738 19524 22744 19536
rect 22796 19524 22802 19576
rect 13924 19496 13952 19502
rect 12345 19459 12403 19465
rect 13740 19468 13952 19496
rect 14936 19496 14964 19502
rect 15105 19499 15163 19505
rect 15105 19496 15117 19499
rect 14936 19468 15117 19496
rect 8297 19431 8355 19437
rect 8297 19397 8309 19431
rect 8343 19428 8355 19431
rect 8754 19428 8760 19440
rect 8343 19400 8760 19428
rect 8343 19397 8355 19400
rect 8297 19391 8355 19397
rect 8754 19388 8760 19400
rect 8812 19388 8818 19440
rect 9401 19431 9459 19437
rect 9401 19397 9413 19431
rect 9447 19428 9459 19431
rect 9950 19428 9956 19440
rect 9447 19400 9956 19428
rect 9447 19397 9459 19400
rect 9401 19391 9459 19397
rect 9950 19388 9956 19400
rect 10008 19388 10014 19440
rect 11790 19388 11796 19440
rect 11848 19428 11854 19440
rect 11885 19431 11943 19437
rect 11885 19428 11897 19431
rect 11848 19400 11897 19428
rect 11848 19388 11854 19400
rect 11885 19397 11897 19400
rect 11931 19397 11943 19431
rect 11885 19391 11943 19397
rect 13170 19388 13176 19440
rect 13228 19428 13234 19440
rect 13740 19428 13768 19468
rect 15105 19465 15117 19468
rect 15151 19465 15163 19499
rect 15105 19459 15163 19465
rect 16393 19499 16451 19505
rect 16393 19465 16405 19499
rect 16439 19496 16451 19499
rect 17313 19499 17371 19505
rect 17313 19496 17325 19499
rect 16439 19468 17325 19496
rect 16439 19465 16451 19468
rect 16393 19459 16451 19465
rect 17313 19465 17325 19468
rect 17359 19465 17371 19499
rect 17313 19459 17371 19465
rect 18026 19499 18084 19505
rect 18026 19465 18038 19499
rect 18072 19465 18084 19499
rect 18026 19459 18084 19465
rect 14182 19428 14188 19440
rect 13228 19400 13768 19428
rect 14127 19400 14188 19428
rect 13228 19388 13234 19400
rect 14182 19388 14188 19400
rect 14240 19388 14246 19440
rect 14550 19388 14556 19440
rect 14608 19428 14614 19440
rect 15841 19431 15899 19437
rect 15841 19428 15853 19431
rect 14608 19400 15853 19428
rect 14608 19388 14614 19400
rect 15841 19397 15853 19400
rect 15887 19397 15899 19431
rect 15841 19391 15899 19397
rect 17586 19388 17592 19440
rect 17644 19428 17650 19440
rect 18041 19428 18069 19459
rect 17644 19400 18069 19428
rect 19061 19431 19119 19437
rect 17644 19388 17650 19400
rect 19061 19397 19073 19431
rect 19107 19428 19119 19431
rect 19242 19428 19248 19440
rect 19107 19400 19248 19428
rect 19107 19397 19119 19400
rect 19061 19391 19119 19397
rect 19242 19388 19248 19400
rect 19300 19388 19306 19440
rect 5796 19264 23000 19360
rect 6914 19224 6920 19236
rect 6859 19196 6920 19224
rect 6914 19184 6920 19196
rect 6972 19184 6978 19236
rect 10318 19224 10324 19236
rect 10263 19196 10324 19224
rect 10318 19184 10324 19196
rect 10376 19184 10382 19236
rect 15933 19227 15991 19233
rect 15933 19193 15945 19227
rect 15979 19224 15991 19227
rect 17586 19224 17592 19236
rect 15979 19196 16344 19224
rect 15979 19193 15991 19196
rect 15933 19187 15991 19193
rect 10505 19159 10563 19165
rect 10505 19125 10517 19159
rect 10551 19156 10563 19159
rect 11241 19159 11299 19165
rect 11241 19156 11253 19159
rect 10551 19128 11253 19156
rect 10551 19125 10563 19128
rect 10505 19119 10563 19125
rect 11241 19125 11253 19128
rect 11287 19125 11299 19159
rect 11241 19119 11299 19125
rect 12066 19116 12072 19168
rect 12124 19156 12130 19168
rect 12322 19159 12380 19165
rect 12322 19156 12334 19159
rect 12124 19128 12334 19156
rect 12124 19116 12130 19128
rect 12322 19125 12334 19128
rect 12368 19125 12380 19159
rect 12322 19119 12380 19125
rect 12986 19116 12992 19168
rect 13044 19156 13050 19168
rect 13357 19159 13415 19165
rect 13357 19156 13369 19159
rect 13044 19128 13369 19156
rect 13044 19116 13050 19128
rect 13357 19125 13369 19128
rect 13403 19125 13415 19159
rect 13357 19119 13415 19125
rect 14182 19116 14188 19168
rect 14240 19116 14246 19168
rect 14826 19116 14832 19168
rect 14884 19159 14956 19168
rect 14884 19125 14910 19159
rect 14944 19125 14956 19159
rect 16316 19156 16344 19196
rect 17052 19196 17592 19224
rect 17052 19156 17080 19196
rect 17586 19184 17592 19196
rect 17644 19184 17650 19236
rect 21085 19227 21143 19233
rect 21085 19193 21097 19227
rect 21131 19224 21143 19227
rect 22186 19224 22192 19236
rect 21131 19196 21312 19224
rect 21131 19193 21143 19196
rect 21085 19187 21143 19193
rect 16316 19128 17080 19156
rect 14884 19116 14956 19125
rect 19242 19116 19248 19168
rect 19300 19156 19306 19168
rect 20050 19159 20108 19165
rect 20050 19156 20062 19159
rect 19300 19128 20062 19156
rect 19300 19116 19306 19128
rect 20050 19125 20062 19128
rect 20096 19125 20108 19159
rect 21284 19156 21312 19196
rect 21744 19196 22192 19224
rect 21744 19156 21772 19196
rect 22186 19184 22192 19196
rect 22244 19184 22250 19236
rect 21284 19128 21772 19156
rect 20050 19119 20108 19125
rect 8938 19048 8944 19100
rect 8996 19088 9002 19100
rect 9677 19091 9735 19097
rect 9677 19088 9689 19091
rect 8996 19060 9689 19088
rect 8996 19048 9002 19060
rect 9677 19057 9689 19060
rect 9723 19057 9735 19091
rect 9950 19088 9956 19100
rect 9895 19060 9956 19088
rect 9677 19051 9735 19057
rect 9950 19048 9956 19060
rect 10008 19048 10014 19100
rect 11514 19088 11520 19100
rect 11348 19060 11520 19088
rect 6733 19023 6791 19029
rect 6733 18989 6745 19023
rect 6779 19020 6791 19023
rect 6914 19020 6920 19032
rect 6779 18992 6920 19020
rect 6779 18989 6791 18992
rect 6733 18983 6791 18989
rect 6914 18980 6920 18992
rect 6972 18980 6978 19032
rect 10226 18980 10232 19032
rect 10284 19020 10290 19032
rect 10689 19023 10747 19029
rect 10689 19020 10701 19023
rect 10284 18992 10701 19020
rect 10284 18980 10290 18992
rect 10689 18989 10701 18992
rect 10735 19020 10747 19023
rect 10962 19020 10968 19032
rect 10735 18992 10968 19020
rect 10735 18989 10747 18992
rect 10689 18983 10747 18989
rect 10962 18980 10968 18992
rect 11020 18980 11026 19032
rect 11241 19023 11299 19029
rect 11241 18989 11253 19023
rect 11287 19020 11299 19023
rect 11348 19020 11376 19060
rect 11514 19048 11520 19060
rect 11572 19088 11578 19100
rect 11701 19091 11759 19097
rect 11701 19088 11713 19091
rect 11572 19060 11713 19088
rect 11572 19048 11578 19060
rect 11701 19057 11713 19060
rect 11747 19057 11759 19091
rect 11974 19088 11980 19100
rect 11919 19060 11980 19088
rect 11701 19051 11759 19057
rect 11974 19048 11980 19060
rect 12032 19048 12038 19100
rect 14200 19088 14228 19116
rect 14550 19088 14556 19100
rect 13110 19060 14228 19088
rect 14495 19060 14556 19088
rect 14550 19048 14556 19060
rect 14608 19048 14614 19100
rect 16114 19088 16120 19100
rect 15686 19060 16120 19088
rect 16114 19048 16120 19060
rect 16172 19048 16178 19100
rect 20162 19048 20168 19100
rect 20220 19048 20226 19100
rect 11606 19020 11612 19032
rect 11287 18992 11376 19020
rect 11551 18992 11612 19020
rect 11287 18989 11299 18992
rect 11241 18983 11299 18989
rect 11606 18980 11612 18992
rect 11664 18980 11670 19032
rect 11790 18980 11796 19032
rect 11848 18980 11854 19032
rect 13354 19020 13360 19032
rect 13202 18992 13360 19020
rect 13354 18980 13360 18992
rect 13412 18980 13418 19032
rect 17126 19020 17132 19032
rect 15778 18992 17132 19020
rect 17126 18980 17132 18992
rect 17184 18980 17190 19032
rect 17221 19023 17279 19029
rect 17221 18989 17233 19023
rect 17267 19020 17279 19023
rect 17310 19020 17316 19032
rect 17267 18992 17316 19020
rect 17267 18989 17279 18992
rect 17221 18983 17279 18989
rect 17310 18980 17316 18992
rect 17368 18980 17374 19032
rect 17482 19023 17540 19029
rect 17482 18989 17494 19023
rect 17528 19020 17540 19023
rect 17862 19020 17868 19032
rect 17528 18992 17868 19020
rect 17528 18989 17540 18992
rect 17482 18983 17540 18989
rect 17862 18980 17868 18992
rect 17920 18980 17926 19032
rect 20346 18980 20352 19032
rect 20404 18980 20410 19032
rect 22738 18980 22744 19032
rect 22796 19020 22802 19032
rect 22833 19023 22891 19029
rect 22833 19020 22845 19023
rect 22796 18992 22845 19020
rect 22796 18980 22802 18992
rect 22833 18989 22845 18992
rect 22879 18989 22891 19023
rect 22833 18983 22891 18989
rect 11425 18955 11483 18961
rect 5736 18924 6316 18952
rect 5736 18680 5764 18924
rect 6288 18884 6316 18924
rect 11425 18921 11437 18955
rect 11471 18952 11483 18955
rect 11808 18952 11836 18980
rect 11471 18924 11836 18952
rect 22572 18955 22630 18961
rect 11471 18921 11483 18924
rect 11425 18915 11483 18921
rect 22572 18921 22584 18955
rect 22618 18952 22630 18955
rect 22618 18924 23520 18952
rect 22618 18921 22630 18924
rect 22572 18915 22630 18921
rect 6457 18887 6515 18893
rect 6457 18884 6469 18887
rect 6288 18856 6469 18884
rect 6457 18853 6469 18856
rect 6503 18853 6515 18887
rect 6457 18847 6515 18853
rect 9493 18887 9551 18893
rect 9493 18853 9505 18887
rect 9539 18884 9551 18887
rect 9950 18884 9956 18896
rect 9539 18856 9956 18884
rect 9539 18853 9551 18856
rect 9493 18847 9551 18853
rect 9950 18844 9956 18856
rect 10008 18844 10014 18896
rect 10873 18887 10931 18893
rect 10873 18853 10885 18887
rect 10919 18884 10931 18887
rect 10962 18884 10968 18896
rect 10919 18856 10968 18884
rect 10919 18853 10931 18856
rect 10873 18847 10931 18853
rect 10962 18844 10968 18856
rect 11020 18844 11026 18896
rect 17770 18844 17776 18896
rect 17828 18884 17834 18896
rect 18598 18884 18604 18896
rect 17828 18856 18604 18884
rect 17828 18844 17834 18856
rect 18598 18844 18604 18856
rect 18656 18844 18662 18896
rect 19705 18887 19763 18893
rect 19705 18853 19717 18887
rect 19751 18884 19763 18887
rect 20898 18884 20904 18896
rect 19751 18856 20904 18884
rect 19751 18853 19763 18856
rect 19705 18847 19763 18853
rect 20898 18844 20904 18856
rect 20956 18844 20962 18896
rect 21266 18844 21272 18896
rect 21324 18884 21330 18896
rect 23492 18893 23520 18924
rect 21453 18887 21511 18893
rect 21453 18884 21465 18887
rect 21324 18856 21465 18884
rect 21324 18844 21330 18856
rect 21453 18853 21465 18856
rect 21499 18853 21511 18887
rect 21453 18847 21511 18853
rect 23477 18887 23535 18893
rect 23477 18853 23489 18887
rect 23523 18853 23535 18887
rect 23477 18847 23535 18853
rect 5796 18720 23000 18816
rect 6089 18683 6147 18689
rect 6089 18680 6101 18683
rect 5736 18652 6101 18680
rect 6089 18649 6101 18652
rect 6135 18649 6147 18683
rect 6089 18643 6147 18649
rect 8297 18683 8355 18689
rect 8297 18649 8309 18683
rect 8343 18680 8355 18683
rect 8754 18680 8760 18692
rect 8343 18652 8760 18680
rect 8343 18649 8355 18652
rect 8297 18643 8355 18649
rect 8754 18640 8760 18652
rect 8812 18640 8818 18692
rect 12069 18683 12127 18689
rect 12069 18649 12081 18683
rect 12115 18680 12127 18683
rect 12158 18680 12164 18692
rect 12115 18652 12164 18680
rect 12115 18649 12127 18652
rect 12069 18643 12127 18649
rect 12158 18640 12164 18652
rect 12216 18640 12222 18692
rect 12529 18683 12587 18689
rect 12529 18649 12541 18683
rect 12575 18680 12587 18683
rect 13170 18680 13176 18692
rect 12575 18652 13176 18680
rect 12575 18649 12587 18652
rect 12529 18643 12587 18649
rect 13170 18640 13176 18652
rect 13228 18640 13234 18692
rect 19797 18683 19855 18689
rect 19797 18649 19809 18683
rect 19843 18680 19855 18683
rect 20070 18680 20076 18692
rect 19843 18652 20076 18680
rect 19843 18649 19855 18652
rect 19797 18643 19855 18649
rect 20070 18640 20076 18652
rect 20128 18640 20134 18692
rect 20898 18640 20904 18692
rect 20956 18680 20962 18692
rect 21821 18683 21879 18689
rect 21821 18680 21833 18683
rect 20956 18652 21833 18680
rect 20956 18640 20962 18652
rect 21821 18649 21833 18652
rect 21867 18649 21879 18683
rect 21821 18643 21879 18649
rect 22281 18683 22339 18689
rect 22281 18649 22293 18683
rect 22327 18680 22339 18683
rect 22922 18680 22928 18692
rect 22327 18652 22928 18680
rect 22327 18649 22339 18652
rect 22281 18643 22339 18649
rect 22922 18640 22928 18652
rect 22980 18640 22986 18692
rect 14001 18615 14059 18621
rect 14001 18581 14013 18615
rect 14047 18612 14059 18615
rect 14826 18612 14832 18624
rect 14047 18584 14832 18612
rect 14047 18581 14059 18584
rect 6730 18544 6736 18556
rect 6675 18516 6736 18544
rect 6730 18504 6736 18516
rect 6788 18504 6794 18556
rect 7653 18547 7711 18553
rect 7653 18513 7665 18547
rect 7699 18544 7711 18547
rect 7852 18550 8984 18578
rect 14001 18575 14059 18581
rect 14826 18572 14832 18584
rect 14884 18572 14890 18624
rect 16114 18572 16120 18624
rect 16172 18612 16178 18624
rect 17052 18615 17110 18621
rect 17052 18612 17064 18615
rect 16172 18584 17064 18612
rect 16172 18572 16178 18584
rect 17052 18581 17064 18584
rect 17098 18581 17110 18615
rect 17052 18575 17110 18581
rect 17586 18572 17592 18624
rect 17644 18612 17650 18624
rect 17681 18615 17739 18621
rect 17681 18612 17693 18615
rect 17644 18584 17693 18612
rect 17644 18572 17650 18584
rect 17681 18581 17693 18584
rect 17727 18581 17739 18615
rect 17681 18575 17739 18581
rect 17770 18572 17776 18624
rect 17828 18612 17834 18624
rect 17828 18584 17889 18612
rect 17828 18572 17834 18584
rect 20162 18572 20168 18624
rect 20220 18612 20226 18624
rect 20334 18615 20392 18621
rect 20334 18612 20346 18615
rect 20220 18584 20346 18612
rect 20220 18572 20226 18584
rect 20334 18581 20346 18584
rect 20380 18581 20392 18615
rect 20334 18575 20392 18581
rect 7852 18544 7880 18550
rect 7699 18516 7880 18544
rect 8956 18544 8984 18550
rect 9122 18544 9128 18556
rect 8956 18516 9128 18544
rect 7699 18513 7711 18516
rect 7653 18507 7711 18513
rect 9122 18504 9128 18516
rect 9180 18504 9186 18556
rect 10962 18553 10968 18556
rect 10950 18547 10968 18553
rect 10950 18544 10962 18547
rect 10907 18516 10962 18544
rect 10950 18513 10962 18516
rect 10950 18507 10968 18513
rect 10962 18504 10968 18507
rect 11020 18504 11026 18556
rect 13446 18504 13452 18556
rect 13504 18504 13510 18556
rect 15562 18504 15568 18556
rect 15620 18544 15626 18556
rect 17497 18547 17555 18553
rect 17497 18544 17509 18547
rect 15620 18516 17509 18544
rect 15620 18504 15626 18516
rect 17497 18513 17509 18516
rect 17543 18513 17555 18547
rect 17862 18544 17868 18556
rect 17807 18516 17868 18544
rect 17497 18507 17555 18513
rect 17862 18504 17868 18516
rect 17920 18504 17926 18556
rect 19337 18547 19395 18553
rect 19337 18513 19349 18547
rect 19383 18544 19395 18547
rect 20548 18550 21128 18578
rect 21634 18572 21640 18624
rect 21692 18572 21698 18624
rect 20548 18544 20576 18550
rect 19383 18516 20576 18544
rect 21100 18544 21128 18550
rect 21652 18544 21680 18572
rect 21100 18516 21680 18544
rect 22097 18547 22155 18553
rect 19383 18513 19395 18516
rect 19337 18507 19395 18513
rect 22097 18513 22109 18547
rect 22143 18544 22155 18547
rect 22186 18544 22192 18556
rect 22143 18516 22192 18544
rect 22143 18513 22155 18516
rect 22097 18507 22155 18513
rect 22186 18504 22192 18516
rect 22244 18544 22250 18556
rect 22922 18544 22928 18556
rect 22244 18516 22928 18544
rect 22244 18504 22250 18516
rect 22922 18504 22928 18516
rect 22980 18504 22986 18556
rect 6641 18479 6699 18485
rect 6641 18445 6653 18479
rect 6687 18445 6699 18479
rect 6641 18439 6699 18445
rect 7929 18479 7987 18485
rect 7929 18445 7941 18479
rect 7975 18476 7987 18479
rect 7975 18448 8248 18476
rect 7975 18445 7987 18448
rect 7929 18439 7987 18445
rect 6656 18408 6684 18439
rect 7469 18411 7527 18417
rect 7469 18408 7481 18411
rect 6656 18380 7481 18408
rect 7469 18377 7481 18380
rect 7515 18377 7527 18411
rect 8220 18408 8248 18448
rect 8662 18436 8668 18488
rect 8720 18476 8726 18488
rect 8757 18479 8815 18485
rect 8757 18476 8769 18479
rect 8720 18448 8769 18476
rect 8720 18436 8726 18448
rect 8757 18445 8769 18448
rect 8803 18445 8815 18479
rect 9030 18476 9036 18488
rect 8975 18448 9036 18476
rect 8757 18439 8815 18445
rect 9030 18436 9036 18448
rect 9088 18436 9094 18488
rect 10686 18476 10692 18488
rect 10631 18448 10692 18476
rect 10686 18436 10692 18448
rect 10744 18436 10750 18488
rect 14550 18476 14556 18488
rect 13662 18448 14556 18476
rect 14550 18436 14556 18448
rect 14608 18436 14614 18488
rect 17310 18436 17316 18488
rect 17368 18476 17374 18488
rect 17678 18476 17684 18488
rect 17368 18448 17684 18476
rect 17368 18436 17374 18448
rect 17678 18436 17684 18448
rect 17736 18436 17742 18488
rect 19613 18479 19671 18485
rect 19613 18445 19625 18479
rect 19659 18476 19671 18479
rect 19659 18448 19840 18476
rect 19659 18445 19671 18448
rect 19613 18439 19671 18445
rect 8573 18411 8631 18417
rect 8573 18408 8585 18411
rect 8220 18380 8585 18408
rect 7469 18371 7527 18377
rect 8573 18377 8585 18380
rect 8619 18377 8631 18411
rect 8573 18371 8631 18377
rect 12874 18411 12932 18417
rect 12874 18377 12886 18411
rect 12920 18408 12932 18411
rect 12986 18408 12992 18420
rect 12920 18380 12992 18408
rect 12920 18377 12932 18380
rect 12874 18371 12932 18377
rect 12986 18368 12992 18380
rect 13044 18368 13050 18420
rect 6546 18300 6552 18352
rect 6604 18340 6610 18352
rect 6917 18343 6975 18349
rect 6917 18340 6929 18343
rect 6604 18312 6929 18340
rect 6604 18300 6610 18312
rect 6917 18309 6929 18312
rect 6963 18309 6975 18343
rect 6917 18303 6975 18309
rect 8846 18300 8852 18352
rect 8904 18340 8910 18352
rect 9401 18343 9459 18349
rect 9401 18340 9413 18343
rect 8904 18312 9413 18340
rect 8904 18300 8910 18312
rect 9401 18309 9413 18312
rect 9447 18309 9459 18343
rect 9401 18303 9459 18309
rect 15746 18300 15752 18352
rect 15804 18340 15810 18352
rect 15933 18343 15991 18349
rect 15933 18340 15945 18343
rect 15804 18312 15945 18340
rect 15804 18300 15810 18312
rect 15933 18309 15945 18312
rect 15979 18309 15991 18343
rect 15933 18303 15991 18309
rect 18049 18343 18107 18349
rect 18049 18309 18061 18343
rect 18095 18340 18107 18343
rect 18414 18340 18420 18352
rect 18095 18312 18420 18340
rect 18095 18309 18107 18312
rect 18049 18303 18107 18309
rect 18414 18300 18420 18312
rect 18472 18300 18478 18352
rect 18874 18300 18880 18352
rect 18932 18340 18938 18352
rect 18969 18343 19027 18349
rect 18969 18340 18981 18343
rect 18932 18312 18981 18340
rect 18932 18300 18938 18312
rect 18969 18309 18981 18312
rect 19015 18309 19027 18343
rect 19812 18340 19840 18448
rect 19886 18436 19892 18488
rect 19944 18476 19950 18488
rect 20073 18479 20131 18485
rect 20073 18476 20085 18479
rect 19944 18448 20085 18476
rect 19944 18436 19950 18448
rect 20073 18445 20085 18448
rect 20119 18445 20131 18479
rect 20073 18439 20131 18445
rect 20346 18340 20352 18352
rect 19812 18312 20352 18340
rect 18969 18303 19027 18309
rect 20346 18300 20352 18312
rect 20404 18300 20410 18352
rect 21453 18343 21511 18349
rect 21453 18309 21465 18343
rect 21499 18340 21511 18343
rect 21818 18340 21824 18352
rect 21499 18312 21824 18340
rect 21499 18309 21511 18312
rect 21453 18303 21511 18309
rect 21818 18300 21824 18312
rect 21876 18300 21882 18352
rect 5796 18176 23000 18272
rect 7837 18139 7895 18145
rect 7837 18105 7849 18139
rect 7883 18136 7895 18139
rect 8846 18136 8852 18148
rect 7883 18108 8064 18136
rect 7883 18105 7895 18108
rect 7837 18099 7895 18105
rect 6733 18071 6791 18077
rect 6733 18037 6745 18071
rect 6779 18068 6791 18071
rect 7466 18068 7472 18080
rect 6779 18040 7472 18068
rect 6779 18037 6791 18040
rect 6733 18031 6791 18037
rect 7466 18028 7472 18040
rect 7524 18028 7530 18080
rect 8036 18068 8064 18108
rect 8680 18108 8852 18136
rect 8680 18068 8708 18108
rect 8846 18096 8852 18108
rect 8904 18096 8910 18148
rect 9030 18096 9036 18148
rect 9088 18136 9094 18148
rect 9677 18139 9735 18145
rect 9677 18136 9689 18139
rect 9088 18108 9689 18136
rect 9088 18096 9094 18108
rect 9677 18105 9689 18108
rect 9723 18105 9735 18139
rect 9677 18099 9735 18105
rect 8036 18040 8708 18068
rect 11974 18028 11980 18080
rect 12032 18068 12038 18080
rect 12176 18074 12848 18102
rect 13262 18096 13268 18148
rect 13320 18136 13326 18148
rect 16301 18139 16359 18145
rect 16301 18136 16313 18139
rect 13320 18108 15148 18136
rect 13320 18096 13326 18108
rect 12176 18068 12204 18074
rect 12032 18040 12204 18068
rect 12820 18068 12848 18074
rect 13012 18071 13070 18077
rect 13012 18068 13024 18071
rect 12820 18040 13024 18068
rect 12032 18028 12038 18040
rect 13012 18037 13024 18040
rect 13058 18037 13070 18071
rect 15120 18068 15148 18108
rect 15856 18108 16313 18136
rect 15856 18068 15884 18108
rect 16301 18105 16313 18108
rect 16347 18105 16359 18139
rect 16301 18099 16359 18105
rect 21177 18139 21235 18145
rect 21177 18105 21189 18139
rect 21223 18136 21235 18139
rect 26418 18136 26424 18148
rect 21223 18108 26424 18136
rect 21223 18105 21235 18108
rect 21177 18099 21235 18105
rect 26418 18096 26424 18108
rect 26476 18096 26482 18148
rect 15120 18040 15884 18068
rect 16025 18071 16083 18077
rect 13012 18031 13070 18037
rect 16025 18037 16037 18071
rect 16071 18068 16083 18071
rect 16482 18068 16488 18080
rect 16071 18040 16488 18068
rect 16071 18037 16083 18040
rect 16025 18031 16083 18037
rect 16482 18028 16488 18040
rect 16540 18028 16546 18080
rect 17678 18068 17684 18080
rect 17623 18040 17684 18068
rect 17678 18028 17684 18040
rect 17736 18028 17742 18080
rect 22744 18012 22796 18018
rect 9950 17960 9956 18012
rect 10008 18000 10014 18012
rect 10008 17972 10069 18000
rect 10428 17972 11192 18000
rect 10008 17960 10014 17972
rect 6549 17935 6607 17941
rect 6549 17901 6561 17935
rect 6595 17932 6607 17935
rect 6914 17932 6920 17944
rect 6595 17904 6920 17932
rect 6595 17901 6607 17904
rect 6549 17895 6607 17901
rect 6914 17892 6920 17904
rect 6972 17932 6978 17944
rect 7561 17935 7619 17941
rect 7561 17932 7573 17935
rect 6972 17904 7573 17932
rect 6972 17892 6978 17904
rect 7561 17901 7573 17904
rect 7607 17932 7619 17935
rect 9582 17932 9588 17944
rect 7607 17904 9588 17932
rect 7607 17901 7619 17904
rect 7561 17895 7619 17901
rect 9582 17892 9588 17904
rect 9640 17892 9646 17944
rect 9766 17892 9772 17944
rect 9824 17932 9830 17944
rect 9861 17935 9919 17941
rect 9861 17932 9873 17935
rect 9824 17904 9873 17932
rect 9824 17892 9830 17904
rect 9861 17901 9873 17904
rect 9907 17901 9919 17935
rect 9861 17895 9919 17901
rect 10226 17892 10232 17944
rect 10284 17932 10290 17944
rect 10428 17932 10456 17972
rect 10284 17904 10456 17932
rect 11164 17932 11192 17972
rect 11330 17960 11336 18012
rect 11388 18000 11394 18012
rect 11793 18003 11851 18009
rect 11793 18000 11805 18003
rect 11388 17972 11805 18000
rect 11388 17960 11394 17972
rect 11793 17969 11805 17972
rect 11839 17969 11851 18003
rect 11793 17963 11851 17969
rect 11885 18003 11943 18009
rect 11885 17969 11897 18003
rect 11931 18000 11943 18003
rect 12066 18000 12072 18012
rect 11931 17972 12072 18000
rect 11931 17969 11943 17972
rect 11885 17963 11943 17969
rect 12066 17960 12072 17972
rect 12124 17960 12130 18012
rect 12250 17960 12256 18012
rect 12308 17960 12314 18012
rect 16577 18003 16635 18009
rect 16577 17969 16589 18003
rect 16623 17969 16635 18003
rect 22741 18000 22744 18009
rect 22680 17972 22744 18000
rect 16577 17963 16635 17969
rect 22741 17963 22744 17972
rect 11609 17935 11667 17941
rect 11609 17932 11621 17935
rect 11164 17904 11621 17932
rect 10284 17892 10290 17904
rect 11609 17901 11621 17904
rect 11655 17901 11667 17935
rect 11609 17895 11667 17901
rect 12158 17892 12164 17944
rect 12216 17892 12222 17944
rect 14001 17935 14059 17941
rect 14001 17901 14013 17935
rect 14047 17932 14059 17935
rect 15473 17935 15531 17941
rect 14047 17904 14412 17932
rect 14047 17901 14059 17904
rect 14001 17895 14059 17901
rect 14274 17873 14280 17876
rect 14262 17867 14280 17873
rect 14262 17864 14274 17867
rect 14219 17836 14274 17864
rect 14262 17833 14274 17836
rect 14262 17827 14280 17833
rect 14274 17824 14280 17827
rect 14332 17824 14338 17876
rect 14384 17864 14412 17904
rect 15473 17901 15485 17935
rect 15519 17932 15531 17935
rect 15562 17932 15568 17944
rect 15519 17904 15568 17932
rect 15519 17901 15531 17904
rect 15473 17895 15531 17901
rect 15562 17892 15568 17904
rect 15620 17892 15626 17944
rect 15746 17932 15752 17944
rect 15691 17904 15752 17932
rect 15746 17892 15752 17904
rect 15804 17892 15810 17944
rect 15838 17892 15844 17944
rect 15896 17932 15902 17944
rect 15896 17904 15957 17932
rect 15896 17892 15902 17904
rect 16022 17892 16028 17944
rect 16080 17932 16086 17944
rect 16592 17932 16620 17963
rect 22796 17963 22799 18009
rect 22744 17954 22796 17960
rect 19800 17944 19852 17950
rect 16080 17904 16620 17932
rect 16080 17892 16086 17904
rect 17310 17892 17316 17944
rect 17368 17892 17374 17944
rect 19797 17932 19800 17941
rect 19736 17904 19800 17932
rect 19797 17895 19800 17904
rect 19852 17895 19855 17941
rect 20058 17935 20116 17941
rect 20058 17901 20070 17935
rect 20104 17932 20116 17935
rect 21269 17935 21327 17941
rect 21269 17932 21281 17935
rect 20104 17904 20300 17932
rect 20104 17901 20116 17904
rect 20058 17895 20116 17901
rect 19800 17886 19852 17892
rect 14458 17864 14464 17876
rect 14384 17836 14464 17864
rect 14458 17824 14464 17836
rect 14516 17824 14522 17876
rect 15657 17867 15715 17873
rect 15657 17833 15669 17867
rect 15703 17864 15715 17867
rect 16298 17864 16304 17876
rect 15703 17836 16304 17864
rect 15703 17833 15715 17836
rect 15657 17827 15715 17833
rect 16298 17824 16304 17836
rect 16356 17824 16362 17876
rect 20272 17864 20300 17904
rect 20824 17904 21281 17932
rect 20824 17864 20852 17904
rect 21269 17901 21281 17904
rect 21315 17932 21327 17935
rect 21450 17932 21456 17944
rect 21315 17904 21456 17932
rect 21315 17901 21327 17904
rect 21269 17895 21327 17901
rect 21450 17892 21456 17904
rect 21508 17892 21514 17944
rect 22462 17932 22468 17944
rect 22520 17941 22526 17944
rect 22520 17935 22538 17941
rect 22419 17904 22468 17932
rect 22462 17892 22468 17904
rect 22526 17901 22538 17935
rect 22520 17895 22538 17901
rect 22520 17892 22526 17895
rect 20272 17836 20852 17864
rect 7098 17756 7104 17808
rect 7156 17796 7162 17808
rect 7377 17799 7435 17805
rect 7377 17796 7389 17799
rect 7156 17768 7389 17796
rect 7156 17756 7162 17768
rect 7377 17765 7389 17768
rect 7423 17765 7435 17799
rect 7377 17759 7435 17765
rect 10318 17756 10324 17808
rect 10376 17796 10382 17808
rect 10505 17799 10563 17805
rect 10505 17796 10517 17799
rect 10376 17768 10517 17796
rect 10376 17756 10382 17768
rect 10505 17765 10517 17768
rect 10551 17765 10563 17799
rect 10505 17759 10563 17765
rect 10962 17756 10968 17808
rect 11020 17796 11026 17808
rect 11425 17799 11483 17805
rect 11425 17796 11437 17799
rect 11020 17768 11437 17796
rect 11020 17756 11026 17768
rect 11425 17765 11437 17768
rect 11471 17765 11483 17799
rect 13354 17796 13360 17808
rect 13299 17768 13360 17796
rect 11425 17759 11483 17765
rect 13354 17756 13360 17768
rect 13412 17756 13418 17808
rect 14826 17756 14832 17808
rect 14884 17796 14890 17808
rect 15381 17799 15439 17805
rect 15381 17796 15393 17799
rect 14884 17768 15393 17796
rect 14884 17756 14890 17768
rect 15381 17765 15393 17768
rect 15427 17765 15439 17799
rect 15381 17759 15439 17765
rect 21177 17799 21235 17805
rect 21177 17765 21189 17799
rect 21223 17796 21235 17799
rect 21450 17796 21456 17808
rect 21223 17768 21456 17796
rect 21223 17765 21235 17768
rect 21177 17759 21235 17765
rect 21450 17756 21456 17768
rect 21508 17756 21514 17808
rect 5796 17632 23000 17728
rect 9582 17552 9588 17604
rect 9640 17592 9646 17604
rect 12161 17595 12219 17601
rect 9640 17564 10456 17592
rect 9640 17552 9646 17564
rect 9401 17527 9459 17533
rect 9401 17493 9413 17527
rect 9447 17524 9459 17527
rect 9766 17524 9772 17536
rect 9447 17496 9772 17524
rect 9447 17493 9459 17496
rect 9401 17487 9459 17493
rect 9766 17484 9772 17496
rect 9824 17524 9830 17536
rect 9824 17496 10180 17524
rect 9824 17484 9830 17496
rect 10152 17468 10180 17496
rect 7193 17459 7251 17465
rect 7193 17425 7205 17459
rect 7239 17456 7251 17459
rect 7282 17456 7288 17468
rect 7239 17428 7288 17456
rect 7239 17425 7251 17428
rect 7193 17419 7251 17425
rect 7282 17416 7288 17428
rect 7340 17416 7346 17468
rect 7466 17465 7472 17468
rect 7454 17459 7472 17465
rect 7454 17456 7466 17459
rect 7411 17428 7466 17456
rect 7454 17425 7466 17428
rect 7454 17419 7472 17425
rect 7466 17416 7472 17419
rect 7524 17416 7530 17468
rect 8846 17416 8852 17468
rect 8904 17456 8910 17468
rect 9125 17459 9183 17465
rect 9125 17456 9137 17459
rect 8904 17428 9137 17456
rect 8904 17416 8910 17428
rect 9125 17425 9137 17428
rect 9171 17425 9183 17459
rect 9125 17419 9183 17425
rect 9217 17459 9275 17465
rect 9217 17425 9229 17459
rect 9263 17425 9275 17459
rect 9217 17419 9275 17425
rect 6546 17388 6552 17400
rect 6491 17360 6552 17388
rect 6546 17348 6552 17360
rect 6604 17348 6610 17400
rect 6641 17391 6699 17397
rect 6641 17357 6653 17391
rect 6687 17388 6699 17391
rect 9232 17388 9260 17419
rect 10134 17416 10140 17468
rect 10192 17416 10198 17468
rect 10428 17465 10456 17564
rect 12161 17561 12173 17595
rect 12207 17592 12219 17595
rect 12250 17592 12256 17604
rect 12207 17564 12256 17592
rect 12207 17561 12219 17564
rect 12161 17555 12219 17561
rect 12250 17552 12256 17564
rect 12308 17592 12314 17604
rect 14737 17595 14795 17601
rect 12308 17564 12940 17592
rect 12308 17552 12314 17564
rect 12912 17524 12940 17564
rect 14737 17561 14749 17595
rect 14783 17592 14795 17595
rect 21818 17592 21824 17604
rect 14783 17564 14964 17592
rect 14783 17561 14795 17564
rect 14737 17555 14795 17561
rect 13618 17527 13676 17533
rect 13618 17524 13630 17527
rect 11256 17496 11928 17524
rect 12912 17496 13630 17524
rect 10413 17459 10471 17465
rect 10413 17425 10425 17459
rect 10459 17425 10471 17459
rect 10413 17419 10471 17425
rect 10686 17416 10692 17468
rect 10744 17456 10750 17468
rect 10781 17459 10839 17465
rect 10781 17456 10793 17459
rect 10744 17428 10793 17456
rect 10744 17416 10750 17428
rect 10781 17425 10793 17428
rect 10827 17425 10839 17459
rect 10781 17419 10839 17425
rect 11042 17459 11100 17465
rect 11042 17425 11054 17459
rect 11088 17456 11100 17459
rect 11256 17456 11284 17496
rect 11088 17428 11284 17456
rect 11900 17456 11928 17496
rect 13618 17493 13630 17496
rect 13664 17493 13676 17527
rect 13618 17487 13676 17493
rect 14090 17484 14096 17536
rect 14148 17524 14154 17536
rect 14936 17524 14964 17564
rect 20272 17564 20760 17592
rect 15381 17527 15439 17533
rect 15381 17524 15393 17527
rect 14148 17496 14596 17524
rect 14936 17496 15393 17524
rect 14148 17484 14154 17496
rect 12897 17459 12955 17465
rect 12897 17456 12909 17459
rect 11900 17428 12112 17456
rect 11088 17425 11100 17428
rect 11042 17419 11100 17425
rect 6687 17360 7236 17388
rect 6687 17357 6699 17360
rect 6641 17351 6699 17357
rect 6822 17252 6828 17264
rect 6767 17224 6828 17252
rect 6822 17212 6828 17224
rect 6880 17212 6886 17264
rect 7208 17252 7236 17360
rect 8864 17360 9260 17388
rect 10229 17391 10287 17397
rect 8573 17255 8631 17261
rect 8573 17252 8585 17255
rect 7208 17224 8585 17252
rect 8573 17221 8585 17224
rect 8619 17252 8631 17255
rect 8864 17252 8892 17360
rect 10229 17357 10241 17391
rect 10275 17388 10287 17391
rect 10318 17388 10324 17400
rect 10275 17360 10324 17388
rect 10275 17357 10287 17360
rect 10229 17351 10287 17357
rect 10318 17348 10324 17360
rect 10376 17348 10382 17400
rect 12084 17388 12112 17428
rect 12728 17428 12909 17456
rect 12728 17388 12756 17428
rect 12897 17425 12909 17428
rect 12943 17425 12955 17459
rect 12897 17419 12955 17425
rect 12986 17416 12992 17468
rect 13044 17456 13050 17468
rect 13081 17459 13139 17465
rect 13081 17456 13093 17459
rect 13044 17428 13093 17456
rect 13044 17416 13050 17428
rect 13081 17425 13093 17428
rect 13127 17425 13139 17459
rect 13081 17419 13139 17425
rect 13357 17459 13415 17465
rect 13357 17425 13369 17459
rect 13403 17456 13415 17459
rect 14458 17456 14464 17468
rect 13403 17428 14464 17456
rect 13403 17425 13415 17428
rect 13357 17419 13415 17425
rect 14458 17416 14464 17428
rect 14516 17416 14522 17468
rect 14568 17456 14596 17496
rect 15381 17493 15393 17496
rect 15427 17493 15439 17527
rect 15381 17487 15439 17493
rect 18340 17496 18920 17524
rect 15289 17459 15347 17465
rect 15289 17456 15301 17459
rect 14568 17428 15301 17456
rect 15289 17425 15301 17428
rect 15335 17425 15347 17459
rect 15289 17419 15347 17425
rect 15473 17459 15531 17465
rect 15473 17425 15485 17459
rect 15519 17456 15531 17459
rect 15519 17428 15608 17456
rect 15519 17425 15531 17428
rect 15473 17419 15531 17425
rect 12084 17360 12756 17388
rect 13265 17323 13323 17329
rect 13265 17289 13277 17323
rect 13311 17320 13323 17323
rect 13354 17320 13360 17332
rect 13311 17292 13360 17320
rect 13311 17289 13323 17292
rect 13265 17283 13323 17289
rect 13354 17280 13360 17292
rect 13412 17280 13418 17332
rect 8619 17224 8892 17252
rect 8619 17221 8631 17224
rect 8573 17215 8631 17221
rect 9030 17212 9036 17264
rect 9088 17252 9094 17264
rect 9125 17255 9183 17261
rect 9125 17252 9137 17255
rect 9088 17224 9137 17252
rect 9088 17212 9094 17224
rect 9125 17221 9137 17224
rect 9171 17221 9183 17255
rect 9125 17215 9183 17221
rect 10318 17212 10324 17264
rect 10376 17252 10382 17264
rect 10597 17255 10655 17261
rect 10597 17252 10609 17255
rect 10376 17224 10609 17252
rect 10376 17212 10382 17224
rect 10597 17221 10609 17224
rect 10643 17221 10655 17255
rect 10597 17215 10655 17221
rect 14734 17212 14740 17264
rect 14792 17252 14798 17264
rect 15105 17255 15163 17261
rect 15105 17252 15117 17255
rect 14792 17224 15117 17252
rect 14792 17212 14798 17224
rect 15105 17221 15117 17224
rect 15151 17221 15163 17255
rect 15304 17252 15332 17419
rect 15580 17388 15608 17428
rect 15654 17416 15660 17468
rect 15712 17456 15718 17468
rect 15712 17428 15773 17456
rect 15948 17428 16988 17456
rect 15712 17416 15718 17428
rect 15948 17388 15976 17428
rect 15580 17360 15976 17388
rect 16960 17388 16988 17428
rect 17678 17416 17684 17468
rect 17736 17456 17742 17468
rect 17865 17459 17923 17465
rect 17865 17456 17877 17459
rect 17736 17428 17877 17456
rect 17736 17416 17742 17428
rect 17865 17425 17877 17428
rect 17911 17425 17923 17459
rect 17865 17419 17923 17425
rect 18126 17459 18184 17465
rect 18126 17425 18138 17459
rect 18172 17456 18184 17459
rect 18340 17456 18368 17496
rect 18172 17428 18368 17456
rect 18172 17425 18184 17428
rect 18126 17419 18184 17425
rect 17126 17388 17132 17400
rect 16960 17360 17132 17388
rect 17126 17348 17132 17360
rect 17184 17348 17190 17400
rect 18892 17388 18920 17496
rect 19702 17484 19708 17536
rect 19760 17524 19766 17536
rect 19760 17496 19821 17524
rect 19760 17484 19766 17496
rect 19518 17456 19524 17468
rect 19463 17428 19524 17456
rect 19518 17416 19524 17428
rect 19576 17416 19582 17468
rect 19613 17459 19671 17465
rect 19613 17425 19625 17459
rect 19659 17456 19671 17459
rect 20272 17456 20300 17564
rect 20732 17524 20760 17564
rect 21376 17564 21824 17592
rect 21376 17524 21404 17564
rect 21818 17552 21824 17564
rect 21876 17552 21882 17604
rect 20732 17496 21404 17524
rect 22186 17456 22192 17468
rect 22244 17465 22250 17468
rect 22244 17459 22262 17465
rect 19659 17428 20300 17456
rect 22143 17428 22192 17456
rect 19659 17425 19671 17428
rect 19613 17419 19671 17425
rect 22186 17416 22192 17428
rect 22250 17425 22262 17459
rect 22244 17419 22262 17425
rect 22465 17459 22523 17465
rect 22465 17425 22477 17459
rect 22511 17456 22523 17459
rect 22738 17456 22744 17468
rect 22511 17428 22744 17456
rect 22511 17425 22523 17428
rect 22465 17419 22523 17425
rect 22244 17416 22250 17419
rect 22738 17416 22744 17428
rect 22796 17416 22802 17468
rect 18892 17360 19472 17388
rect 19444 17354 19472 17360
rect 16132 17292 16712 17320
rect 15838 17252 15844 17264
rect 15304 17224 15844 17252
rect 15105 17215 15163 17221
rect 15838 17212 15844 17224
rect 15896 17252 15902 17264
rect 16132 17252 16160 17292
rect 15896 17224 16160 17252
rect 16684 17252 16712 17292
rect 16850 17252 16856 17264
rect 16684 17224 16856 17252
rect 15896 17212 15902 17224
rect 16850 17212 16856 17224
rect 16908 17252 16914 17264
rect 17052 17258 17724 17286
rect 19058 17280 19064 17332
rect 19116 17320 19122 17332
rect 19245 17323 19303 17329
rect 19444 17326 20576 17354
rect 19245 17320 19257 17323
rect 19116 17292 19257 17320
rect 19116 17280 19122 17292
rect 19245 17289 19257 17292
rect 19291 17289 19303 17323
rect 20548 17320 20576 17326
rect 21082 17320 21088 17332
rect 20548 17292 21088 17320
rect 19245 17283 19303 17289
rect 21082 17280 21088 17292
rect 21140 17280 21146 17332
rect 17052 17252 17080 17258
rect 16908 17224 17080 17252
rect 17696 17252 17724 17258
rect 17862 17252 17868 17264
rect 17696 17224 17868 17252
rect 16908 17212 16914 17224
rect 17862 17212 17868 17224
rect 17920 17212 17926 17264
rect 18598 17212 18604 17264
rect 18656 17252 18662 17264
rect 19337 17255 19395 17261
rect 19337 17252 19349 17255
rect 18656 17224 19349 17252
rect 18656 17212 18662 17224
rect 19337 17221 19349 17224
rect 19383 17221 19395 17255
rect 19337 17215 19395 17221
rect 20073 17255 20131 17261
rect 20073 17221 20085 17255
rect 20119 17252 20131 17255
rect 20162 17252 20168 17264
rect 20119 17224 20168 17252
rect 20119 17221 20131 17224
rect 20073 17215 20131 17221
rect 20162 17212 20168 17224
rect 20220 17212 20226 17264
rect 5796 17088 23000 17184
rect 9493 17051 9551 17057
rect 9493 17017 9505 17051
rect 9539 17048 9551 17051
rect 10134 17048 10140 17060
rect 9539 17020 10140 17048
rect 9539 17017 9551 17020
rect 9493 17011 9551 17017
rect 10134 17008 10140 17020
rect 10192 17008 10198 17060
rect 11330 17048 11336 17060
rect 11275 17020 11336 17048
rect 11330 17008 11336 17020
rect 11388 17008 11394 17060
rect 11974 17048 11980 17060
rect 11919 17020 11980 17048
rect 11974 17008 11980 17020
rect 12032 17008 12038 17060
rect 14277 17051 14335 17057
rect 14277 17017 14289 17051
rect 14323 17048 14335 17051
rect 15286 17048 15292 17060
rect 14323 17020 15292 17048
rect 14323 17017 14335 17020
rect 14277 17011 14335 17017
rect 15286 17008 15292 17020
rect 15344 17008 15350 17060
rect 16298 17008 16304 17060
rect 16356 17048 16362 17060
rect 16761 17051 16819 17057
rect 16761 17048 16773 17051
rect 16356 17020 16773 17048
rect 16356 17008 16362 17020
rect 16761 17017 16773 17020
rect 16807 17017 16819 17051
rect 16761 17011 16819 17017
rect 19702 17008 19708 17060
rect 19760 17048 19766 17060
rect 20165 17051 20223 17057
rect 20165 17048 20177 17051
rect 19760 17020 20177 17048
rect 19760 17008 19766 17020
rect 20165 17017 20177 17020
rect 20211 17017 20223 17051
rect 20165 17011 20223 17017
rect 12066 16940 12072 16992
rect 12124 16980 12130 16992
rect 13004 16983 13062 16989
rect 13004 16980 13016 16983
rect 12124 16952 13016 16980
rect 12124 16940 12130 16952
rect 13004 16949 13016 16952
rect 13050 16949 13062 16983
rect 13004 16943 13062 16949
rect 10870 16912 10876 16924
rect 10815 16884 10876 16912
rect 10870 16872 10876 16884
rect 10928 16872 10934 16924
rect 11701 16915 11759 16921
rect 11701 16881 11713 16915
rect 11747 16912 11759 16915
rect 11747 16884 11928 16912
rect 11747 16881 11759 16884
rect 11701 16875 11759 16881
rect 11900 16856 11928 16884
rect 12894 16872 12900 16924
rect 12952 16872 12958 16924
rect 14274 16912 14280 16924
rect 14016 16884 14280 16912
rect 10318 16804 10324 16856
rect 10376 16844 10382 16856
rect 10612 16847 10670 16853
rect 10612 16844 10624 16847
rect 10376 16816 10624 16844
rect 10376 16804 10382 16816
rect 10612 16813 10624 16816
rect 10658 16813 10670 16847
rect 10612 16807 10670 16813
rect 11517 16847 11575 16853
rect 11517 16813 11529 16847
rect 11563 16844 11575 16847
rect 11606 16844 11612 16856
rect 11563 16816 11612 16844
rect 11563 16813 11575 16816
rect 11517 16807 11575 16813
rect 11606 16804 11612 16816
rect 11664 16804 11670 16856
rect 11790 16844 11796 16856
rect 11735 16816 11796 16844
rect 11790 16804 11796 16816
rect 11848 16804 11854 16856
rect 11882 16804 11888 16856
rect 11940 16844 11946 16856
rect 11940 16816 12190 16844
rect 11940 16804 11946 16816
rect 13262 16804 13268 16856
rect 13320 16844 13326 16856
rect 14016 16853 14044 16884
rect 14274 16872 14280 16884
rect 14332 16872 14338 16924
rect 18138 16912 18144 16924
rect 18083 16884 18144 16912
rect 18138 16872 18144 16884
rect 18196 16912 18202 16924
rect 18785 16915 18843 16921
rect 18785 16912 18797 16915
rect 18196 16884 18797 16912
rect 18196 16872 18202 16884
rect 18785 16881 18797 16884
rect 18831 16881 18843 16915
rect 18785 16875 18843 16881
rect 20070 16872 20076 16924
rect 20128 16912 20134 16924
rect 23474 16912 23480 16924
rect 20128 16884 23480 16912
rect 20128 16872 20134 16884
rect 23474 16872 23480 16884
rect 23532 16872 23538 16924
rect 13909 16847 13967 16853
rect 13909 16844 13921 16847
rect 13320 16816 13921 16844
rect 13320 16804 13326 16816
rect 13909 16813 13921 16816
rect 13955 16813 13967 16847
rect 13909 16807 13967 16813
rect 14001 16847 14059 16853
rect 14001 16813 14013 16847
rect 14047 16813 14059 16847
rect 14001 16807 14059 16813
rect 14090 16804 14096 16856
rect 14148 16844 14154 16856
rect 14369 16847 14427 16853
rect 14148 16816 14209 16844
rect 14148 16804 14154 16816
rect 14369 16813 14381 16847
rect 14415 16844 14427 16847
rect 14458 16844 14464 16856
rect 14415 16816 14464 16844
rect 14415 16813 14427 16816
rect 14369 16807 14427 16813
rect 14458 16804 14464 16816
rect 14516 16804 14522 16856
rect 14642 16853 14648 16856
rect 14630 16847 14648 16853
rect 14630 16844 14642 16847
rect 14587 16816 14642 16844
rect 14630 16813 14642 16816
rect 14630 16807 14648 16813
rect 14642 16804 14648 16807
rect 14700 16804 14706 16856
rect 15562 16844 15568 16856
rect 15396 16816 15568 16844
rect 13633 16779 13691 16785
rect 13633 16745 13645 16779
rect 13679 16776 13691 16779
rect 15396 16776 15424 16816
rect 15562 16804 15568 16816
rect 15620 16804 15626 16856
rect 16040 16816 16528 16844
rect 13679 16748 15424 16776
rect 15841 16779 15899 16785
rect 13679 16745 13691 16748
rect 13633 16739 13691 16745
rect 15841 16745 15853 16779
rect 15887 16776 15899 16779
rect 16040 16776 16068 16816
rect 15887 16748 16068 16776
rect 16500 16776 16528 16816
rect 18414 16804 18420 16856
rect 18472 16844 18478 16856
rect 19046 16847 19104 16853
rect 19046 16844 19058 16847
rect 18472 16816 19058 16844
rect 18472 16804 18478 16816
rect 19046 16813 19058 16816
rect 19092 16813 19104 16847
rect 20898 16844 20904 16856
rect 20843 16816 20904 16844
rect 19046 16807 19104 16813
rect 20898 16804 20904 16816
rect 20956 16804 20962 16856
rect 16666 16776 16672 16788
rect 16500 16748 16672 16776
rect 15887 16745 15899 16748
rect 15841 16739 15899 16745
rect 16666 16736 16672 16748
rect 16724 16736 16730 16788
rect 17770 16736 17776 16788
rect 17828 16776 17834 16788
rect 17880 16779 17938 16785
rect 17880 16776 17892 16779
rect 17828 16748 17892 16776
rect 17828 16736 17834 16748
rect 17880 16745 17892 16748
rect 17926 16745 17938 16779
rect 20714 16776 20720 16788
rect 20659 16748 20720 16776
rect 17880 16739 17938 16745
rect 20714 16736 20720 16748
rect 20772 16736 20778 16788
rect 20809 16779 20867 16785
rect 20809 16745 20821 16779
rect 20855 16776 20867 16779
rect 21450 16776 21456 16788
rect 20855 16748 21456 16776
rect 20855 16745 20867 16748
rect 20809 16739 20867 16745
rect 21450 16736 21456 16748
rect 21508 16736 21514 16788
rect 13078 16668 13084 16720
rect 13136 16708 13142 16720
rect 13357 16711 13415 16717
rect 13357 16708 13369 16711
rect 13136 16680 13369 16708
rect 13136 16668 13142 16680
rect 13357 16677 13369 16680
rect 13403 16677 13415 16711
rect 13357 16671 13415 16677
rect 20070 16668 20076 16720
rect 20128 16708 20134 16720
rect 20162 16708 20168 16720
rect 20128 16680 20168 16708
rect 20128 16668 20134 16680
rect 20162 16668 20168 16680
rect 20220 16708 20226 16720
rect 20441 16711 20499 16717
rect 20441 16708 20453 16711
rect 20220 16680 20453 16708
rect 20220 16668 20226 16680
rect 20441 16677 20453 16680
rect 20487 16677 20499 16711
rect 20441 16671 20499 16677
rect 20990 16668 20996 16720
rect 21048 16708 21054 16720
rect 21177 16711 21235 16717
rect 21177 16708 21189 16711
rect 21048 16680 21189 16708
rect 21048 16668 21054 16680
rect 21177 16677 21189 16680
rect 21223 16677 21235 16711
rect 21177 16671 21235 16677
rect 5796 16544 23000 16640
rect 8757 16507 8815 16513
rect 8757 16473 8769 16507
rect 8803 16504 8815 16507
rect 8846 16504 8852 16516
rect 8803 16476 8852 16504
rect 8803 16473 8815 16476
rect 8757 16467 8815 16473
rect 8846 16464 8852 16476
rect 8904 16464 8910 16516
rect 11606 16464 11612 16516
rect 11664 16504 11670 16516
rect 11793 16507 11851 16513
rect 11793 16504 11805 16507
rect 11664 16476 11805 16504
rect 11664 16464 11670 16476
rect 11793 16473 11805 16476
rect 11839 16473 11851 16507
rect 11793 16467 11851 16473
rect 13078 16464 13084 16516
rect 13136 16504 13142 16516
rect 13173 16507 13231 16513
rect 13173 16504 13185 16507
rect 13136 16476 13185 16504
rect 13136 16464 13142 16476
rect 13173 16473 13185 16476
rect 13219 16473 13231 16507
rect 13173 16467 13231 16473
rect 13262 16464 13268 16516
rect 13320 16504 13326 16516
rect 13357 16507 13415 16513
rect 13357 16504 13369 16507
rect 13320 16476 13369 16504
rect 13320 16464 13326 16476
rect 13357 16473 13369 16476
rect 13403 16473 13415 16507
rect 13357 16467 13415 16473
rect 15746 16464 15752 16516
rect 15804 16504 15810 16516
rect 15804 16476 16068 16504
rect 15804 16464 15810 16476
rect 10588 16449 10646 16455
rect 7009 16439 7067 16445
rect 7009 16405 7021 16439
rect 7055 16436 7067 16439
rect 7638 16439 7696 16445
rect 7638 16436 7650 16439
rect 7055 16408 7650 16436
rect 7055 16405 7067 16408
rect 7009 16399 7067 16405
rect 7638 16405 7650 16408
rect 7684 16405 7696 16439
rect 7638 16399 7696 16405
rect 7926 16396 7932 16448
rect 7984 16436 7990 16448
rect 7984 16408 9168 16436
rect 10588 16415 10600 16449
rect 10634 16436 10646 16449
rect 10962 16436 10968 16448
rect 10634 16415 10968 16436
rect 10588 16409 10968 16415
rect 10603 16408 10968 16409
rect 7984 16396 7990 16408
rect 6178 16368 6184 16380
rect 6123 16340 6184 16368
rect 6178 16328 6184 16340
rect 6236 16328 6242 16380
rect 6825 16371 6883 16377
rect 6825 16337 6837 16371
rect 6871 16368 6883 16371
rect 6914 16368 6920 16380
rect 6871 16340 6920 16368
rect 6871 16337 6883 16340
rect 6825 16331 6883 16337
rect 6914 16328 6920 16340
rect 6972 16328 6978 16380
rect 7282 16328 7288 16380
rect 7340 16368 7346 16380
rect 7377 16371 7435 16377
rect 7377 16368 7389 16371
rect 7340 16340 7389 16368
rect 7340 16328 7346 16340
rect 7377 16337 7389 16340
rect 7423 16337 7435 16371
rect 9030 16368 9036 16380
rect 8975 16340 9036 16368
rect 7377 16331 7435 16337
rect 9030 16328 9036 16340
rect 9088 16328 9094 16380
rect 9140 16377 9168 16408
rect 10962 16396 10968 16408
rect 11020 16396 11026 16448
rect 12802 16396 12808 16448
rect 12860 16396 12866 16448
rect 14476 16439 14534 16445
rect 14476 16405 14488 16439
rect 14522 16436 14534 16439
rect 14826 16436 14832 16448
rect 14522 16408 14832 16436
rect 14522 16405 14534 16408
rect 14476 16399 14534 16405
rect 14826 16396 14832 16408
rect 14884 16396 14890 16448
rect 15378 16445 15384 16448
rect 15366 16439 15384 16445
rect 15366 16436 15378 16439
rect 15323 16408 15378 16436
rect 15366 16405 15378 16408
rect 15366 16399 15384 16405
rect 15378 16396 15384 16399
rect 15436 16396 15442 16448
rect 9125 16371 9183 16377
rect 9125 16337 9137 16371
rect 9171 16337 9183 16371
rect 9125 16331 9183 16337
rect 10321 16371 10379 16377
rect 10321 16337 10333 16371
rect 10367 16368 10379 16371
rect 10594 16368 10600 16380
rect 10367 16340 10600 16368
rect 10367 16337 10379 16340
rect 10321 16331 10379 16337
rect 10594 16328 10600 16340
rect 10652 16328 10658 16380
rect 11606 16328 11612 16380
rect 11664 16368 11670 16380
rect 11793 16371 11851 16377
rect 11793 16368 11805 16371
rect 11664 16340 11805 16368
rect 11664 16328 11670 16340
rect 11793 16337 11805 16340
rect 11839 16337 11851 16371
rect 11793 16331 11851 16337
rect 11885 16371 11943 16377
rect 11885 16337 11897 16371
rect 11931 16368 11943 16371
rect 11974 16368 11980 16380
rect 11931 16340 11980 16368
rect 11931 16337 11943 16340
rect 11885 16331 11943 16337
rect 11974 16328 11980 16340
rect 12032 16328 12038 16380
rect 12820 16368 12848 16396
rect 12897 16371 12955 16377
rect 12897 16368 12909 16371
rect 12820 16340 12909 16368
rect 12897 16337 12909 16340
rect 12943 16368 12955 16371
rect 13354 16368 13360 16380
rect 12943 16340 13360 16368
rect 12943 16337 12955 16340
rect 12897 16331 12955 16337
rect 13354 16328 13360 16340
rect 13412 16328 13418 16380
rect 14737 16371 14795 16377
rect 14737 16337 14749 16371
rect 14783 16368 14795 16371
rect 15105 16371 15163 16377
rect 15105 16368 15117 16371
rect 14783 16340 15117 16368
rect 14783 16337 14795 16340
rect 14737 16331 14795 16337
rect 15105 16337 15117 16340
rect 15151 16368 15163 16371
rect 15930 16368 15936 16380
rect 15151 16340 15936 16368
rect 15151 16337 15163 16340
rect 15105 16331 15163 16337
rect 15930 16328 15936 16340
rect 15988 16328 15994 16380
rect 16040 16368 16068 16476
rect 16666 16464 16672 16516
rect 16724 16504 16730 16516
rect 17313 16507 17371 16513
rect 16724 16476 16988 16504
rect 16724 16464 16730 16476
rect 16960 16445 16988 16476
rect 17313 16473 17325 16507
rect 17359 16504 17371 16507
rect 17770 16504 17776 16516
rect 17359 16476 17776 16504
rect 17359 16473 17371 16476
rect 17313 16467 17371 16473
rect 17770 16464 17776 16476
rect 17828 16464 17834 16516
rect 19889 16507 19947 16513
rect 19889 16473 19901 16507
rect 19935 16504 19947 16507
rect 20714 16504 20720 16516
rect 19935 16476 20720 16504
rect 19935 16473 19947 16476
rect 19889 16467 19947 16473
rect 20714 16464 20720 16476
rect 20772 16464 20778 16516
rect 21453 16507 21511 16513
rect 21453 16473 21465 16507
rect 21499 16504 21511 16507
rect 21634 16504 21640 16516
rect 21499 16476 21640 16504
rect 21499 16473 21511 16476
rect 21453 16467 21511 16473
rect 21634 16464 21640 16476
rect 21692 16464 21698 16516
rect 22005 16507 22063 16513
rect 22005 16473 22017 16507
rect 22051 16504 22063 16507
rect 22186 16504 22192 16516
rect 22051 16476 22192 16504
rect 22051 16473 22063 16476
rect 22005 16467 22063 16473
rect 22186 16464 22192 16476
rect 22244 16464 22250 16516
rect 22370 16464 22376 16516
rect 22428 16504 22434 16516
rect 22465 16507 22523 16513
rect 22465 16504 22477 16507
rect 22428 16476 22477 16504
rect 22428 16464 22434 16476
rect 22465 16473 22477 16476
rect 22511 16473 22523 16507
rect 22465 16467 22523 16473
rect 16577 16439 16635 16445
rect 16577 16405 16589 16439
rect 16623 16436 16635 16439
rect 16853 16439 16911 16445
rect 16853 16436 16865 16439
rect 16623 16408 16865 16436
rect 16623 16405 16635 16408
rect 16577 16399 16635 16405
rect 16853 16405 16865 16408
rect 16899 16405 16911 16439
rect 16853 16399 16911 16405
rect 16945 16439 17003 16445
rect 16945 16405 16957 16439
rect 16991 16405 17003 16439
rect 16945 16399 17003 16405
rect 18598 16396 18604 16448
rect 18656 16436 18662 16448
rect 20346 16445 20352 16448
rect 18770 16439 18828 16445
rect 18770 16436 18782 16439
rect 18656 16408 18782 16436
rect 18656 16396 18662 16408
rect 18770 16405 18782 16408
rect 18816 16405 18828 16439
rect 20334 16439 20352 16445
rect 20334 16436 20346 16439
rect 20291 16408 20346 16436
rect 18770 16399 18828 16405
rect 20334 16405 20346 16408
rect 20334 16399 20352 16405
rect 20346 16396 20352 16399
rect 20404 16396 20410 16448
rect 16666 16368 16672 16380
rect 16040 16340 16672 16368
rect 16666 16328 16672 16340
rect 16724 16328 16730 16380
rect 17037 16371 17095 16377
rect 17037 16368 17049 16371
rect 16868 16340 17049 16368
rect 16868 16312 16896 16340
rect 17037 16337 17049 16340
rect 17083 16337 17095 16371
rect 17037 16331 17095 16337
rect 19886 16328 19892 16380
rect 19944 16368 19950 16380
rect 20073 16371 20131 16377
rect 20073 16368 20085 16371
rect 19944 16340 20085 16368
rect 19944 16328 19950 16340
rect 20073 16337 20085 16340
rect 20119 16337 20131 16371
rect 20073 16331 20131 16337
rect 6273 16303 6331 16309
rect 6273 16269 6285 16303
rect 6319 16300 6331 16303
rect 8846 16300 8852 16312
rect 6319 16272 6776 16300
rect 8791 16272 8852 16300
rect 6319 16269 6331 16272
rect 6273 16263 6331 16269
rect 6748 16232 6776 16272
rect 8846 16260 8852 16272
rect 8904 16260 8910 16312
rect 9401 16303 9459 16309
rect 9401 16269 9413 16303
rect 9447 16300 9459 16303
rect 9858 16300 9864 16312
rect 9447 16272 9864 16300
rect 9447 16269 9459 16272
rect 9401 16263 9459 16269
rect 9858 16260 9864 16272
rect 9916 16300 9922 16312
rect 9953 16303 10011 16309
rect 9953 16300 9965 16303
rect 9916 16272 9965 16300
rect 9916 16260 9922 16272
rect 9953 16269 9965 16272
rect 9999 16269 10011 16303
rect 9953 16263 10011 16269
rect 16850 16260 16856 16312
rect 16908 16260 16914 16312
rect 17954 16260 17960 16312
rect 18012 16300 18018 16312
rect 18509 16303 18567 16309
rect 18509 16300 18521 16303
rect 18012 16272 18521 16300
rect 18012 16260 18018 16272
rect 18509 16269 18521 16272
rect 18555 16269 18567 16303
rect 18509 16263 18567 16269
rect 22189 16303 22247 16309
rect 22189 16269 22201 16303
rect 22235 16300 22247 16303
rect 22278 16300 22284 16312
rect 22235 16272 22284 16300
rect 22235 16269 22247 16272
rect 22189 16263 22247 16269
rect 22278 16260 22284 16272
rect 22336 16300 22342 16312
rect 22922 16300 22928 16312
rect 22336 16272 22928 16300
rect 22336 16260 22342 16272
rect 22922 16260 22928 16272
rect 22980 16260 22986 16312
rect 9214 16232 9220 16244
rect 6748 16204 7420 16232
rect 9159 16204 9220 16232
rect 7392 16164 7420 16204
rect 9214 16192 9220 16204
rect 9272 16192 9278 16244
rect 9769 16235 9827 16241
rect 9769 16201 9781 16235
rect 9815 16232 9827 16235
rect 10226 16232 10232 16244
rect 9815 16204 10232 16232
rect 9815 16201 9827 16204
rect 9769 16195 9827 16201
rect 10226 16192 10232 16204
rect 10284 16192 10290 16244
rect 11701 16235 11759 16241
rect 11701 16201 11713 16235
rect 11747 16232 11759 16235
rect 11882 16232 11888 16244
rect 11747 16204 11888 16232
rect 11747 16201 11759 16204
rect 11701 16195 11759 16201
rect 11882 16192 11888 16204
rect 11940 16232 11946 16244
rect 12161 16235 12219 16241
rect 12161 16232 12173 16235
rect 11940 16204 12173 16232
rect 11940 16192 11946 16204
rect 12161 16201 12173 16204
rect 12207 16201 12219 16235
rect 12161 16195 12219 16201
rect 8757 16167 8815 16173
rect 8757 16164 8769 16167
rect 7392 16136 8769 16164
rect 8757 16133 8769 16136
rect 8803 16133 8815 16167
rect 8757 16127 8815 16133
rect 9030 16124 9036 16176
rect 9088 16164 9094 16176
rect 9125 16167 9183 16173
rect 9125 16164 9137 16167
rect 9088 16136 9137 16164
rect 9088 16124 9094 16136
rect 9125 16133 9137 16136
rect 9171 16133 9183 16167
rect 9125 16127 9183 16133
rect 9585 16167 9643 16173
rect 9585 16133 9597 16167
rect 9631 16164 9643 16167
rect 10042 16164 10048 16176
rect 9631 16136 10048 16164
rect 9631 16133 9643 16136
rect 9585 16127 9643 16133
rect 10042 16124 10048 16136
rect 10100 16124 10106 16176
rect 10137 16167 10195 16173
rect 10137 16133 10149 16167
rect 10183 16164 10195 16167
rect 10962 16164 10968 16176
rect 10183 16136 10968 16164
rect 10183 16133 10195 16136
rect 10137 16127 10195 16133
rect 10962 16124 10968 16136
rect 11020 16124 11026 16176
rect 12710 16164 12716 16176
rect 12655 16136 12716 16164
rect 12710 16124 12716 16136
rect 12768 16124 12774 16176
rect 21266 16124 21272 16176
rect 21324 16164 21330 16176
rect 21453 16167 21511 16173
rect 21453 16164 21465 16167
rect 21324 16136 21465 16164
rect 21324 16124 21330 16136
rect 21453 16133 21465 16136
rect 21499 16133 21511 16167
rect 21453 16127 21511 16133
rect 5796 16000 23000 16096
rect 6914 15920 6920 15972
rect 6972 15960 6978 15972
rect 8573 15963 8631 15969
rect 6972 15932 8064 15960
rect 6972 15920 6978 15932
rect 8036 15892 8064 15932
rect 8573 15929 8585 15963
rect 8619 15960 8631 15963
rect 8846 15960 8852 15972
rect 8619 15932 8852 15960
rect 8619 15929 8631 15932
rect 8573 15923 8631 15929
rect 8846 15920 8852 15932
rect 8904 15920 8910 15972
rect 9401 15963 9459 15969
rect 9401 15929 9413 15963
rect 9447 15960 9459 15963
rect 11146 15960 11152 15972
rect 9447 15932 11152 15960
rect 9447 15929 9459 15932
rect 9401 15923 9459 15929
rect 11146 15920 11152 15932
rect 11204 15920 11210 15972
rect 11790 15960 11796 15972
rect 11735 15932 11796 15960
rect 11790 15920 11796 15932
rect 11848 15920 11854 15972
rect 12986 15920 12992 15972
rect 13044 15960 13050 15972
rect 13449 15963 13507 15969
rect 13449 15960 13461 15963
rect 13044 15932 13461 15960
rect 13044 15920 13050 15932
rect 13449 15929 13461 15932
rect 13495 15960 13507 15963
rect 13495 15932 14044 15960
rect 13495 15929 13507 15932
rect 13449 15923 13507 15929
rect 9030 15892 9036 15904
rect 8036 15864 8616 15892
rect 8975 15864 9036 15892
rect 6917 15759 6975 15765
rect 6917 15725 6929 15759
rect 6963 15756 6975 15759
rect 7190 15756 7196 15768
rect 6963 15728 7196 15756
rect 6963 15725 6975 15728
rect 6917 15719 6975 15725
rect 7190 15716 7196 15728
rect 7248 15716 7254 15768
rect 7466 15716 7472 15768
rect 7524 15716 7530 15768
rect 7926 15716 7932 15768
rect 7984 15756 7990 15768
rect 8481 15759 8539 15765
rect 8481 15756 8493 15759
rect 7984 15728 8493 15756
rect 7984 15716 7990 15728
rect 8481 15725 8493 15728
rect 8527 15725 8539 15759
rect 8588 15756 8616 15864
rect 9030 15852 9036 15864
rect 9088 15852 9094 15904
rect 8938 15756 8944 15768
rect 8588 15728 8944 15756
rect 8481 15719 8539 15725
rect 8938 15716 8944 15728
rect 8996 15756 9002 15768
rect 9217 15759 9275 15765
rect 9217 15756 9229 15759
rect 8996 15728 9229 15756
rect 8996 15716 9002 15728
rect 9217 15725 9229 15728
rect 9263 15725 9275 15759
rect 9490 15756 9496 15768
rect 9435 15728 9496 15756
rect 9217 15719 9275 15725
rect 9490 15716 9496 15728
rect 9548 15716 9554 15768
rect 9754 15759 9812 15765
rect 9754 15725 9766 15759
rect 9800 15756 9812 15759
rect 10042 15756 10048 15768
rect 9800 15728 10048 15756
rect 9800 15725 9812 15728
rect 9754 15719 9812 15725
rect 10042 15716 10048 15728
rect 10100 15716 10106 15768
rect 10778 15716 10784 15768
rect 10836 15756 10842 15768
rect 10965 15759 11023 15765
rect 10965 15756 10977 15759
rect 10836 15728 10977 15756
rect 10836 15716 10842 15728
rect 10965 15725 10977 15728
rect 11011 15725 11023 15759
rect 11425 15759 11483 15765
rect 11425 15756 11437 15759
rect 10965 15719 11023 15725
rect 11348 15728 11437 15756
rect 7184 15682 7242 15688
rect 7184 15648 7196 15682
rect 7230 15679 7242 15682
rect 7484 15679 7512 15716
rect 7230 15651 7512 15679
rect 7230 15648 7242 15651
rect 10410 15648 10416 15700
rect 10468 15688 10474 15700
rect 11348 15688 11376 15728
rect 11425 15725 11437 15728
rect 11471 15756 11483 15759
rect 11606 15756 11612 15768
rect 11471 15728 11612 15756
rect 11471 15725 11483 15728
rect 11425 15719 11483 15725
rect 11606 15716 11612 15728
rect 11664 15716 11670 15768
rect 12069 15759 12127 15765
rect 12069 15725 12081 15759
rect 12115 15756 12127 15759
rect 12342 15756 12348 15768
rect 12115 15728 12348 15756
rect 12115 15725 12127 15728
rect 12069 15719 12127 15725
rect 12342 15716 12348 15728
rect 12400 15716 12406 15768
rect 12434 15688 12440 15700
rect 10468 15660 11376 15688
rect 12330 15682 12440 15688
rect 10468 15648 10474 15660
rect 12330 15648 12342 15682
rect 12376 15660 12440 15682
rect 12376 15648 12388 15660
rect 12434 15648 12440 15660
rect 12492 15648 12498 15700
rect 14016 15688 14044 15932
rect 16850 15852 16856 15904
rect 16908 15892 16914 15904
rect 16908 15864 17816 15892
rect 16908 15852 16914 15864
rect 16666 15824 16672 15836
rect 16611 15796 16672 15824
rect 16666 15784 16672 15796
rect 16724 15784 16730 15836
rect 17788 15824 17816 15864
rect 18432 15864 18828 15892
rect 18432 15824 18460 15864
rect 17788 15796 18460 15824
rect 14369 15759 14427 15765
rect 14369 15725 14381 15759
rect 14415 15756 14427 15759
rect 14458 15756 14464 15768
rect 14415 15728 14464 15756
rect 14415 15725 14427 15728
rect 14369 15719 14427 15725
rect 14458 15716 14464 15728
rect 14516 15716 14522 15768
rect 16485 15759 16543 15765
rect 16485 15725 16497 15759
rect 16531 15756 16543 15759
rect 16942 15756 16948 15768
rect 16531 15728 16948 15756
rect 16531 15725 16543 15728
rect 16485 15719 16543 15725
rect 16942 15716 16948 15728
rect 17000 15716 17006 15768
rect 17316 15700 17368 15706
rect 14630 15691 14688 15697
rect 14630 15688 14642 15691
rect 14016 15660 14642 15688
rect 14630 15657 14642 15660
rect 14676 15657 14688 15691
rect 14630 15651 14688 15657
rect 14844 15660 15608 15688
rect 7184 15642 7242 15648
rect 12330 15642 12388 15648
rect 8297 15623 8355 15629
rect 8297 15589 8309 15623
rect 8343 15620 8355 15623
rect 8754 15620 8760 15632
rect 8343 15592 8760 15620
rect 8343 15589 8355 15592
rect 8297 15583 8355 15589
rect 8754 15580 8760 15592
rect 8812 15580 8818 15632
rect 10226 15580 10232 15632
rect 10284 15620 10290 15632
rect 11333 15623 11391 15629
rect 11333 15620 11345 15623
rect 10284 15592 11345 15620
rect 10284 15580 10290 15592
rect 11333 15589 11345 15592
rect 11379 15589 11391 15623
rect 11333 15583 11391 15589
rect 14274 15580 14280 15632
rect 14332 15620 14338 15632
rect 14844 15620 14872 15660
rect 14332 15592 14872 15620
rect 15580 15620 15608 15660
rect 17420 15688 17448 15742
rect 18598 15716 18604 15768
rect 18656 15756 18662 15768
rect 18693 15759 18751 15765
rect 18693 15756 18705 15759
rect 18656 15728 18705 15756
rect 18656 15716 18662 15728
rect 18693 15725 18705 15728
rect 18739 15725 18751 15759
rect 18800 15756 18828 15864
rect 19429 15827 19487 15833
rect 19429 15793 19441 15827
rect 19475 15824 19487 15827
rect 20070 15824 20076 15836
rect 19475 15796 20076 15824
rect 19475 15793 19487 15796
rect 19429 15787 19487 15793
rect 20070 15784 20076 15796
rect 20128 15784 20134 15836
rect 22738 15824 22744 15836
rect 22683 15796 22744 15824
rect 22738 15784 22744 15796
rect 22796 15784 22802 15836
rect 18969 15759 19027 15765
rect 18969 15756 18981 15759
rect 18800 15728 18981 15756
rect 18693 15719 18751 15725
rect 18969 15725 18981 15728
rect 19015 15725 19027 15759
rect 18969 15719 19027 15725
rect 17368 15660 17448 15688
rect 17316 15642 17368 15648
rect 15749 15623 15807 15629
rect 15749 15620 15761 15623
rect 15580 15592 15761 15620
rect 14332 15580 14338 15592
rect 15749 15589 15761 15592
rect 15795 15589 15807 15623
rect 17770 15620 17776 15632
rect 17715 15592 17776 15620
rect 15749 15583 15807 15589
rect 17770 15580 17776 15592
rect 17828 15580 17834 15632
rect 18984 15620 19012 15719
rect 19058 15716 19064 15768
rect 19116 15756 19122 15768
rect 20824 15759 20882 15765
rect 19116 15728 19177 15756
rect 19116 15716 19122 15728
rect 20824 15725 20836 15759
rect 20870 15756 20882 15759
rect 20990 15756 20996 15768
rect 20870 15728 20996 15756
rect 20870 15725 20882 15728
rect 20824 15719 20882 15725
rect 20990 15716 20996 15728
rect 21048 15716 21054 15768
rect 21085 15759 21143 15765
rect 21085 15725 21097 15759
rect 21131 15756 21143 15759
rect 21450 15756 21456 15768
rect 21131 15728 21456 15756
rect 21131 15725 21143 15728
rect 21085 15719 21143 15725
rect 21450 15716 21456 15728
rect 21508 15716 21514 15768
rect 19153 15691 19211 15697
rect 19153 15657 19165 15691
rect 19199 15688 19211 15691
rect 19613 15691 19671 15697
rect 19613 15688 19625 15691
rect 19199 15660 19625 15688
rect 19199 15657 19211 15660
rect 19153 15651 19211 15657
rect 19613 15657 19625 15660
rect 19659 15657 19671 15691
rect 19613 15651 19671 15657
rect 21910 15648 21916 15700
rect 21968 15688 21974 15700
rect 22480 15691 22538 15697
rect 22480 15688 22492 15691
rect 21968 15660 22492 15688
rect 21968 15648 21974 15660
rect 22480 15657 22492 15660
rect 22526 15657 22538 15691
rect 22480 15651 22538 15657
rect 19058 15620 19064 15632
rect 18984 15592 19064 15620
rect 19058 15580 19064 15592
rect 19116 15580 19122 15632
rect 21361 15623 21419 15629
rect 21361 15589 21373 15623
rect 21407 15620 21419 15623
rect 21726 15620 21732 15632
rect 21407 15592 21732 15620
rect 21407 15589 21419 15592
rect 21361 15583 21419 15589
rect 21726 15580 21732 15592
rect 21784 15580 21790 15632
rect 5796 15456 23000 15552
rect 6089 15419 6147 15425
rect 6089 15385 6101 15419
rect 6135 15416 6147 15419
rect 6178 15416 6184 15428
rect 6135 15388 6184 15416
rect 6135 15385 6147 15388
rect 6089 15379 6147 15385
rect 6178 15376 6184 15388
rect 6236 15376 6242 15428
rect 9214 15376 9220 15428
rect 9272 15416 9278 15428
rect 9953 15419 10011 15425
rect 9953 15416 9965 15419
rect 9272 15388 9965 15416
rect 9272 15376 9278 15388
rect 9953 15385 9965 15388
rect 9999 15385 10011 15419
rect 9953 15379 10011 15385
rect 16301 15419 16359 15425
rect 16301 15385 16313 15419
rect 16347 15385 16359 15419
rect 16301 15379 16359 15385
rect 8312 15351 8370 15357
rect 8312 15317 8324 15351
rect 8358 15348 8370 15351
rect 9033 15351 9091 15357
rect 9033 15348 9045 15351
rect 8358 15320 9045 15348
rect 8358 15317 8370 15320
rect 8312 15311 8370 15317
rect 9033 15317 9045 15320
rect 9079 15317 9091 15351
rect 9033 15311 9091 15317
rect 12066 15308 12072 15360
rect 12124 15348 12130 15360
rect 12161 15351 12219 15357
rect 12161 15348 12173 15351
rect 12124 15320 12173 15348
rect 12124 15308 12130 15320
rect 12161 15317 12173 15320
rect 12207 15317 12219 15351
rect 15182 15351 15240 15357
rect 15182 15348 15194 15351
rect 12161 15311 12219 15317
rect 14016 15320 15194 15348
rect 6549 15283 6607 15289
rect 6549 15249 6561 15283
rect 6595 15280 6607 15283
rect 6822 15280 6828 15292
rect 6595 15252 6828 15280
rect 6595 15249 6607 15252
rect 6549 15243 6607 15249
rect 6822 15240 6828 15252
rect 6880 15240 6886 15292
rect 7101 15283 7159 15289
rect 7101 15280 7113 15283
rect 6932 15252 7113 15280
rect 6273 15215 6331 15221
rect 6273 15181 6285 15215
rect 6319 15212 6331 15215
rect 6932 15212 6960 15252
rect 7101 15249 7113 15252
rect 7147 15280 7159 15283
rect 7926 15280 7932 15292
rect 7147 15252 7932 15280
rect 7147 15249 7159 15252
rect 7101 15243 7159 15249
rect 7926 15240 7932 15252
rect 7984 15240 7990 15292
rect 8573 15283 8631 15289
rect 8573 15249 8585 15283
rect 8619 15280 8631 15283
rect 8662 15280 8668 15292
rect 8619 15252 8668 15280
rect 8619 15249 8631 15252
rect 8573 15243 8631 15249
rect 8662 15240 8668 15252
rect 8720 15240 8726 15292
rect 8849 15283 8907 15289
rect 8849 15249 8861 15283
rect 8895 15280 8907 15283
rect 8938 15280 8944 15292
rect 8895 15252 8944 15280
rect 8895 15249 8907 15252
rect 8849 15243 8907 15249
rect 8938 15240 8944 15252
rect 8996 15240 9002 15292
rect 10137 15283 10195 15289
rect 10137 15249 10149 15283
rect 10183 15280 10195 15283
rect 10226 15280 10232 15292
rect 10183 15252 10232 15280
rect 10183 15249 10195 15252
rect 10137 15243 10195 15249
rect 10226 15240 10232 15252
rect 10284 15240 10290 15292
rect 10321 15283 10379 15289
rect 10321 15249 10333 15283
rect 10367 15280 10379 15283
rect 10778 15280 10784 15292
rect 10367 15252 10784 15280
rect 10367 15249 10379 15252
rect 10321 15243 10379 15249
rect 10778 15240 10784 15252
rect 10836 15280 10842 15292
rect 10836 15252 10994 15280
rect 10836 15240 10842 15252
rect 11882 15240 11888 15292
rect 11940 15240 11946 15292
rect 12618 15240 12624 15292
rect 12676 15280 12682 15292
rect 14016 15280 14044 15320
rect 15182 15317 15194 15320
rect 15228 15317 15240 15351
rect 16316 15348 16344 15379
rect 16942 15376 16948 15428
rect 17000 15416 17006 15428
rect 17497 15419 17555 15425
rect 17497 15416 17509 15419
rect 17000 15388 17509 15416
rect 17000 15376 17006 15388
rect 17497 15385 17509 15388
rect 17543 15385 17555 15419
rect 17497 15379 17555 15385
rect 18966 15376 18972 15428
rect 19024 15416 19030 15428
rect 22005 15419 22063 15425
rect 22005 15416 22017 15419
rect 19024 15388 19196 15416
rect 19024 15376 19030 15388
rect 16669 15351 16727 15357
rect 16669 15348 16681 15351
rect 16316 15320 16681 15348
rect 15182 15311 15240 15317
rect 16669 15317 16681 15320
rect 16715 15317 16727 15351
rect 19168 15348 19196 15388
rect 20916 15388 21404 15416
rect 20916 15348 20944 15388
rect 19168 15320 20944 15348
rect 16669 15311 16727 15317
rect 21082 15308 21088 15360
rect 21140 15348 21146 15360
rect 21192 15351 21250 15357
rect 21192 15348 21204 15351
rect 21140 15320 21204 15348
rect 21140 15308 21146 15320
rect 21192 15317 21204 15320
rect 21238 15317 21250 15351
rect 21376 15348 21404 15388
rect 21836 15388 22017 15416
rect 21836 15348 21864 15388
rect 22005 15385 22017 15388
rect 22051 15385 22063 15419
rect 22005 15379 22063 15385
rect 21376 15320 21864 15348
rect 21192 15311 21250 15317
rect 14734 15280 14740 15292
rect 12676 15252 14044 15280
rect 14306 15252 14740 15280
rect 12676 15240 12682 15252
rect 14734 15240 14740 15252
rect 14792 15240 14798 15292
rect 15654 15240 15660 15292
rect 15712 15280 15718 15292
rect 16393 15283 16451 15289
rect 16393 15280 16405 15283
rect 15712 15252 16405 15280
rect 15712 15240 15718 15252
rect 16393 15249 16405 15252
rect 16439 15249 16451 15283
rect 16577 15283 16635 15289
rect 16577 15280 16589 15283
rect 16393 15243 16451 15249
rect 16500 15252 16589 15280
rect 6319 15184 6960 15212
rect 6319 15181 6331 15184
rect 6273 15175 6331 15181
rect 10410 15172 10416 15224
rect 10468 15212 10474 15224
rect 10686 15212 10692 15224
rect 10468 15184 10529 15212
rect 10631 15184 10692 15212
rect 10468 15172 10474 15184
rect 10686 15172 10692 15184
rect 10744 15172 10750 15224
rect 11790 15172 11796 15224
rect 11848 15172 11854 15224
rect 13170 15212 13176 15224
rect 13115 15184 13176 15212
rect 13170 15172 13176 15184
rect 13228 15172 13234 15224
rect 16022 15172 16028 15224
rect 16080 15212 16086 15224
rect 16500 15212 16528 15252
rect 16577 15249 16589 15252
rect 16623 15249 16635 15283
rect 16577 15243 16635 15249
rect 16761 15283 16819 15289
rect 16761 15249 16773 15283
rect 16807 15280 16819 15283
rect 16850 15280 16856 15292
rect 16807 15252 16856 15280
rect 16807 15249 16819 15252
rect 16761 15243 16819 15249
rect 16850 15240 16856 15252
rect 16908 15240 16914 15292
rect 18598 15240 18604 15292
rect 18656 15280 18662 15292
rect 18770 15283 18828 15289
rect 18770 15280 18782 15283
rect 18656 15252 18782 15280
rect 18656 15240 18662 15252
rect 18770 15249 18782 15252
rect 18816 15249 18828 15283
rect 18770 15243 18828 15249
rect 16080 15184 16528 15212
rect 16080 15172 16086 15184
rect 17954 15172 17960 15224
rect 18012 15212 18018 15224
rect 18509 15215 18567 15221
rect 18509 15212 18521 15215
rect 18012 15184 18521 15212
rect 18012 15172 18018 15184
rect 18509 15181 18521 15184
rect 18555 15181 18567 15215
rect 21450 15212 21456 15224
rect 21395 15184 21456 15212
rect 18509 15175 18567 15181
rect 21450 15172 21456 15184
rect 21508 15172 21514 15224
rect 22278 15212 22284 15224
rect 22223 15184 22284 15212
rect 22278 15172 22284 15184
rect 22336 15172 22342 15224
rect 6917 15147 6975 15153
rect 6917 15113 6929 15147
rect 6963 15144 6975 15147
rect 8665 15147 8723 15153
rect 8665 15144 8677 15147
rect 6963 15116 7696 15144
rect 6963 15113 6975 15116
rect 6917 15107 6975 15113
rect 7668 15076 7696 15116
rect 8588 15116 8677 15144
rect 8588 15076 8616 15116
rect 8665 15113 8677 15116
rect 8711 15113 8723 15147
rect 8665 15107 8723 15113
rect 11042 15147 11100 15153
rect 11042 15113 11054 15147
rect 11088 15113 11100 15147
rect 13357 15147 13415 15153
rect 13357 15144 13369 15147
rect 11042 15107 11100 15113
rect 13188 15116 13369 15144
rect 7668 15048 8616 15076
rect 11057 15076 11085 15107
rect 11330 15076 11336 15088
rect 11057 15048 11336 15076
rect 11330 15036 11336 15048
rect 11388 15036 11394 15088
rect 12802 15036 12808 15088
rect 12860 15076 12866 15088
rect 13188 15076 13216 15116
rect 13357 15113 13369 15116
rect 13403 15113 13415 15147
rect 14458 15144 14464 15156
rect 14403 15116 14464 15144
rect 13357 15107 13415 15113
rect 13556 15082 14228 15110
rect 14458 15104 14464 15116
rect 14516 15104 14522 15156
rect 19794 15104 19800 15156
rect 19852 15144 19858 15156
rect 20073 15147 20131 15153
rect 20073 15144 20085 15147
rect 19852 15116 20085 15144
rect 19852 15104 19858 15116
rect 20073 15113 20085 15116
rect 20119 15113 20131 15147
rect 20073 15107 20131 15113
rect 13556 15076 13584 15082
rect 12860 15048 13584 15076
rect 14200 15076 14228 15082
rect 15930 15076 15936 15088
rect 14200 15048 15936 15076
rect 12860 15036 12866 15048
rect 15930 15036 15936 15048
rect 15988 15076 15994 15088
rect 16298 15076 16304 15088
rect 15988 15048 16304 15076
rect 15988 15036 15994 15048
rect 16298 15036 16304 15048
rect 16356 15036 16362 15088
rect 16945 15079 17003 15085
rect 16945 15045 16957 15079
rect 16991 15076 17003 15079
rect 17310 15076 17316 15088
rect 16991 15048 17316 15076
rect 16991 15045 17003 15048
rect 16945 15039 17003 15045
rect 17310 15036 17316 15048
rect 17368 15036 17374 15088
rect 19889 15079 19947 15085
rect 19889 15045 19901 15079
rect 19935 15076 19947 15079
rect 19978 15076 19984 15088
rect 19935 15048 19984 15076
rect 19935 15045 19947 15048
rect 19889 15039 19947 15045
rect 19978 15036 19984 15048
rect 20036 15036 20042 15088
rect 22462 15076 22468 15088
rect 22407 15048 22468 15076
rect 22462 15036 22468 15048
rect 22520 15036 22526 15088
rect 5796 14912 23000 15008
rect 8757 14875 8815 14881
rect 8757 14841 8769 14875
rect 8803 14872 8815 14875
rect 10134 14872 10140 14884
rect 8803 14844 10140 14872
rect 8803 14841 8815 14844
rect 8757 14835 8815 14841
rect 10134 14832 10140 14844
rect 10192 14832 10198 14884
rect 10321 14875 10379 14881
rect 10321 14841 10333 14875
rect 10367 14872 10379 14875
rect 10410 14872 10416 14884
rect 10367 14844 10416 14872
rect 10367 14841 10379 14844
rect 10321 14835 10379 14841
rect 10410 14832 10416 14844
rect 10468 14832 10474 14884
rect 10686 14832 10692 14884
rect 10744 14872 10750 14884
rect 10744 14844 10916 14872
rect 10744 14832 10750 14844
rect 9030 14764 9036 14816
rect 9088 14804 9094 14816
rect 9286 14807 9344 14813
rect 9286 14804 9298 14807
rect 9088 14776 9298 14804
rect 9088 14764 9094 14776
rect 9286 14773 9298 14776
rect 9332 14773 9344 14807
rect 10888 14804 10916 14844
rect 11348 14844 12480 14872
rect 11348 14804 11376 14844
rect 10888 14776 11376 14804
rect 12452 14804 12480 14844
rect 17402 14832 17408 14884
rect 17460 14872 17466 14884
rect 17589 14875 17647 14881
rect 17589 14872 17601 14875
rect 17460 14844 17601 14872
rect 17460 14832 17466 14844
rect 17589 14841 17601 14844
rect 17635 14841 17647 14875
rect 17589 14835 17647 14841
rect 20901 14875 20959 14881
rect 20901 14841 20913 14875
rect 20947 14872 20959 14875
rect 20990 14872 20996 14884
rect 20947 14844 20996 14872
rect 20947 14841 20959 14844
rect 20901 14835 20959 14841
rect 20990 14832 20996 14844
rect 21048 14832 21054 14884
rect 13633 14807 13691 14813
rect 13633 14804 13645 14807
rect 12452 14776 13645 14804
rect 9286 14767 9344 14773
rect 13633 14773 13645 14776
rect 13679 14773 13691 14807
rect 13633 14767 13691 14773
rect 20346 14764 20352 14816
rect 20404 14804 20410 14816
rect 21361 14807 21419 14813
rect 21361 14804 21373 14807
rect 20404 14776 21373 14804
rect 20404 14764 20410 14776
rect 21361 14773 21373 14776
rect 21407 14773 21419 14807
rect 21361 14767 21419 14773
rect 22744 14748 22796 14754
rect 6914 14736 6920 14748
rect 6859 14708 6920 14736
rect 6914 14696 6920 14708
rect 6972 14696 6978 14748
rect 8404 14708 9154 14736
rect 6730 14628 6736 14680
rect 6788 14668 6794 14680
rect 8404 14677 8432 14708
rect 18230 14696 18236 14748
rect 18288 14696 18294 14748
rect 18782 14736 18788 14748
rect 18727 14708 18788 14736
rect 18782 14696 18788 14708
rect 18840 14696 18846 14748
rect 20438 14696 20444 14748
rect 20496 14736 20502 14748
rect 22741 14736 22744 14745
rect 20496 14708 20576 14736
rect 22680 14708 22744 14736
rect 20496 14696 20502 14708
rect 7178 14671 7236 14677
rect 7178 14668 7190 14671
rect 6788 14640 7190 14668
rect 6788 14628 6794 14640
rect 7178 14637 7190 14640
rect 7224 14637 7236 14671
rect 7178 14631 7236 14637
rect 8389 14671 8447 14677
rect 8389 14637 8401 14671
rect 8435 14637 8447 14671
rect 10870 14668 10876 14680
rect 10166 14640 10876 14668
rect 8389 14631 8447 14637
rect 10870 14628 10876 14640
rect 10928 14628 10934 14680
rect 10962 14628 10968 14680
rect 11020 14668 11026 14680
rect 12176 14671 12234 14677
rect 12176 14668 12188 14671
rect 11020 14640 11468 14668
rect 11020 14628 11026 14640
rect 11440 14600 11468 14640
rect 11992 14640 12188 14668
rect 11992 14600 12020 14640
rect 12176 14637 12188 14640
rect 12222 14637 12234 14671
rect 12176 14631 12234 14637
rect 12342 14628 12348 14680
rect 12400 14668 12406 14680
rect 12437 14671 12495 14677
rect 12437 14668 12449 14671
rect 12400 14640 12449 14668
rect 12400 14628 12406 14640
rect 12437 14637 12449 14640
rect 12483 14637 12495 14671
rect 12437 14631 12495 14637
rect 13354 14628 13360 14680
rect 13412 14668 13418 14680
rect 13817 14671 13875 14677
rect 13817 14668 13829 14671
rect 13412 14640 13829 14668
rect 13412 14628 13418 14640
rect 13817 14637 13829 14640
rect 13863 14637 13875 14671
rect 14458 14668 14464 14680
rect 14403 14640 14464 14668
rect 13817 14631 13875 14637
rect 14458 14628 14464 14640
rect 14516 14628 14522 14680
rect 16206 14668 16212 14680
rect 16151 14640 16212 14668
rect 16206 14628 16212 14640
rect 16264 14628 16270 14680
rect 16482 14677 16488 14680
rect 16470 14671 16488 14677
rect 16470 14668 16482 14671
rect 16427 14640 16482 14668
rect 16470 14637 16482 14640
rect 16470 14631 16488 14637
rect 16482 14628 16488 14631
rect 16540 14628 16546 14680
rect 18230 14671 18294 14696
rect 17328 14640 18092 14668
rect 14722 14603 14780 14609
rect 14722 14600 14734 14603
rect 7392 14572 8156 14600
rect 11440 14572 12020 14600
rect 14568 14572 14734 14600
rect 7392 14566 7420 14572
rect 6546 14492 6552 14544
rect 6604 14532 6610 14544
rect 6748 14538 7420 14566
rect 6748 14532 6776 14538
rect 6604 14504 6776 14532
rect 8128 14532 8156 14572
rect 14568 14544 14596 14572
rect 14722 14569 14734 14572
rect 14768 14569 14780 14603
rect 14722 14563 14780 14569
rect 15194 14560 15200 14612
rect 15252 14600 15258 14612
rect 17328 14600 17356 14640
rect 15252 14572 16068 14600
rect 15252 14560 15258 14572
rect 16040 14566 16068 14572
rect 16592 14572 17356 14600
rect 18064 14600 18092 14640
rect 18230 14637 18245 14671
rect 18279 14637 18294 14671
rect 18230 14631 18294 14637
rect 18506 14628 18512 14680
rect 18564 14628 18570 14680
rect 20070 14628 20076 14680
rect 20128 14668 20134 14680
rect 20245 14671 20303 14677
rect 20245 14668 20257 14671
rect 20128 14640 20257 14668
rect 20128 14628 20134 14640
rect 20245 14637 20257 14640
rect 20291 14668 20303 14671
rect 20346 14668 20352 14680
rect 20291 14640 20352 14668
rect 20291 14637 20303 14640
rect 20245 14631 20303 14637
rect 20346 14628 20352 14640
rect 20404 14628 20410 14680
rect 20548 14677 20576 14708
rect 22741 14699 22744 14708
rect 22796 14699 22799 14745
rect 22744 14690 22796 14696
rect 20533 14671 20591 14677
rect 20533 14637 20545 14671
rect 20579 14637 20591 14671
rect 22462 14668 22468 14680
rect 22520 14677 22526 14680
rect 22520 14671 22538 14677
rect 20533 14631 20591 14637
rect 20625 14654 20683 14660
rect 20625 14620 20637 14654
rect 20671 14620 20683 14654
rect 22419 14640 22468 14668
rect 22462 14628 22468 14640
rect 22526 14637 22538 14671
rect 22520 14631 22538 14637
rect 22520 14628 22526 14631
rect 20625 14614 20683 14620
rect 18598 14600 18604 14612
rect 18064 14572 18604 14600
rect 16592 14566 16620 14572
rect 8297 14535 8355 14541
rect 8297 14532 8309 14535
rect 8128 14504 8309 14532
rect 6604 14492 6610 14504
rect 8297 14501 8309 14504
rect 8343 14501 8355 14535
rect 8297 14495 8355 14501
rect 13446 14492 13452 14544
rect 13504 14532 13510 14544
rect 14001 14535 14059 14541
rect 14001 14532 14013 14535
rect 13504 14504 14013 14532
rect 13504 14492 13510 14504
rect 14001 14501 14013 14504
rect 14047 14501 14059 14535
rect 14001 14495 14059 14501
rect 14550 14492 14556 14544
rect 14608 14492 14614 14544
rect 15838 14532 15844 14544
rect 15783 14504 15844 14532
rect 15838 14492 15844 14504
rect 15896 14492 15902 14544
rect 16040 14538 16620 14566
rect 18598 14560 18604 14572
rect 18656 14560 18662 14612
rect 18966 14560 18972 14612
rect 19024 14603 19099 14612
rect 19024 14569 19053 14603
rect 19087 14569 19099 14603
rect 19024 14560 19099 14569
rect 19978 14560 19984 14612
rect 20036 14600 20042 14612
rect 20441 14603 20499 14609
rect 20441 14600 20453 14603
rect 20036 14572 20453 14600
rect 20036 14560 20042 14572
rect 20441 14569 20453 14572
rect 20487 14569 20499 14603
rect 20441 14563 20499 14569
rect 20640 14544 20668 14614
rect 20162 14532 20168 14544
rect 20107 14504 20168 14532
rect 20162 14492 20168 14504
rect 20220 14492 20226 14544
rect 20622 14492 20628 14544
rect 20680 14492 20686 14544
rect 5796 14368 23000 14464
rect 10594 14288 10600 14340
rect 10652 14328 10658 14340
rect 10781 14331 10839 14337
rect 10781 14328 10793 14331
rect 10652 14300 10793 14328
rect 10652 14288 10658 14300
rect 10781 14297 10793 14300
rect 10827 14297 10839 14331
rect 10781 14291 10839 14297
rect 11790 14288 11796 14340
rect 11848 14328 11854 14340
rect 14093 14331 14151 14337
rect 14093 14328 14105 14331
rect 11848 14300 12020 14328
rect 11848 14288 11854 14300
rect 11992 14294 12020 14300
rect 12820 14300 14105 14328
rect 12820 14294 12848 14300
rect 11992 14266 12848 14294
rect 14093 14297 14105 14300
rect 14139 14328 14151 14331
rect 14550 14328 14556 14340
rect 14139 14300 14556 14328
rect 14139 14297 14151 14300
rect 14093 14291 14151 14297
rect 14550 14288 14556 14300
rect 14608 14288 14614 14340
rect 17126 14288 17132 14340
rect 17184 14328 17190 14340
rect 17497 14331 17555 14337
rect 17497 14328 17509 14331
rect 17184 14300 17509 14328
rect 17184 14288 17190 14300
rect 17497 14297 17509 14300
rect 17543 14297 17555 14331
rect 18966 14328 18972 14340
rect 18911 14300 18972 14328
rect 17497 14291 17555 14297
rect 18966 14288 18972 14300
rect 19024 14288 19030 14340
rect 21910 14288 21916 14340
rect 21968 14328 21974 14340
rect 22005 14331 22063 14337
rect 22005 14328 22017 14331
rect 21968 14300 22017 14328
rect 21968 14288 21974 14300
rect 22005 14297 22017 14300
rect 22051 14297 22063 14331
rect 22005 14291 22063 14297
rect 12974 14263 13032 14269
rect 12974 14229 12986 14263
rect 13020 14260 13032 14263
rect 13446 14260 13452 14272
rect 13020 14232 13452 14260
rect 13020 14229 13032 14232
rect 12974 14223 13032 14229
rect 13446 14220 13452 14232
rect 13504 14220 13510 14272
rect 14274 14220 14280 14272
rect 14332 14260 14338 14272
rect 14461 14263 14519 14269
rect 14461 14260 14473 14263
rect 14332 14232 14473 14260
rect 14332 14220 14338 14232
rect 14461 14229 14473 14232
rect 14507 14229 14519 14263
rect 14461 14223 14519 14229
rect 15752 14204 15804 14210
rect 6546 14192 6552 14204
rect 6491 14164 6552 14192
rect 6546 14152 6552 14164
rect 6604 14152 6610 14204
rect 7282 14152 7288 14204
rect 7340 14192 7346 14204
rect 7837 14195 7895 14201
rect 7837 14192 7849 14195
rect 7340 14164 7849 14192
rect 7340 14152 7346 14164
rect 7837 14161 7849 14164
rect 7883 14161 7895 14195
rect 7837 14155 7895 14161
rect 7926 14152 7932 14204
rect 7984 14192 7990 14204
rect 8098 14195 8156 14201
rect 8098 14192 8110 14195
rect 7984 14164 8110 14192
rect 7984 14152 7990 14164
rect 8098 14161 8110 14164
rect 8144 14161 8156 14195
rect 8098 14155 8156 14161
rect 11146 14152 11152 14204
rect 11204 14192 11210 14204
rect 11900 14195 11958 14201
rect 11900 14192 11912 14195
rect 11204 14164 11912 14192
rect 11204 14152 11210 14164
rect 11900 14161 11912 14164
rect 11946 14192 11958 14195
rect 12802 14192 12808 14204
rect 11946 14164 12808 14192
rect 11946 14161 11958 14164
rect 11900 14155 11958 14161
rect 12802 14152 12808 14164
rect 12860 14152 12866 14204
rect 14185 14195 14243 14201
rect 14185 14161 14197 14195
rect 14231 14161 14243 14195
rect 14366 14192 14372 14204
rect 14311 14164 14372 14192
rect 14185 14155 14243 14161
rect 6641 14127 6699 14133
rect 6641 14093 6653 14127
rect 6687 14124 6699 14127
rect 6914 14124 6920 14136
rect 6687 14096 6920 14124
rect 6687 14093 6699 14096
rect 6641 14087 6699 14093
rect 6914 14084 6920 14096
rect 6972 14084 6978 14136
rect 12161 14127 12219 14133
rect 12161 14093 12173 14127
rect 12207 14124 12219 14127
rect 12342 14124 12348 14136
rect 12207 14096 12348 14124
rect 12207 14093 12219 14096
rect 12161 14087 12219 14093
rect 12342 14084 12348 14096
rect 12400 14124 12406 14136
rect 12713 14127 12771 14133
rect 12713 14124 12725 14127
rect 12400 14096 12725 14124
rect 12400 14084 12406 14096
rect 12713 14093 12725 14096
rect 12759 14093 12771 14127
rect 14200 14124 14228 14155
rect 14366 14152 14372 14164
rect 14424 14152 14430 14204
rect 14550 14192 14556 14204
rect 14495 14164 14556 14192
rect 14550 14152 14556 14164
rect 14608 14152 14614 14204
rect 14829 14195 14887 14201
rect 14829 14161 14841 14195
rect 14875 14192 14887 14195
rect 15194 14192 15200 14204
rect 14875 14164 15200 14192
rect 14875 14161 14887 14164
rect 14829 14155 14887 14161
rect 15194 14152 15200 14164
rect 15252 14152 15258 14204
rect 16761 14195 16819 14201
rect 16761 14161 16773 14195
rect 16807 14192 16819 14195
rect 16942 14192 16948 14204
rect 16807 14164 16948 14192
rect 16807 14161 16819 14164
rect 16761 14155 16819 14161
rect 16942 14152 16948 14164
rect 17000 14152 17006 14204
rect 18598 14192 18604 14204
rect 18656 14201 18662 14204
rect 18656 14195 18674 14201
rect 18555 14164 18604 14192
rect 18598 14152 18604 14164
rect 18662 14161 18674 14195
rect 18656 14155 18674 14161
rect 18656 14152 18662 14155
rect 18782 14152 18788 14204
rect 18840 14192 18846 14204
rect 18877 14195 18935 14201
rect 18877 14192 18889 14195
rect 18840 14164 18889 14192
rect 18840 14152 18846 14164
rect 18877 14161 18889 14164
rect 18923 14161 18935 14195
rect 18877 14155 18935 14161
rect 19058 14152 19064 14204
rect 19116 14192 19122 14204
rect 19245 14195 19303 14201
rect 19245 14192 19257 14195
rect 19116 14164 19257 14192
rect 19116 14152 19122 14164
rect 19245 14161 19257 14164
rect 19291 14161 19303 14195
rect 19245 14155 19303 14161
rect 19337 14195 19395 14201
rect 19337 14161 19349 14195
rect 19383 14161 19395 14195
rect 19337 14155 19395 14161
rect 19429 14195 19487 14201
rect 19429 14161 19441 14195
rect 19475 14161 19487 14195
rect 19429 14155 19487 14161
rect 19613 14195 19671 14201
rect 19613 14161 19625 14195
rect 19659 14192 19671 14195
rect 20346 14192 20352 14204
rect 19659 14164 20352 14192
rect 19659 14161 19671 14164
rect 19613 14155 19671 14161
rect 15752 14146 15804 14152
rect 15562 14124 15568 14136
rect 14200 14096 14412 14124
rect 12713 14087 12771 14093
rect 14384 14056 14412 14096
rect 15212 14096 15568 14124
rect 15212 14056 15240 14096
rect 15562 14084 15568 14096
rect 15620 14084 15626 14136
rect 16574 14084 16580 14136
rect 16632 14124 16638 14136
rect 16632 14096 16693 14124
rect 16632 14084 16638 14096
rect 15470 14056 15476 14068
rect 14384 14028 15240 14056
rect 15415 14028 15476 14056
rect 15470 14016 15476 14028
rect 15528 14016 15534 14068
rect 6273 13991 6331 13997
rect 6273 13988 6285 13991
rect 5736 13960 6285 13988
rect 5736 13784 5764 13960
rect 6273 13957 6285 13960
rect 6319 13957 6331 13991
rect 6273 13951 6331 13957
rect 9122 13948 9128 14000
rect 9180 13988 9186 14000
rect 9217 13991 9275 13997
rect 9217 13988 9229 13991
rect 9180 13960 9229 13988
rect 9180 13948 9186 13960
rect 9217 13957 9229 13960
rect 9263 13957 9275 13991
rect 9217 13951 9275 13957
rect 10781 13991 10839 13997
rect 10781 13957 10793 13991
rect 10827 13988 10839 13991
rect 11790 13988 11796 14000
rect 10827 13960 11796 13988
rect 10827 13957 10839 13960
rect 10781 13951 10839 13957
rect 11790 13948 11796 13960
rect 11848 13948 11854 14000
rect 19352 13988 19380 14155
rect 19444 14124 19472 14155
rect 20346 14152 20352 14164
rect 20404 14152 20410 14204
rect 21266 14192 21272 14204
rect 21324 14201 21330 14204
rect 21324 14195 21342 14201
rect 21223 14164 21272 14192
rect 21266 14152 21272 14164
rect 21330 14161 21342 14195
rect 21324 14155 21342 14161
rect 21324 14152 21330 14155
rect 21450 14152 21456 14204
rect 21508 14192 21514 14204
rect 21545 14195 21603 14201
rect 21545 14192 21557 14195
rect 21508 14164 21557 14192
rect 21508 14152 21514 14164
rect 21545 14161 21557 14164
rect 21591 14161 21603 14195
rect 21545 14155 21603 14161
rect 22189 14195 22247 14201
rect 22189 14161 22201 14195
rect 22235 14192 22247 14195
rect 22278 14192 22284 14204
rect 22235 14164 22284 14192
rect 22235 14161 22247 14164
rect 22189 14155 22247 14161
rect 22278 14152 22284 14164
rect 22336 14152 22342 14204
rect 19886 14124 19892 14136
rect 19444 14096 19892 14124
rect 19886 14084 19892 14096
rect 19944 14084 19950 14136
rect 22373 14059 22431 14065
rect 22373 14025 22385 14059
rect 22419 14056 22431 14059
rect 23109 14059 23167 14065
rect 23109 14056 23121 14059
rect 22419 14028 23121 14056
rect 22419 14025 22431 14028
rect 22373 14019 22431 14025
rect 23109 14025 23121 14028
rect 23155 14025 23167 14059
rect 23109 14019 23167 14025
rect 20073 13991 20131 13997
rect 20073 13988 20085 13991
rect 19352 13960 20085 13988
rect 20073 13957 20085 13960
rect 20119 13988 20131 13991
rect 22922 13988 22928 14000
rect 20119 13960 22928 13988
rect 20119 13957 20131 13960
rect 20073 13951 20131 13957
rect 22922 13948 22928 13960
rect 22980 13948 22986 14000
rect 5796 13824 23000 13920
rect 6181 13787 6239 13793
rect 6181 13784 6193 13787
rect 5736 13756 6193 13784
rect 6181 13753 6193 13756
rect 6227 13753 6239 13787
rect 6181 13747 6239 13753
rect 6641 13787 6699 13793
rect 6641 13753 6653 13787
rect 6687 13784 6699 13787
rect 6730 13784 6736 13796
rect 6687 13756 6736 13784
rect 6687 13753 6699 13756
rect 6641 13747 6699 13753
rect 6730 13744 6736 13756
rect 6788 13744 6794 13796
rect 7653 13787 7711 13793
rect 7653 13753 7665 13787
rect 7699 13784 7711 13787
rect 7926 13784 7932 13796
rect 7699 13756 7932 13784
rect 7699 13753 7711 13756
rect 7653 13747 7711 13753
rect 7926 13744 7932 13756
rect 7984 13744 7990 13796
rect 9030 13744 9036 13796
rect 9088 13784 9094 13796
rect 9309 13787 9367 13793
rect 9309 13784 9321 13787
rect 9088 13756 9321 13784
rect 9088 13744 9094 13756
rect 9309 13753 9321 13756
rect 9355 13753 9367 13787
rect 9309 13747 9367 13753
rect 11241 13787 11299 13793
rect 11241 13753 11253 13787
rect 11287 13784 11299 13787
rect 11330 13784 11336 13796
rect 11287 13756 11336 13784
rect 11287 13753 11299 13756
rect 11241 13747 11299 13753
rect 11330 13744 11336 13756
rect 11388 13744 11394 13796
rect 14366 13744 14372 13796
rect 14424 13784 14430 13796
rect 16209 13787 16267 13793
rect 16209 13784 16221 13787
rect 14424 13756 14596 13784
rect 14424 13744 14430 13756
rect 10226 13676 10232 13728
rect 10284 13716 10290 13728
rect 10344 13719 10402 13725
rect 10344 13716 10356 13719
rect 10284 13688 10356 13716
rect 10284 13676 10290 13688
rect 10344 13685 10356 13688
rect 10390 13685 10402 13719
rect 10344 13679 10402 13685
rect 10778 13676 10784 13728
rect 10836 13716 10842 13728
rect 12276 13719 12334 13725
rect 12276 13716 12288 13719
rect 10836 13688 12288 13716
rect 10836 13676 10842 13688
rect 12276 13685 12288 13688
rect 12322 13685 12334 13719
rect 12276 13679 12334 13685
rect 12805 13719 12863 13725
rect 12805 13685 12817 13719
rect 12851 13716 12863 13719
rect 13817 13719 13875 13725
rect 13817 13716 13829 13719
rect 12851 13688 13829 13716
rect 12851 13685 12863 13688
rect 12805 13679 12863 13685
rect 13817 13685 13829 13688
rect 13863 13685 13875 13719
rect 13817 13679 13875 13685
rect 12532 13660 12584 13666
rect 6362 13608 6368 13660
rect 6420 13648 6426 13660
rect 6733 13651 6791 13657
rect 6733 13648 6745 13651
rect 6420 13620 6745 13648
rect 6420 13608 6426 13620
rect 6733 13617 6745 13620
rect 6779 13617 6791 13651
rect 9122 13648 9128 13660
rect 6733 13611 6791 13617
rect 6840 13620 9128 13648
rect 6840 13589 6868 13620
rect 9122 13608 9128 13620
rect 9180 13648 9186 13660
rect 9180 13620 9591 13648
rect 12466 13620 12532 13648
rect 9180 13608 9186 13620
rect 12710 13608 12716 13660
rect 12768 13648 12774 13660
rect 12897 13651 12955 13657
rect 12897 13648 12909 13651
rect 12768 13620 12909 13648
rect 12768 13608 12774 13620
rect 12897 13617 12909 13620
rect 12943 13617 12955 13651
rect 14568 13648 14596 13756
rect 16040 13756 16221 13784
rect 16040 13648 16068 13756
rect 16209 13753 16221 13756
rect 16255 13753 16267 13787
rect 18322 13784 18328 13796
rect 18267 13756 18328 13784
rect 16209 13747 16267 13753
rect 18322 13744 18328 13756
rect 18380 13744 18386 13796
rect 20165 13787 20223 13793
rect 20165 13753 20177 13787
rect 20211 13784 20223 13787
rect 21726 13784 21732 13796
rect 20211 13756 21732 13784
rect 20211 13753 20223 13756
rect 20165 13747 20223 13753
rect 21726 13744 21732 13756
rect 21784 13744 21790 13796
rect 20257 13719 20315 13725
rect 20257 13716 20269 13719
rect 19812 13688 20269 13716
rect 18788 13660 18840 13666
rect 14568 13620 16068 13648
rect 17589 13651 17647 13657
rect 12897 13611 12955 13617
rect 17589 13617 17601 13651
rect 17635 13648 17647 13651
rect 17954 13648 17960 13660
rect 17635 13620 17960 13648
rect 17635 13617 17647 13620
rect 17589 13611 17647 13617
rect 17954 13608 17960 13620
rect 18012 13608 18018 13660
rect 18785 13648 18788 13657
rect 18724 13620 18788 13648
rect 18785 13611 18788 13620
rect 18840 13611 18843 13657
rect 12532 13602 12584 13608
rect 18788 13602 18840 13608
rect 6457 13583 6515 13589
rect 6457 13549 6469 13583
rect 6503 13549 6515 13583
rect 6457 13543 6515 13549
rect 6825 13583 6883 13589
rect 6825 13549 6837 13583
rect 6871 13549 6883 13583
rect 6825 13543 6883 13549
rect 6178 13404 6184 13456
rect 6236 13444 6242 13456
rect 6472 13444 6500 13543
rect 6730 13472 6736 13524
rect 6788 13512 6794 13524
rect 6840 13512 6868 13543
rect 6914 13540 6920 13592
rect 6972 13580 6978 13592
rect 7009 13583 7067 13589
rect 7009 13580 7021 13583
rect 6972 13552 7021 13580
rect 6972 13540 6978 13552
rect 7009 13549 7021 13552
rect 7055 13549 7067 13583
rect 7009 13543 7067 13549
rect 7469 13583 7527 13589
rect 7469 13549 7481 13583
rect 7515 13549 7527 13583
rect 7469 13543 7527 13549
rect 6788 13484 6868 13512
rect 6788 13472 6794 13484
rect 7484 13444 7512 13543
rect 9490 13540 9496 13592
rect 9548 13540 9554 13592
rect 10962 13540 10968 13592
rect 11020 13580 11026 13592
rect 13081 13583 13139 13589
rect 13081 13580 13093 13583
rect 11020 13552 11454 13580
rect 12636 13552 13093 13580
rect 11020 13540 11026 13552
rect 10686 13444 10692 13456
rect 6236 13416 7512 13444
rect 10631 13416 10692 13444
rect 6236 13404 6242 13416
rect 10686 13404 10692 13416
rect 10744 13404 10750 13456
rect 11606 13404 11612 13456
rect 11664 13444 11670 13456
rect 12636 13444 12664 13552
rect 13081 13549 13093 13552
rect 13127 13580 13139 13583
rect 13354 13580 13360 13592
rect 13127 13552 13360 13580
rect 13127 13549 13139 13552
rect 13081 13543 13139 13549
rect 13354 13540 13360 13552
rect 13412 13580 13418 13592
rect 14001 13583 14059 13589
rect 14001 13580 14013 13583
rect 13412 13552 14013 13580
rect 13412 13540 13418 13552
rect 14001 13549 14013 13552
rect 14047 13549 14059 13583
rect 14001 13543 14059 13549
rect 17770 13540 17776 13592
rect 17828 13580 17834 13592
rect 18141 13583 18199 13589
rect 18141 13580 18153 13583
rect 17828 13552 18153 13580
rect 17828 13540 17834 13552
rect 18141 13549 18153 13552
rect 18187 13549 18199 13583
rect 18141 13543 18199 13549
rect 17126 13472 17132 13524
rect 17184 13512 17190 13524
rect 17328 13515 17386 13521
rect 17328 13512 17340 13515
rect 17184 13484 17340 13512
rect 17184 13472 17190 13484
rect 17328 13481 17340 13484
rect 17374 13481 17386 13515
rect 17328 13475 17386 13481
rect 19046 13515 19104 13521
rect 19046 13481 19058 13515
rect 19092 13512 19104 13515
rect 19812 13512 19840 13688
rect 20257 13685 20269 13688
rect 20303 13685 20315 13719
rect 20257 13679 20315 13685
rect 21361 13719 21419 13725
rect 21361 13685 21373 13719
rect 21407 13685 21419 13719
rect 19886 13608 19892 13660
rect 19944 13648 19950 13660
rect 20456 13654 20944 13682
rect 21361 13679 21419 13685
rect 20456 13648 20484 13654
rect 19944 13620 20484 13648
rect 20916 13648 20944 13654
rect 21376 13648 21404 13679
rect 22744 13660 22796 13666
rect 22741 13648 22744 13657
rect 20916 13620 21404 13648
rect 22680 13620 22744 13648
rect 19944 13608 19950 13620
rect 22741 13611 22744 13620
rect 22796 13611 22799 13657
rect 22744 13602 22796 13608
rect 20438 13580 20444 13592
rect 20383 13552 20444 13580
rect 20438 13540 20444 13552
rect 20496 13540 20502 13592
rect 20714 13540 20720 13592
rect 20772 13580 20778 13592
rect 20809 13583 20867 13589
rect 20809 13580 20821 13583
rect 20772 13552 20821 13580
rect 20772 13540 20778 13552
rect 20809 13549 20821 13552
rect 20855 13549 20867 13583
rect 22462 13580 22468 13592
rect 22520 13589 22526 13592
rect 22520 13583 22538 13589
rect 22419 13552 22468 13580
rect 20809 13543 20867 13549
rect 22462 13540 22468 13552
rect 22526 13549 22538 13583
rect 22520 13543 22538 13549
rect 22520 13540 22526 13543
rect 20530 13512 20536 13524
rect 19092 13484 19840 13512
rect 20475 13484 20536 13512
rect 19092 13481 19104 13484
rect 19046 13475 19104 13481
rect 20530 13472 20536 13484
rect 20588 13472 20594 13524
rect 20625 13515 20683 13521
rect 20625 13481 20637 13515
rect 20671 13481 20683 13515
rect 20625 13475 20683 13481
rect 11664 13416 12664 13444
rect 11664 13404 11670 13416
rect 12986 13404 12992 13456
rect 13044 13444 13050 13456
rect 13265 13447 13323 13453
rect 13265 13444 13277 13447
rect 13044 13416 13277 13444
rect 13044 13404 13050 13416
rect 13265 13413 13277 13416
rect 13311 13413 13323 13447
rect 13265 13407 13323 13413
rect 13446 13404 13452 13456
rect 13504 13444 13510 13456
rect 14185 13447 14243 13453
rect 14185 13444 14197 13447
rect 13504 13416 14197 13444
rect 13504 13404 13510 13416
rect 14185 13413 14197 13416
rect 14231 13413 14243 13447
rect 14185 13407 14243 13413
rect 20162 13404 20168 13456
rect 20220 13444 20226 13456
rect 20640 13444 20668 13475
rect 20220 13416 20668 13444
rect 20220 13404 20226 13416
rect 5796 13280 23000 13376
rect 6641 13243 6699 13249
rect 6641 13209 6653 13243
rect 6687 13240 6699 13243
rect 6914 13240 6920 13252
rect 6687 13212 6920 13240
rect 6687 13209 6699 13212
rect 6641 13203 6699 13209
rect 6914 13200 6920 13212
rect 6972 13200 6978 13252
rect 8665 13243 8723 13249
rect 8665 13209 8677 13243
rect 8711 13240 8723 13243
rect 9490 13240 9496 13252
rect 8711 13212 8892 13240
rect 8711 13209 8723 13212
rect 8665 13203 8723 13209
rect 8864 13172 8892 13212
rect 9324 13212 9496 13240
rect 9324 13172 9352 13212
rect 9490 13200 9496 13212
rect 9548 13240 9554 13252
rect 9548 13212 9720 13240
rect 9548 13200 9554 13212
rect 9692 13206 9720 13212
rect 10428 13212 10916 13240
rect 10428 13206 10456 13212
rect 9692 13178 10456 13206
rect 7760 13144 8432 13172
rect 8864 13144 9352 13172
rect 10597 13175 10655 13181
rect 6362 13064 6368 13116
rect 6420 13104 6426 13116
rect 6549 13107 6607 13113
rect 6549 13104 6561 13107
rect 6420 13076 6561 13104
rect 6420 13064 6426 13076
rect 6549 13073 6561 13076
rect 6595 13073 6607 13107
rect 6730 13104 6736 13116
rect 6675 13076 6736 13104
rect 6549 13067 6607 13073
rect 6730 13064 6736 13076
rect 6788 13064 6794 13116
rect 7546 13107 7604 13113
rect 7546 13073 7558 13107
rect 7592 13104 7604 13107
rect 7760 13104 7788 13144
rect 7592 13076 7788 13104
rect 8404 13104 8432 13144
rect 10597 13141 10609 13175
rect 10643 13172 10655 13175
rect 10778 13172 10784 13184
rect 10643 13144 10784 13172
rect 10643 13141 10655 13144
rect 10597 13135 10655 13141
rect 10778 13132 10784 13144
rect 10836 13132 10842 13184
rect 10045 13107 10103 13113
rect 10045 13104 10057 13107
rect 8404 13076 8616 13104
rect 7592 13073 7604 13076
rect 7546 13067 7604 13073
rect 7282 13036 7288 13048
rect 7227 13008 7288 13036
rect 7282 12996 7288 13008
rect 7340 12996 7346 13048
rect 8588 13036 8616 13076
rect 9876 13076 10057 13104
rect 9876 13036 9904 13076
rect 10045 13073 10057 13076
rect 10091 13073 10103 13107
rect 10888 13090 10916 13212
rect 12526 13200 12532 13252
rect 12584 13240 12590 13252
rect 14185 13243 14243 13249
rect 14185 13240 14197 13243
rect 12584 13212 14197 13240
rect 12584 13200 12590 13212
rect 14185 13209 14197 13212
rect 14231 13209 14243 13243
rect 14185 13203 14243 13209
rect 15933 13243 15991 13249
rect 15933 13209 15945 13243
rect 15979 13240 15991 13243
rect 16022 13240 16028 13252
rect 15979 13212 16028 13240
rect 15979 13209 15991 13212
rect 15933 13203 15991 13209
rect 16022 13200 16028 13212
rect 16080 13200 16086 13252
rect 17310 13200 17316 13252
rect 17368 13240 17374 13252
rect 20073 13243 20131 13249
rect 17368 13212 17448 13240
rect 17368 13200 17374 13212
rect 12161 13175 12219 13181
rect 12161 13141 12173 13175
rect 12207 13172 12219 13175
rect 12710 13172 12716 13184
rect 12207 13144 12716 13172
rect 12207 13141 12219 13144
rect 12161 13135 12219 13141
rect 12710 13132 12716 13144
rect 12768 13132 12774 13184
rect 13066 13175 13124 13181
rect 13066 13141 13078 13175
rect 13112 13172 13124 13175
rect 13446 13172 13452 13184
rect 13112 13144 13452 13172
rect 13112 13141 13124 13144
rect 13066 13135 13124 13141
rect 13446 13132 13452 13144
rect 13504 13132 13510 13184
rect 14550 13132 14556 13184
rect 14608 13172 14614 13184
rect 15381 13175 15439 13181
rect 15381 13172 15393 13175
rect 14608 13144 15393 13172
rect 14608 13132 14614 13144
rect 15381 13141 15393 13144
rect 15427 13141 15439 13175
rect 15381 13135 15439 13141
rect 15473 13175 15531 13181
rect 15473 13141 15485 13175
rect 15519 13172 15531 13175
rect 16114 13172 16120 13184
rect 15519 13144 16120 13172
rect 15519 13141 15531 13144
rect 15473 13135 15531 13141
rect 16114 13132 16120 13144
rect 16172 13132 16178 13184
rect 17420 13172 17448 13212
rect 20073 13209 20085 13243
rect 20119 13240 20131 13243
rect 20530 13240 20536 13252
rect 20119 13212 20536 13240
rect 20119 13209 20131 13212
rect 20073 13203 20131 13209
rect 20530 13200 20536 13212
rect 20588 13200 20594 13252
rect 21726 13200 21732 13252
rect 21784 13240 21790 13252
rect 21784 13212 21956 13240
rect 21784 13200 21790 13212
rect 18616 13175 18674 13181
rect 18616 13172 18628 13175
rect 17420 13144 18628 13172
rect 18616 13141 18628 13144
rect 18662 13141 18674 13175
rect 18616 13135 18674 13141
rect 21200 13175 21258 13181
rect 21200 13141 21212 13175
rect 21246 13172 21258 13175
rect 21634 13172 21640 13184
rect 21246 13144 21640 13172
rect 21246 13141 21258 13144
rect 21200 13135 21258 13141
rect 21634 13132 21640 13144
rect 21692 13132 21698 13184
rect 21928 13181 21956 13212
rect 21913 13175 21971 13181
rect 21913 13141 21925 13175
rect 21959 13141 21971 13175
rect 21913 13135 21971 13141
rect 10045 13067 10103 13073
rect 13354 13064 13360 13116
rect 13412 13104 13418 13116
rect 15286 13104 15292 13116
rect 13412 13076 13860 13104
rect 15231 13076 15292 13104
rect 13412 13064 13418 13076
rect 11980 13048 12032 13054
rect 10229 13039 10287 13045
rect 10229 13036 10241 13039
rect 8588 13008 9904 13036
rect 10060 13008 10241 13036
rect 10060 12980 10088 13008
rect 10229 13005 10241 13008
rect 10275 13005 10287 13039
rect 10229 12999 10287 13005
rect 10413 13039 10471 13045
rect 10413 13005 10425 13039
rect 10459 13036 10471 13039
rect 10686 13036 10692 13048
rect 10459 13008 10692 13036
rect 10459 13005 10471 13008
rect 10413 12999 10471 13005
rect 10686 12996 10692 13008
rect 10744 12996 10750 13048
rect 11914 13008 11980 13036
rect 12342 12996 12348 13048
rect 12400 13036 12406 13048
rect 12805 13039 12863 13045
rect 12805 13036 12817 13039
rect 12400 13008 12817 13036
rect 12400 12996 12406 13008
rect 12805 13005 12817 13008
rect 12851 13005 12863 13039
rect 13832 13036 13860 13076
rect 15286 13064 15292 13076
rect 15344 13064 15350 13116
rect 15562 13064 15568 13116
rect 15620 13104 15626 13116
rect 15657 13107 15715 13113
rect 15657 13104 15669 13107
rect 15620 13076 15669 13104
rect 15620 13064 15626 13076
rect 15657 13073 15669 13076
rect 15703 13073 15715 13107
rect 15657 13067 15715 13073
rect 17052 13107 17110 13113
rect 17052 13073 17064 13107
rect 17098 13104 17110 13107
rect 17218 13104 17224 13116
rect 17098 13076 17224 13104
rect 17098 13073 17110 13076
rect 17052 13067 17110 13073
rect 17218 13064 17224 13076
rect 17276 13064 17282 13116
rect 17313 13107 17371 13113
rect 17313 13073 17325 13107
rect 17359 13104 17371 13107
rect 17494 13104 17500 13116
rect 17359 13076 17500 13104
rect 17359 13073 17371 13076
rect 17313 13067 17371 13073
rect 17494 13064 17500 13076
rect 17552 13064 17558 13116
rect 18782 13064 18788 13116
rect 18840 13104 18846 13116
rect 18877 13107 18935 13113
rect 18877 13104 18889 13107
rect 18840 13076 18889 13104
rect 18840 13064 18846 13076
rect 18877 13073 18889 13076
rect 18923 13073 18935 13107
rect 18877 13067 18935 13073
rect 20438 13064 20444 13116
rect 20496 13104 20502 13116
rect 21729 13107 21787 13113
rect 21729 13104 21741 13107
rect 20496 13076 21741 13104
rect 20496 13064 20502 13076
rect 21729 13073 21741 13076
rect 21775 13073 21787 13107
rect 21729 13067 21787 13073
rect 21818 13064 21824 13116
rect 21876 13104 21882 13116
rect 21876 13076 21937 13104
rect 21876 13064 21882 13076
rect 22002 13064 22008 13116
rect 22060 13104 22066 13116
rect 22097 13107 22155 13113
rect 22097 13104 22109 13107
rect 22060 13076 22109 13104
rect 22060 13064 22066 13076
rect 22097 13073 22109 13076
rect 22143 13073 22155 13107
rect 22097 13067 22155 13073
rect 14737 13039 14795 13045
rect 14737 13036 14749 13039
rect 13832 13008 14749 13036
rect 12805 12999 12863 13005
rect 14737 13005 14749 13008
rect 14783 13005 14795 13039
rect 21450 13036 21456 13048
rect 21395 13008 21456 13036
rect 14737 12999 14795 13005
rect 11980 12990 12032 12996
rect 10042 12928 10048 12980
rect 10100 12928 10106 12980
rect 10778 12928 10784 12980
rect 10836 12968 10842 12980
rect 11724 12971 11782 12977
rect 11724 12968 11736 12971
rect 10836 12940 11736 12968
rect 10836 12928 10842 12940
rect 11724 12937 11736 12940
rect 11770 12937 11782 12971
rect 14752 12968 14780 12999
rect 14936 12974 15792 13002
rect 21450 12996 21456 13008
rect 21508 12996 21514 13048
rect 14936 12968 14964 12974
rect 14752 12940 14964 12968
rect 15764 12968 15792 12974
rect 15764 12940 16436 12968
rect 11724 12931 11782 12937
rect 15105 12903 15163 12909
rect 15105 12869 15117 12903
rect 15151 12900 15163 12903
rect 15654 12900 15660 12912
rect 15151 12872 15660 12900
rect 15151 12869 15163 12872
rect 15105 12863 15163 12869
rect 15654 12860 15660 12872
rect 15712 12860 15718 12912
rect 16408 12900 16436 12940
rect 17034 12900 17040 12912
rect 16408 12872 17040 12900
rect 17034 12860 17040 12872
rect 17092 12860 17098 12912
rect 17494 12900 17500 12912
rect 17439 12872 17500 12900
rect 17494 12860 17500 12872
rect 17552 12860 17558 12912
rect 20162 12860 20168 12912
rect 20220 12900 20226 12912
rect 21545 12903 21603 12909
rect 21545 12900 21557 12903
rect 20220 12872 21557 12900
rect 20220 12860 20226 12872
rect 21545 12869 21557 12872
rect 21591 12869 21603 12903
rect 21545 12863 21603 12869
rect 5796 12736 23000 12832
rect 8757 12699 8815 12705
rect 8757 12665 8769 12699
rect 8803 12696 8815 12699
rect 10226 12696 10232 12708
rect 8803 12668 8984 12696
rect 8803 12665 8815 12668
rect 8757 12659 8815 12665
rect 8956 12662 8984 12668
rect 9600 12668 10232 12696
rect 9600 12662 9628 12668
rect 8956 12634 9628 12662
rect 10226 12656 10232 12668
rect 10284 12656 10290 12708
rect 11885 12699 11943 12705
rect 11885 12665 11897 12699
rect 11931 12696 11943 12699
rect 11974 12696 11980 12708
rect 11931 12668 11980 12696
rect 11931 12665 11943 12668
rect 11885 12659 11943 12665
rect 11974 12656 11980 12668
rect 12032 12696 12038 12708
rect 12032 12668 13676 12696
rect 12032 12656 12038 12668
rect 9792 12631 9850 12637
rect 9792 12597 9804 12631
rect 9838 12628 9850 12631
rect 10410 12628 10416 12640
rect 9838 12600 10416 12628
rect 9838 12597 9850 12600
rect 9792 12591 9850 12597
rect 10410 12588 10416 12600
rect 10468 12588 10474 12640
rect 7926 12560 7932 12572
rect 7484 12532 7932 12560
rect 6365 12495 6423 12501
rect 6365 12461 6377 12495
rect 6411 12492 6423 12495
rect 6411 12464 6500 12492
rect 6411 12461 6423 12464
rect 6365 12455 6423 12461
rect 6472 12424 6500 12464
rect 6546 12452 6552 12504
rect 6604 12492 6610 12504
rect 7101 12495 7159 12501
rect 6604 12464 6665 12492
rect 6604 12452 6610 12464
rect 7101 12461 7113 12495
rect 7147 12492 7159 12495
rect 7484 12492 7512 12532
rect 7926 12520 7932 12532
rect 7984 12560 7990 12572
rect 13262 12560 13268 12572
rect 7984 12532 9062 12560
rect 13207 12532 13268 12560
rect 7984 12520 7990 12532
rect 13262 12520 13268 12532
rect 13320 12520 13326 12572
rect 13648 12560 13676 12668
rect 16758 12656 16764 12708
rect 16816 12696 16822 12708
rect 17126 12696 17132 12708
rect 16816 12668 16988 12696
rect 17071 12668 17132 12696
rect 16816 12656 16822 12668
rect 16040 12600 16620 12628
rect 13648 12532 13768 12560
rect 7147 12464 7512 12492
rect 7147 12461 7159 12464
rect 7101 12455 7159 12461
rect 8846 12452 8852 12504
rect 8904 12492 8910 12504
rect 12986 12492 12992 12504
rect 13044 12501 13050 12504
rect 13044 12495 13062 12501
rect 8904 12464 8970 12492
rect 12943 12464 12992 12492
rect 8904 12452 8910 12464
rect 12986 12452 12992 12464
rect 13050 12461 13062 12495
rect 13044 12455 13062 12461
rect 13044 12452 13050 12455
rect 13446 12452 13452 12504
rect 13504 12492 13510 12504
rect 13633 12495 13691 12501
rect 13633 12492 13645 12495
rect 13504 12464 13645 12492
rect 13504 12452 13510 12464
rect 13633 12461 13645 12464
rect 13679 12461 13691 12495
rect 13740 12492 13768 12532
rect 15838 12520 15844 12572
rect 15896 12560 15902 12572
rect 16040 12560 16068 12600
rect 15896 12532 16068 12560
rect 16592 12560 16620 12600
rect 16592 12532 16896 12560
rect 15896 12520 15902 12532
rect 13894 12495 13952 12501
rect 13894 12492 13906 12495
rect 13740 12464 13906 12492
rect 13633 12455 13691 12461
rect 13894 12461 13906 12464
rect 13940 12461 13952 12495
rect 13894 12455 13952 12461
rect 15562 12452 15568 12504
rect 15620 12492 15626 12504
rect 16577 12495 16635 12501
rect 16577 12492 16589 12495
rect 15620 12464 16589 12492
rect 15620 12452 15626 12464
rect 16577 12461 16589 12464
rect 16623 12461 16635 12495
rect 16577 12455 16635 12461
rect 16758 12452 16764 12504
rect 16816 12452 16822 12504
rect 16868 12501 16896 12532
rect 16960 12501 16988 12668
rect 17126 12656 17132 12668
rect 17184 12656 17190 12708
rect 21634 12656 21640 12708
rect 21692 12696 21698 12708
rect 22741 12699 22799 12705
rect 22741 12696 22753 12699
rect 21692 12668 22753 12696
rect 21692 12656 21698 12668
rect 22741 12665 22753 12668
rect 22787 12696 22799 12699
rect 22922 12696 22928 12708
rect 22787 12668 22928 12696
rect 22787 12665 22799 12668
rect 22741 12659 22799 12665
rect 22922 12656 22928 12668
rect 22980 12656 22986 12708
rect 18601 12563 18659 12569
rect 18601 12529 18613 12563
rect 18647 12560 18659 12563
rect 18782 12560 18788 12572
rect 18647 12532 18788 12560
rect 18647 12529 18659 12532
rect 18601 12523 18659 12529
rect 18782 12520 18788 12532
rect 18840 12520 18846 12572
rect 16853 12495 16911 12501
rect 16853 12461 16865 12495
rect 16899 12461 16911 12495
rect 16853 12455 16911 12461
rect 16945 12495 17003 12501
rect 16945 12461 16957 12495
rect 16991 12492 17003 12495
rect 17126 12492 17132 12504
rect 16991 12464 17132 12492
rect 16991 12461 17003 12464
rect 16945 12455 17003 12461
rect 17126 12452 17132 12464
rect 17184 12452 17190 12504
rect 20162 12492 20168 12504
rect 19168 12464 19932 12492
rect 20107 12464 20168 12492
rect 6730 12424 6736 12436
rect 6472 12396 6736 12424
rect 6730 12384 6736 12396
rect 6788 12424 6794 12436
rect 6917 12427 6975 12433
rect 6917 12424 6929 12427
rect 6788 12396 6929 12424
rect 6788 12384 6794 12396
rect 6917 12393 6929 12396
rect 6963 12393 6975 12427
rect 6917 12387 6975 12393
rect 18340 12427 18398 12433
rect 18340 12393 18352 12427
rect 18386 12424 18398 12427
rect 18966 12424 18972 12436
rect 18386 12396 18972 12424
rect 18386 12393 18398 12396
rect 6362 12356 6368 12368
rect 5736 12328 6368 12356
rect 5736 12152 5764 12328
rect 6362 12316 6368 12328
rect 6420 12356 6426 12368
rect 6457 12359 6515 12365
rect 6457 12356 6469 12359
rect 6420 12328 6469 12356
rect 6420 12316 6426 12328
rect 6457 12325 6469 12328
rect 6503 12325 6515 12359
rect 6457 12319 6515 12325
rect 10137 12359 10195 12365
rect 10137 12325 10149 12359
rect 10183 12356 10195 12359
rect 10226 12356 10232 12368
rect 10183 12328 10232 12356
rect 10183 12325 10195 12328
rect 10137 12319 10195 12325
rect 10226 12316 10232 12328
rect 10284 12316 10290 12368
rect 15013 12359 15071 12365
rect 15013 12325 15025 12359
rect 15059 12356 15071 12359
rect 15212 12362 16620 12390
rect 18340 12387 18398 12393
rect 18966 12384 18972 12396
rect 19024 12384 19030 12436
rect 15212 12356 15240 12362
rect 15059 12328 15240 12356
rect 16592 12356 16620 12362
rect 16758 12356 16764 12368
rect 16592 12328 16764 12356
rect 15059 12325 15071 12328
rect 15013 12319 15071 12325
rect 16758 12316 16764 12328
rect 16816 12316 16822 12368
rect 17221 12359 17279 12365
rect 17221 12325 17233 12359
rect 17267 12356 17279 12359
rect 17954 12356 17960 12368
rect 17267 12328 17960 12356
rect 17267 12325 17279 12328
rect 17221 12319 17279 12325
rect 17954 12316 17960 12328
rect 18012 12356 18018 12368
rect 19168 12356 19196 12464
rect 19904 12390 19932 12464
rect 20162 12452 20168 12464
rect 20220 12452 20226 12504
rect 21082 12492 21088 12504
rect 21027 12464 21088 12492
rect 21082 12452 21088 12464
rect 21140 12492 21146 12504
rect 21361 12495 21419 12501
rect 21361 12492 21373 12495
rect 21140 12464 21373 12492
rect 21140 12452 21146 12464
rect 21361 12461 21373 12464
rect 21407 12461 21419 12495
rect 21361 12455 21419 12461
rect 22480 12464 23060 12492
rect 21634 12433 21640 12436
rect 21622 12427 21640 12433
rect 21622 12424 21634 12427
rect 21579 12396 21634 12424
rect 21622 12393 21634 12396
rect 19904 12362 20944 12390
rect 21622 12387 21640 12393
rect 21634 12384 21640 12387
rect 21692 12384 21698 12436
rect 22480 12424 22508 12464
rect 21836 12396 22508 12424
rect 18012 12328 19196 12356
rect 20916 12356 20944 12362
rect 21836 12356 21864 12396
rect 20916 12328 21864 12356
rect 23032 12356 23060 12464
rect 28718 12356 28724 12368
rect 23032 12328 28724 12356
rect 18012 12316 18018 12328
rect 28718 12316 28724 12328
rect 28776 12316 28782 12368
rect 5796 12192 23000 12288
rect 6273 12155 6331 12161
rect 6273 12152 6285 12155
rect 5736 12124 6285 12152
rect 6273 12121 6285 12124
rect 6319 12121 6331 12155
rect 6273 12115 6331 12121
rect 6549 12155 6607 12161
rect 6549 12121 6561 12155
rect 6595 12152 6607 12155
rect 6730 12152 6736 12164
rect 6595 12124 6736 12152
rect 6595 12121 6607 12124
rect 6549 12115 6607 12121
rect 6730 12112 6736 12124
rect 6788 12112 6794 12164
rect 8846 12152 8852 12164
rect 8791 12124 8852 12152
rect 8846 12112 8852 12124
rect 8904 12152 8910 12164
rect 8904 12124 9076 12152
rect 8904 12112 8910 12124
rect 9048 12084 9076 12124
rect 10428 12124 10916 12152
rect 10428 12118 10456 12124
rect 9508 12090 10456 12118
rect 9508 12084 9536 12090
rect 7944 12056 8524 12084
rect 9048 12056 9536 12084
rect 10597 12087 10655 12093
rect 6546 11976 6552 12028
rect 6604 12016 6610 12028
rect 6641 12019 6699 12025
rect 6641 12016 6653 12019
rect 6604 11988 6653 12016
rect 6604 11976 6610 11988
rect 6641 11985 6653 11988
rect 6687 11985 6699 12019
rect 6641 11979 6699 11985
rect 7730 12019 7788 12025
rect 7730 11985 7742 12019
rect 7776 12016 7788 12019
rect 7944 12016 7972 12056
rect 7776 11988 7972 12016
rect 8496 12016 8524 12056
rect 10597 12053 10609 12087
rect 10643 12084 10655 12087
rect 10778 12084 10784 12096
rect 10643 12056 10784 12084
rect 10643 12053 10655 12056
rect 10597 12047 10655 12053
rect 10778 12044 10784 12056
rect 10836 12044 10842 12096
rect 9861 12019 9919 12025
rect 9861 12016 9873 12019
rect 8496 11988 8708 12016
rect 7776 11985 7788 11988
rect 7730 11979 7788 11985
rect 7282 11908 7288 11960
rect 7340 11948 7346 11960
rect 7469 11951 7527 11957
rect 7469 11948 7481 11951
rect 7340 11920 7481 11948
rect 7340 11908 7346 11920
rect 7469 11917 7481 11920
rect 7515 11917 7527 11951
rect 8680 11948 8708 11988
rect 9692 11988 9873 12016
rect 9692 11948 9720 11988
rect 9861 11985 9873 11988
rect 9907 11985 9919 12019
rect 10888 12002 10916 12124
rect 14550 12112 14556 12164
rect 14608 12152 14614 12164
rect 14737 12155 14795 12161
rect 14737 12152 14749 12155
rect 14608 12124 14749 12152
rect 14608 12112 14614 12124
rect 14737 12121 14749 12124
rect 14783 12121 14795 12155
rect 14737 12115 14795 12121
rect 16758 12112 16764 12164
rect 16816 12152 16822 12164
rect 21545 12155 21603 12161
rect 16816 12124 17080 12152
rect 16816 12112 16822 12124
rect 13262 12084 13268 12096
rect 11900 12056 12296 12084
rect 9861 11979 9919 11985
rect 10042 11948 10048 11960
rect 8680 11920 9720 11948
rect 9987 11920 10048 11948
rect 7469 11911 7527 11917
rect 10042 11908 10048 11920
rect 10100 11908 10106 11960
rect 10226 11948 10232 11960
rect 10171 11920 10232 11948
rect 10226 11908 10232 11920
rect 10284 11908 10290 11960
rect 11900 11934 11928 12056
rect 12268 12016 12296 12056
rect 13096 12056 13268 12084
rect 13096 12016 13124 12056
rect 13262 12044 13268 12056
rect 13320 12084 13326 12096
rect 13618 12087 13676 12093
rect 13618 12084 13630 12087
rect 13320 12056 13630 12084
rect 13320 12044 13326 12056
rect 13618 12053 13630 12056
rect 13664 12053 13676 12087
rect 13618 12047 13676 12053
rect 15182 12087 15240 12093
rect 15182 12053 15194 12087
rect 15228 12084 15240 12087
rect 15654 12084 15660 12096
rect 15228 12056 15660 12084
rect 15228 12053 15240 12056
rect 15182 12047 15240 12053
rect 15654 12044 15660 12056
rect 15712 12044 15718 12096
rect 17052 12093 17080 12124
rect 21545 12121 21557 12155
rect 21591 12152 21603 12155
rect 21634 12152 21640 12164
rect 21591 12124 21640 12152
rect 21591 12121 21603 12124
rect 21545 12115 21603 12121
rect 21634 12112 21640 12124
rect 21692 12112 21698 12164
rect 16393 12087 16451 12093
rect 16393 12053 16405 12087
rect 16439 12084 16451 12087
rect 16945 12087 17003 12093
rect 16945 12084 16957 12087
rect 16439 12056 16957 12084
rect 16439 12053 16451 12056
rect 16393 12047 16451 12053
rect 16945 12053 16957 12056
rect 16991 12053 17003 12087
rect 16945 12047 17003 12053
rect 17037 12087 17095 12093
rect 17037 12053 17049 12087
rect 17083 12053 17095 12087
rect 17037 12047 17095 12053
rect 17494 12044 17500 12096
rect 17552 12084 17558 12096
rect 17865 12087 17923 12093
rect 17865 12084 17877 12087
rect 17552 12056 17877 12084
rect 17552 12044 17558 12056
rect 17865 12053 17877 12056
rect 17911 12053 17923 12087
rect 17865 12047 17923 12053
rect 17954 12044 17960 12096
rect 18012 12084 18018 12096
rect 18770 12087 18828 12093
rect 18012 12056 18073 12084
rect 18012 12044 18018 12056
rect 18770 12053 18782 12087
rect 18816 12084 18828 12087
rect 20070 12084 20076 12096
rect 18816 12056 20076 12084
rect 18816 12053 18828 12056
rect 18770 12047 18828 12053
rect 20070 12044 20076 12056
rect 20128 12044 20134 12096
rect 12268 11988 13124 12016
rect 13357 12019 13415 12025
rect 13357 11985 13369 12019
rect 13403 12016 13415 12019
rect 13446 12016 13452 12028
rect 13403 11988 13452 12016
rect 13403 11985 13415 11988
rect 13357 11979 13415 11985
rect 13446 11976 13452 11988
rect 13504 11976 13510 12028
rect 14921 12019 14979 12025
rect 14921 11985 14933 12019
rect 14967 12016 14979 12019
rect 15470 12016 15476 12028
rect 14967 11988 15476 12016
rect 14967 11985 14979 11988
rect 14921 11979 14979 11985
rect 15470 11976 15476 11988
rect 15528 11976 15534 12028
rect 15562 11976 15568 12028
rect 15620 12016 15626 12028
rect 16761 12019 16819 12025
rect 16761 12016 16773 12019
rect 15620 11988 16773 12016
rect 15620 11976 15626 11988
rect 11980 11960 12032 11966
rect 12069 11951 12127 11957
rect 12069 11948 12081 11951
rect 12032 11920 12081 11948
rect 12069 11917 12081 11920
rect 12115 11917 12127 11951
rect 12069 11911 12127 11917
rect 11980 11902 12032 11908
rect 10594 11840 10600 11892
rect 10652 11880 10658 11892
rect 11724 11883 11782 11889
rect 11724 11880 11736 11883
rect 10652 11852 10824 11880
rect 10652 11840 10658 11852
rect 10796 11846 10824 11852
rect 11532 11852 11736 11880
rect 11532 11846 11560 11852
rect 6362 11812 6368 11824
rect 6307 11784 6368 11812
rect 6362 11772 6368 11784
rect 6420 11772 6426 11824
rect 10796 11818 11560 11846
rect 11724 11849 11736 11852
rect 11770 11849 11782 11883
rect 16500 11880 16528 11988
rect 16761 11985 16773 11988
rect 16807 11985 16819 12019
rect 17126 12016 17132 12028
rect 17071 11988 17132 12016
rect 16761 11979 16819 11985
rect 17126 11976 17132 11988
rect 17184 12016 17190 12028
rect 17773 12019 17831 12025
rect 17773 12016 17785 12019
rect 17184 11988 17785 12016
rect 17184 11976 17190 11988
rect 17773 11985 17785 11988
rect 17819 11985 17831 12019
rect 17773 11979 17831 11985
rect 18141 12019 18199 12025
rect 18141 11985 18153 12019
rect 18187 11985 18199 12019
rect 21174 12016 21180 12028
rect 21232 12025 21238 12028
rect 21232 12019 21250 12025
rect 21131 11988 21180 12016
rect 18141 11979 18199 11985
rect 17310 11880 17316 11892
rect 16500 11852 16804 11880
rect 17255 11852 17316 11880
rect 11724 11843 11782 11849
rect 16776 11812 16804 11852
rect 17310 11840 17316 11852
rect 17368 11840 17374 11892
rect 18156 11880 18184 11979
rect 21174 11976 21180 11988
rect 21238 11985 21250 12019
rect 21232 11979 21250 11985
rect 21232 11976 21238 11979
rect 18506 11948 18512 11960
rect 18451 11920 18512 11948
rect 18506 11908 18512 11920
rect 18564 11908 18570 11960
rect 21450 11948 21456 11960
rect 21395 11920 21456 11948
rect 21450 11908 21456 11920
rect 21508 11908 21514 11960
rect 21729 11951 21787 11957
rect 21729 11917 21741 11951
rect 21775 11948 21787 11951
rect 22186 11948 22192 11960
rect 21775 11920 22192 11948
rect 21775 11917 21787 11920
rect 21729 11911 21787 11917
rect 22186 11908 22192 11920
rect 22244 11908 22250 11960
rect 22388 11920 23060 11948
rect 18230 11880 18236 11892
rect 17420 11852 18236 11880
rect 17420 11812 17448 11852
rect 18230 11840 18236 11852
rect 18288 11840 18294 11892
rect 21913 11883 21971 11889
rect 21913 11849 21925 11883
rect 21959 11880 21971 11883
rect 22388 11880 22416 11920
rect 21959 11852 22416 11880
rect 23032 11880 23060 11920
rect 23661 11883 23719 11889
rect 23661 11880 23673 11883
rect 23032 11852 23673 11880
rect 21959 11849 21971 11852
rect 21913 11843 21971 11849
rect 23661 11849 23673 11852
rect 23707 11849 23719 11883
rect 23661 11843 23719 11849
rect 17586 11812 17592 11824
rect 16776 11784 17448 11812
rect 17531 11784 17592 11812
rect 17586 11772 17592 11784
rect 17644 11772 17650 11824
rect 19889 11815 19947 11821
rect 19889 11781 19901 11815
rect 19935 11812 19947 11815
rect 19978 11812 19984 11824
rect 19935 11784 19984 11812
rect 19935 11781 19947 11784
rect 19889 11775 19947 11781
rect 19978 11772 19984 11784
rect 20036 11772 20042 11824
rect 20073 11815 20131 11821
rect 20073 11781 20085 11815
rect 20119 11812 20131 11815
rect 21726 11812 21732 11824
rect 20119 11784 21732 11812
rect 20119 11781 20131 11784
rect 20073 11775 20131 11781
rect 21726 11772 21732 11784
rect 21784 11772 21790 11824
rect 5796 11648 23000 11744
rect 7926 11568 7932 11620
rect 7984 11608 7990 11620
rect 8297 11611 8355 11617
rect 8297 11608 8309 11611
rect 7984 11580 8309 11608
rect 7984 11568 7990 11580
rect 8297 11577 8309 11580
rect 8343 11577 8355 11611
rect 8297 11571 8355 11577
rect 10410 11568 10416 11620
rect 10468 11608 10474 11620
rect 10597 11611 10655 11617
rect 10597 11608 10609 11611
rect 10468 11580 10609 11608
rect 10468 11568 10474 11580
rect 10597 11577 10609 11580
rect 10643 11577 10655 11611
rect 10597 11571 10655 11577
rect 13262 11568 13268 11620
rect 13320 11608 13326 11620
rect 13449 11611 13507 11617
rect 13449 11608 13461 11611
rect 13320 11580 13461 11608
rect 13320 11568 13326 11580
rect 13449 11577 13461 11580
rect 13495 11577 13507 11611
rect 13449 11571 13507 11577
rect 6362 11500 6368 11552
rect 6420 11540 6426 11552
rect 6457 11543 6515 11549
rect 6457 11540 6469 11543
rect 6420 11512 6469 11540
rect 6420 11500 6426 11512
rect 6457 11509 6469 11512
rect 6503 11509 6515 11543
rect 6457 11503 6515 11509
rect 8846 11500 8852 11552
rect 8904 11540 8910 11552
rect 9562 11543 9620 11549
rect 9562 11540 9574 11543
rect 8904 11512 9574 11540
rect 8904 11500 8910 11512
rect 9562 11509 9574 11512
rect 9608 11509 9620 11543
rect 9562 11503 9620 11509
rect 11425 11543 11483 11549
rect 11425 11509 11437 11543
rect 11471 11540 11483 11543
rect 11974 11540 11980 11552
rect 11471 11512 11980 11540
rect 11471 11509 11483 11512
rect 11425 11503 11483 11509
rect 11974 11500 11980 11512
rect 12032 11500 12038 11552
rect 20165 11543 20223 11549
rect 20165 11509 20177 11543
rect 20211 11540 20223 11543
rect 21634 11540 21640 11552
rect 20211 11512 21640 11540
rect 20211 11509 20223 11512
rect 20165 11503 20223 11509
rect 21634 11500 21640 11512
rect 21692 11500 21698 11552
rect 13998 11472 14004 11484
rect 6178 11364 6184 11416
rect 6236 11404 6242 11416
rect 6638 11404 6644 11416
rect 6236 11376 6644 11404
rect 6236 11364 6242 11376
rect 6638 11364 6644 11376
rect 6696 11364 6702 11416
rect 6917 11407 6975 11413
rect 6917 11373 6929 11407
rect 6963 11404 6975 11407
rect 7190 11404 7196 11416
rect 6963 11376 7196 11404
rect 6963 11373 6975 11376
rect 6917 11367 6975 11373
rect 7190 11364 7196 11376
rect 7248 11364 7254 11416
rect 8662 11364 8668 11416
rect 8720 11404 8726 11416
rect 9416 11404 9444 11458
rect 13943 11444 14004 11472
rect 13998 11432 14004 11444
rect 14056 11432 14062 11484
rect 22738 11472 22744 11484
rect 22683 11444 22744 11472
rect 22738 11432 22744 11444
rect 22796 11432 22802 11484
rect 10502 11404 10508 11416
rect 8720 11376 9444 11404
rect 10442 11376 10508 11404
rect 8720 11364 8726 11376
rect 10502 11364 10508 11376
rect 10560 11364 10566 11416
rect 11606 11404 11612 11416
rect 11551 11376 11612 11404
rect 11606 11364 11612 11376
rect 11664 11364 11670 11416
rect 12069 11407 12127 11413
rect 12069 11373 12081 11407
rect 12115 11404 12127 11407
rect 12342 11404 12348 11416
rect 12115 11376 12348 11404
rect 12115 11373 12127 11376
rect 12069 11367 12127 11373
rect 12342 11364 12348 11376
rect 12400 11364 12406 11416
rect 14262 11407 14320 11413
rect 14262 11373 14274 11407
rect 14308 11404 14320 11407
rect 14550 11404 14556 11416
rect 14308 11376 14556 11404
rect 14308 11373 14320 11376
rect 14262 11367 14320 11373
rect 14550 11364 14556 11376
rect 14608 11364 14614 11416
rect 15470 11404 15476 11416
rect 15415 11376 15476 11404
rect 15470 11364 15476 11376
rect 15528 11364 15534 11416
rect 15838 11404 15844 11416
rect 15783 11376 15844 11404
rect 15838 11364 15844 11376
rect 15896 11364 15902 11416
rect 16850 11404 16856 11416
rect 16795 11376 16856 11404
rect 16850 11364 16856 11376
rect 16908 11364 16914 11416
rect 17114 11407 17172 11413
rect 17114 11373 17126 11407
rect 17160 11404 17172 11407
rect 17586 11404 17592 11416
rect 17160 11376 17592 11404
rect 17160 11373 17172 11376
rect 17114 11367 17172 11373
rect 17586 11364 17592 11376
rect 17644 11364 17650 11416
rect 18782 11404 18788 11416
rect 18064 11376 18552 11404
rect 18727 11376 18788 11404
rect 6825 11339 6883 11345
rect 6825 11305 6837 11339
rect 6871 11336 6883 11339
rect 11793 11339 11851 11345
rect 6871 11330 7231 11336
rect 6871 11308 7185 11330
rect 6871 11305 6883 11308
rect 6825 11299 6883 11305
rect 7173 11296 7185 11308
rect 7219 11296 7231 11330
rect 11793 11305 11805 11339
rect 11839 11336 11851 11339
rect 15657 11339 15715 11345
rect 11839 11330 12383 11336
rect 11839 11308 12337 11330
rect 11839 11305 11851 11308
rect 11793 11299 11851 11305
rect 7173 11290 7231 11296
rect 12325 11296 12337 11308
rect 12371 11296 12383 11330
rect 15657 11305 15669 11339
rect 15703 11305 15715 11339
rect 15657 11299 15715 11305
rect 12325 11290 12383 11296
rect 9030 11228 9036 11280
rect 9088 11268 9094 11280
rect 9217 11271 9275 11277
rect 9217 11268 9229 11271
rect 9088 11240 9229 11268
rect 9088 11228 9094 11240
rect 9217 11237 9229 11240
rect 9263 11237 9275 11271
rect 9217 11231 9275 11237
rect 15381 11271 15439 11277
rect 15381 11237 15393 11271
rect 15427 11268 15439 11271
rect 15672 11268 15700 11299
rect 15746 11296 15752 11348
rect 15804 11336 15810 11348
rect 18064 11336 18092 11376
rect 15804 11308 15865 11336
rect 17880 11308 18092 11336
rect 18524 11336 18552 11376
rect 18782 11364 18788 11376
rect 18840 11364 18846 11416
rect 20625 11407 20683 11413
rect 20625 11404 20637 11407
rect 20456 11376 20637 11404
rect 20456 11348 20484 11376
rect 20625 11373 20637 11376
rect 20671 11373 20683 11407
rect 20625 11367 20683 11373
rect 20993 11407 21051 11413
rect 20993 11373 21005 11407
rect 21039 11404 21051 11407
rect 21174 11404 21180 11416
rect 21039 11376 21180 11404
rect 21039 11373 21051 11376
rect 20993 11367 21051 11373
rect 21174 11364 21180 11376
rect 21232 11364 21238 11416
rect 22480 11407 22538 11413
rect 22480 11373 22492 11407
rect 22526 11404 22538 11407
rect 23845 11407 23903 11413
rect 23845 11404 23857 11407
rect 22526 11376 23857 11404
rect 22526 11373 22538 11376
rect 22480 11367 22538 11373
rect 23845 11373 23857 11376
rect 23891 11373 23903 11407
rect 23845 11367 23903 11373
rect 19046 11339 19104 11345
rect 19046 11336 19058 11339
rect 18524 11308 19058 11336
rect 15804 11296 15810 11308
rect 15427 11240 15700 11268
rect 16209 11271 16267 11277
rect 15427 11237 15439 11240
rect 15381 11231 15439 11237
rect 16209 11237 16221 11271
rect 16255 11268 16267 11271
rect 16408 11274 17172 11302
rect 17880 11280 17908 11308
rect 19046 11305 19058 11308
rect 19092 11305 19104 11339
rect 19046 11299 19104 11305
rect 19150 11296 19156 11348
rect 19208 11336 19214 11348
rect 20349 11339 20407 11345
rect 20349 11336 20361 11339
rect 19208 11308 20361 11336
rect 19208 11296 19214 11308
rect 20349 11305 20361 11308
rect 20395 11305 20407 11339
rect 20349 11299 20407 11305
rect 20438 11296 20444 11348
rect 20496 11296 20502 11348
rect 20530 11296 20536 11348
rect 20588 11336 20594 11348
rect 20717 11339 20775 11345
rect 20717 11336 20729 11339
rect 20588 11308 20729 11336
rect 20588 11296 20594 11308
rect 20717 11305 20729 11308
rect 20763 11305 20775 11339
rect 20717 11299 20775 11305
rect 20806 11296 20812 11348
rect 20864 11336 20870 11348
rect 20864 11308 20925 11336
rect 20864 11296 20870 11308
rect 16408 11268 16436 11274
rect 16255 11240 16436 11268
rect 17144 11268 17172 11274
rect 17310 11268 17316 11280
rect 17144 11240 17316 11268
rect 16255 11237 16267 11240
rect 16209 11231 16267 11237
rect 17310 11228 17316 11240
rect 17368 11228 17374 11280
rect 17862 11228 17868 11280
rect 17920 11228 17926 11280
rect 18046 11228 18052 11280
rect 18104 11268 18110 11280
rect 18233 11271 18291 11277
rect 18233 11268 18245 11271
rect 18104 11240 18245 11268
rect 18104 11228 18110 11240
rect 18233 11237 18245 11240
rect 18279 11237 18291 11271
rect 21358 11268 21364 11280
rect 21303 11240 21364 11268
rect 18233 11231 18291 11237
rect 21358 11228 21364 11240
rect 21416 11228 21422 11280
rect 5796 11104 23000 11200
rect 11330 11024 11336 11076
rect 11388 11064 11394 11076
rect 11885 11067 11943 11073
rect 11885 11064 11897 11067
rect 11388 11036 11897 11064
rect 11388 11024 11394 11036
rect 11885 11033 11897 11036
rect 11931 11033 11943 11067
rect 11885 11027 11943 11033
rect 14737 11067 14795 11073
rect 14737 11033 14749 11067
rect 14783 11064 14795 11067
rect 15746 11064 15752 11076
rect 14783 11036 14964 11064
rect 14783 11033 14795 11036
rect 14737 11027 14795 11033
rect 10413 10999 10471 11005
rect 10413 10965 10425 10999
rect 10459 10996 10471 10999
rect 10594 10996 10600 11008
rect 10459 10968 10600 10996
rect 10459 10965 10471 10968
rect 10413 10959 10471 10965
rect 10594 10956 10600 10968
rect 10652 10956 10658 11008
rect 13618 10999 13676 11005
rect 13618 10996 13630 10999
rect 13280 10968 13630 10996
rect 6638 10888 6644 10940
rect 6696 10928 6702 10940
rect 6825 10931 6883 10937
rect 6825 10928 6837 10931
rect 6696 10900 6837 10928
rect 6696 10888 6702 10900
rect 6825 10897 6837 10900
rect 6871 10897 6883 10931
rect 6825 10891 6883 10897
rect 7009 10931 7067 10937
rect 7009 10897 7021 10931
rect 7055 10928 7067 10931
rect 7546 10931 7604 10937
rect 7546 10928 7558 10931
rect 7055 10900 7558 10928
rect 7055 10897 7067 10900
rect 7009 10891 7067 10897
rect 7546 10897 7558 10900
rect 7592 10897 7604 10931
rect 7546 10891 7604 10897
rect 9125 10931 9183 10937
rect 9125 10897 9137 10931
rect 9171 10928 9183 10931
rect 10042 10928 10048 10940
rect 9171 10900 10048 10928
rect 9171 10897 9183 10900
rect 9125 10891 9183 10897
rect 10042 10888 10048 10900
rect 10100 10888 10106 10940
rect 10502 10888 10508 10940
rect 10560 10928 10566 10940
rect 10560 10900 10718 10928
rect 10560 10888 10566 10900
rect 13280 10872 13308 10968
rect 13618 10965 13630 10968
rect 13664 10965 13676 10999
rect 14936 10996 14964 11036
rect 15488 11036 15752 11064
rect 15488 10996 15516 11036
rect 15746 11024 15752 11036
rect 15804 11024 15810 11076
rect 19705 11067 19763 11073
rect 19705 11033 19717 11067
rect 19751 11064 19763 11067
rect 20806 11064 20812 11076
rect 19751 11036 19932 11064
rect 19751 11033 19763 11036
rect 19705 11027 19763 11033
rect 19904 11030 19932 11036
rect 20640 11036 20812 11064
rect 20640 11030 20668 11036
rect 19904 11002 20668 11030
rect 20806 11024 20812 11036
rect 20864 11024 20870 11076
rect 14936 10968 15516 10996
rect 18800 10968 19380 10996
rect 13618 10959 13676 10965
rect 13357 10931 13415 10937
rect 13357 10897 13369 10931
rect 13403 10928 13415 10931
rect 13446 10928 13452 10940
rect 13403 10900 13452 10928
rect 13403 10897 13415 10900
rect 13357 10891 13415 10897
rect 13446 10888 13452 10900
rect 13504 10888 13510 10940
rect 15930 10888 15936 10940
rect 15988 10928 15994 10940
rect 16316 10931 16374 10937
rect 16316 10928 16328 10931
rect 15988 10900 16328 10928
rect 15988 10888 15994 10900
rect 16316 10897 16328 10900
rect 16362 10897 16374 10931
rect 16316 10891 16374 10897
rect 18325 10931 18383 10937
rect 18325 10897 18337 10931
rect 18371 10928 18383 10931
rect 18414 10928 18420 10940
rect 18371 10900 18420 10928
rect 18371 10897 18383 10900
rect 18325 10891 18383 10897
rect 18414 10888 18420 10900
rect 18472 10888 18478 10940
rect 18586 10931 18644 10937
rect 18586 10897 18598 10931
rect 18632 10928 18644 10931
rect 18800 10928 18828 10968
rect 18632 10900 18828 10928
rect 19352 10928 19380 10968
rect 21082 10956 21088 11008
rect 21140 10996 21146 11008
rect 21200 10999 21258 11005
rect 21200 10996 21212 10999
rect 21140 10968 21212 10996
rect 21140 10956 21146 10968
rect 21200 10965 21212 10968
rect 21246 10996 21258 10999
rect 21358 10996 21364 11008
rect 21246 10968 21364 10996
rect 21246 10965 21258 10968
rect 21200 10959 21258 10965
rect 21358 10956 21364 10968
rect 21416 10956 21422 11008
rect 22296 10968 23244 10996
rect 20162 10928 20168 10940
rect 19352 10900 20168 10928
rect 18632 10897 18644 10900
rect 18586 10891 18644 10897
rect 20162 10888 20168 10900
rect 20220 10888 20226 10940
rect 22097 10931 22155 10937
rect 22097 10897 22109 10931
rect 22143 10928 22155 10931
rect 22296 10928 22324 10968
rect 22143 10900 22324 10928
rect 23216 10928 23244 10968
rect 24029 10931 24087 10937
rect 24029 10928 24041 10931
rect 23216 10900 24041 10928
rect 22143 10897 22155 10900
rect 22097 10891 22155 10897
rect 24029 10897 24041 10900
rect 24075 10897 24087 10931
rect 24029 10891 24087 10897
rect 7282 10860 7288 10872
rect 7227 10832 7288 10860
rect 7282 10820 7288 10832
rect 7340 10820 7346 10872
rect 8941 10863 8999 10869
rect 8941 10829 8953 10863
rect 8987 10860 8999 10863
rect 9030 10860 9036 10872
rect 8987 10832 9036 10860
rect 8987 10829 8999 10832
rect 8941 10823 8999 10829
rect 9030 10820 9036 10832
rect 9088 10820 9094 10872
rect 13262 10860 13268 10872
rect 11730 10832 13268 10860
rect 13262 10820 13268 10832
rect 13320 10820 13326 10872
rect 16577 10863 16635 10869
rect 16577 10829 16589 10863
rect 16623 10860 16635 10863
rect 16850 10860 16856 10872
rect 16623 10832 16856 10860
rect 16623 10829 16635 10832
rect 16577 10823 16635 10829
rect 16850 10820 16856 10832
rect 16908 10820 16914 10872
rect 21450 10860 21456 10872
rect 21395 10832 21456 10860
rect 21450 10820 21456 10832
rect 21508 10820 21514 10872
rect 21910 10820 21916 10872
rect 21968 10860 21974 10872
rect 22005 10863 22063 10869
rect 22005 10860 22017 10863
rect 21968 10832 22017 10860
rect 21968 10820 21974 10832
rect 22005 10829 22017 10832
rect 22051 10829 22063 10863
rect 22005 10823 22063 10829
rect 22465 10863 22523 10869
rect 22465 10829 22477 10863
rect 22511 10860 22523 10863
rect 23109 10863 23167 10869
rect 23109 10860 23121 10863
rect 22511 10832 23121 10860
rect 22511 10829 22523 10832
rect 22465 10823 22523 10829
rect 23109 10829 23121 10832
rect 23155 10829 23167 10863
rect 23109 10823 23167 10829
rect 5736 10764 6408 10792
rect 5736 10520 5764 10764
rect 6380 10724 6408 10764
rect 10870 10752 10876 10804
rect 10928 10792 10934 10804
rect 11540 10795 11598 10801
rect 11540 10792 11552 10795
rect 10928 10764 11552 10792
rect 10928 10752 10934 10764
rect 11540 10761 11552 10764
rect 11586 10761 11598 10795
rect 15197 10795 15255 10801
rect 15197 10792 15209 10795
rect 11540 10755 11598 10761
rect 14476 10764 15209 10792
rect 14476 10736 14504 10764
rect 15197 10761 15209 10764
rect 15243 10761 15255 10795
rect 15197 10755 15255 10761
rect 6549 10727 6607 10733
rect 6549 10724 6561 10727
rect 6380 10696 6561 10724
rect 6549 10693 6561 10696
rect 6595 10693 6607 10727
rect 8662 10724 8668 10736
rect 8607 10696 8668 10724
rect 6549 10687 6607 10693
rect 8662 10684 8668 10696
rect 8720 10684 8726 10736
rect 9030 10684 9036 10736
rect 9088 10724 9094 10736
rect 9309 10727 9367 10733
rect 9309 10724 9321 10727
rect 9088 10696 9321 10724
rect 9088 10684 9094 10696
rect 9309 10693 9321 10696
rect 9355 10693 9367 10727
rect 9309 10687 9367 10693
rect 14458 10684 14464 10736
rect 14516 10684 14522 10736
rect 20073 10727 20131 10733
rect 20073 10693 20085 10727
rect 20119 10724 20131 10727
rect 20530 10724 20536 10736
rect 20119 10696 20536 10724
rect 20119 10693 20131 10696
rect 20073 10687 20131 10693
rect 20530 10684 20536 10696
rect 20588 10724 20594 10736
rect 21560 10730 23060 10758
rect 21560 10724 21588 10730
rect 20588 10696 21588 10724
rect 23032 10724 23060 10730
rect 26234 10724 26240 10736
rect 23032 10696 26240 10724
rect 20588 10684 20594 10696
rect 26234 10684 26240 10696
rect 26292 10684 26298 10736
rect 5796 10560 23000 10656
rect 6641 10523 6699 10529
rect 6641 10520 6653 10523
rect 5736 10492 6653 10520
rect 6641 10489 6653 10492
rect 6687 10489 6699 10523
rect 6641 10483 6699 10489
rect 10502 10480 10508 10532
rect 10560 10520 10566 10532
rect 10597 10523 10655 10529
rect 10597 10520 10609 10523
rect 10560 10492 10609 10520
rect 10560 10480 10566 10492
rect 10597 10489 10609 10492
rect 10643 10489 10655 10523
rect 10597 10483 10655 10489
rect 13262 10480 13268 10532
rect 13320 10520 13326 10532
rect 13449 10523 13507 10529
rect 13449 10520 13461 10523
rect 13320 10492 13461 10520
rect 13320 10480 13326 10492
rect 13449 10489 13461 10492
rect 13495 10489 13507 10523
rect 13449 10483 13507 10489
rect 14001 10523 14059 10529
rect 14001 10489 14013 10523
rect 14047 10520 14059 10523
rect 14550 10520 14556 10532
rect 14047 10492 14556 10520
rect 14047 10489 14059 10492
rect 14001 10483 14059 10489
rect 14550 10480 14556 10492
rect 14608 10480 14614 10532
rect 16114 10480 16120 10532
rect 16172 10520 16178 10532
rect 16209 10523 16267 10529
rect 16209 10520 16221 10523
rect 16172 10492 16221 10520
rect 16172 10480 16178 10492
rect 16209 10489 16221 10492
rect 16255 10489 16267 10523
rect 16209 10483 16267 10489
rect 18230 10480 18236 10532
rect 18288 10520 18294 10532
rect 18325 10523 18383 10529
rect 18325 10520 18337 10523
rect 18288 10492 18337 10520
rect 18288 10480 18294 10492
rect 18325 10489 18337 10492
rect 18371 10520 18383 10523
rect 18371 10492 20208 10520
rect 18371 10489 18383 10492
rect 18325 10483 18383 10489
rect 6549 10455 6607 10461
rect 6549 10421 6561 10455
rect 6595 10452 6607 10455
rect 7009 10455 7067 10461
rect 7009 10452 7021 10455
rect 6595 10424 7021 10452
rect 6595 10421 6607 10424
rect 6549 10415 6607 10421
rect 7009 10421 7021 10424
rect 7055 10452 7067 10455
rect 8662 10452 8668 10464
rect 7055 10424 7328 10452
rect 7055 10421 7067 10424
rect 7009 10415 7067 10421
rect 7300 10384 7328 10424
rect 8496 10424 8668 10452
rect 8496 10384 8524 10424
rect 8662 10412 8668 10424
rect 8720 10412 8726 10464
rect 11330 10452 11336 10464
rect 11275 10424 11336 10452
rect 11330 10412 11336 10424
rect 11388 10412 11394 10464
rect 17678 10452 17684 10464
rect 17623 10424 17684 10452
rect 17678 10412 17684 10424
rect 17736 10412 17742 10464
rect 20180 10452 20208 10492
rect 20254 10480 20260 10532
rect 20312 10520 20318 10532
rect 20312 10492 20373 10520
rect 20312 10480 20318 10492
rect 20180 10424 20944 10452
rect 18788 10396 18840 10402
rect 6380 10356 6960 10384
rect 7300 10356 8524 10384
rect 11517 10387 11575 10393
rect 6273 10319 6331 10325
rect 6273 10316 6285 10319
rect 5736 10288 6285 10316
rect 5736 9976 5764 10288
rect 6273 10285 6285 10288
rect 6319 10316 6331 10319
rect 6380 10316 6408 10356
rect 6319 10288 6408 10316
rect 6319 10285 6331 10288
rect 6273 10279 6331 10285
rect 6822 10276 6828 10328
rect 6880 10276 6886 10328
rect 6932 10316 6960 10356
rect 11517 10353 11529 10387
rect 11563 10384 11575 10387
rect 11606 10384 11612 10396
rect 11563 10356 11612 10384
rect 11563 10353 11575 10356
rect 11517 10347 11575 10353
rect 11606 10344 11612 10356
rect 11664 10344 11670 10396
rect 17954 10344 17960 10396
rect 18012 10344 18018 10396
rect 18785 10384 18788 10393
rect 20916 10393 20944 10424
rect 18724 10356 18788 10384
rect 18785 10347 18788 10356
rect 18840 10347 18843 10393
rect 20901 10387 20959 10393
rect 20901 10353 20913 10387
rect 20947 10384 20959 10387
rect 21266 10384 21272 10396
rect 20947 10356 21272 10384
rect 20947 10353 20959 10356
rect 20901 10347 20959 10353
rect 21266 10344 21272 10356
rect 21324 10344 21330 10396
rect 7101 10319 7159 10325
rect 7101 10316 7113 10319
rect 6932 10288 7113 10316
rect 7101 10285 7113 10288
rect 7147 10285 7159 10319
rect 7101 10279 7159 10285
rect 9122 10276 9128 10328
rect 9180 10316 9186 10328
rect 9217 10319 9275 10325
rect 9217 10316 9229 10319
rect 9180 10288 9229 10316
rect 9180 10276 9186 10288
rect 9217 10285 9229 10288
rect 9263 10285 9275 10319
rect 9217 10279 9275 10285
rect 12069 10319 12127 10325
rect 12069 10285 12081 10319
rect 12115 10316 12127 10319
rect 12342 10316 12348 10328
rect 12115 10288 12348 10316
rect 12115 10285 12127 10288
rect 12069 10279 12127 10285
rect 12342 10276 12348 10288
rect 12400 10276 12406 10328
rect 13262 10276 13268 10328
rect 13320 10316 13326 10328
rect 14182 10316 14188 10328
rect 13320 10288 14188 10316
rect 13320 10276 13326 10288
rect 14182 10276 14188 10288
rect 14240 10276 14246 10328
rect 14369 10319 14427 10325
rect 14369 10285 14381 10319
rect 14415 10316 14427 10319
rect 14458 10316 14464 10328
rect 14415 10288 14464 10316
rect 14415 10285 14427 10288
rect 14369 10279 14427 10285
rect 14458 10276 14464 10288
rect 14516 10276 14522 10328
rect 14553 10319 14611 10325
rect 14553 10285 14565 10319
rect 14599 10316 14611 10319
rect 15286 10316 15292 10328
rect 14599 10288 15292 10316
rect 14599 10285 14611 10288
rect 14553 10279 14611 10285
rect 15286 10276 15292 10288
rect 15344 10276 15350 10328
rect 16025 10319 16083 10325
rect 16025 10285 16037 10319
rect 16071 10316 16083 10319
rect 16850 10316 16856 10328
rect 16071 10288 16856 10316
rect 16071 10285 16083 10288
rect 16025 10279 16083 10285
rect 16850 10276 16856 10288
rect 16908 10316 16914 10328
rect 17589 10319 17647 10325
rect 17589 10316 17601 10319
rect 16908 10288 17601 10316
rect 16908 10276 16914 10288
rect 17589 10285 17601 10288
rect 17635 10285 17647 10319
rect 17589 10279 17647 10285
rect 17865 10319 17923 10325
rect 17865 10285 17877 10319
rect 17911 10316 17923 10319
rect 17972 10316 18000 10344
rect 18788 10338 18840 10344
rect 17911 10288 18000 10316
rect 17911 10285 17923 10288
rect 17865 10279 17923 10285
rect 18046 10276 18052 10328
rect 18104 10316 18110 10328
rect 18104 10288 18165 10316
rect 18104 10276 18110 10288
rect 20346 10276 20352 10328
rect 20404 10316 20410 10328
rect 20441 10319 20499 10325
rect 20441 10316 20453 10319
rect 20404 10288 20453 10316
rect 20404 10276 20410 10288
rect 20441 10285 20453 10288
rect 20487 10285 20499 10319
rect 20622 10316 20628 10328
rect 20567 10288 20628 10316
rect 20441 10279 20499 10285
rect 20622 10276 20628 10288
rect 20680 10276 20686 10328
rect 21361 10319 21419 10325
rect 21361 10285 21373 10319
rect 21407 10316 21419 10319
rect 21450 10316 21456 10328
rect 21407 10288 21456 10316
rect 21407 10285 21419 10288
rect 21361 10279 21419 10285
rect 21450 10276 21456 10288
rect 21508 10276 21514 10328
rect 23198 10316 23204 10328
rect 21560 10288 23204 10316
rect 6365 10251 6423 10257
rect 6365 10217 6377 10251
rect 6411 10248 6423 10251
rect 6840 10248 6868 10276
rect 6411 10220 6868 10248
rect 6411 10217 6423 10220
rect 6365 10211 6423 10217
rect 9030 10208 9036 10260
rect 9088 10248 9094 10260
rect 9478 10251 9536 10257
rect 9478 10248 9490 10251
rect 9088 10220 9490 10248
rect 9088 10208 9094 10220
rect 9478 10217 9490 10220
rect 9524 10217 9536 10251
rect 9478 10211 9536 10217
rect 11793 10251 11851 10257
rect 11793 10217 11805 10251
rect 11839 10248 11851 10251
rect 14277 10251 14335 10257
rect 11839 10242 12383 10248
rect 11839 10220 12337 10242
rect 11839 10217 11851 10220
rect 11793 10211 11851 10217
rect 12325 10208 12337 10220
rect 12371 10208 12383 10242
rect 14277 10217 14289 10251
rect 14323 10217 14335 10251
rect 14277 10211 14335 10217
rect 15764 10251 15822 10257
rect 15764 10217 15776 10251
rect 15810 10248 15822 10251
rect 16114 10248 16120 10260
rect 15810 10220 16120 10248
rect 15810 10217 15822 10220
rect 15764 10211 15822 10217
rect 12325 10202 12383 10208
rect 14292 10180 14320 10211
rect 16114 10208 16120 10220
rect 16172 10208 16178 10260
rect 17310 10248 17316 10260
rect 17368 10257 17374 10260
rect 17368 10251 17386 10257
rect 17267 10220 17316 10248
rect 17310 10208 17316 10220
rect 17374 10217 17386 10251
rect 17957 10251 18015 10257
rect 17957 10248 17969 10251
rect 17368 10211 17386 10217
rect 17512 10220 17969 10248
rect 17368 10208 17374 10211
rect 14550 10180 14556 10192
rect 14292 10152 14556 10180
rect 14550 10140 14556 10152
rect 14608 10140 14614 10192
rect 14645 10183 14703 10189
rect 14645 10149 14657 10183
rect 14691 10180 14703 10183
rect 14918 10180 14924 10192
rect 14691 10152 14924 10180
rect 14691 10149 14703 10152
rect 14645 10143 14703 10149
rect 14918 10140 14924 10152
rect 14976 10140 14982 10192
rect 17218 10140 17224 10192
rect 17276 10180 17282 10192
rect 17512 10180 17540 10220
rect 17957 10217 17969 10220
rect 18003 10217 18015 10251
rect 19046 10251 19104 10257
rect 19046 10248 19058 10251
rect 17957 10211 18015 10217
rect 18524 10220 19058 10248
rect 17276 10152 17540 10180
rect 17276 10140 17282 10152
rect 18138 10140 18144 10192
rect 18196 10180 18202 10192
rect 18524 10180 18552 10220
rect 19046 10217 19058 10220
rect 19092 10217 19104 10251
rect 19046 10211 19104 10217
rect 20533 10251 20591 10257
rect 20533 10217 20545 10251
rect 20579 10248 20591 10251
rect 21560 10248 21588 10288
rect 23198 10276 23204 10288
rect 23256 10276 23262 10328
rect 20579 10220 21588 10248
rect 21622 10251 21680 10257
rect 20579 10217 20591 10220
rect 20533 10211 20591 10217
rect 21622 10217 21634 10251
rect 21668 10248 21680 10251
rect 21910 10248 21916 10260
rect 21668 10220 21916 10248
rect 21668 10217 21680 10220
rect 21622 10211 21680 10217
rect 21910 10208 21916 10220
rect 21968 10208 21974 10260
rect 18196 10152 18552 10180
rect 20165 10183 20223 10189
rect 18196 10140 18202 10152
rect 20165 10149 20177 10183
rect 20211 10180 20223 10183
rect 20806 10180 20812 10192
rect 20211 10152 20812 10180
rect 20211 10149 20223 10152
rect 20165 10143 20223 10149
rect 20806 10140 20812 10152
rect 20864 10140 20870 10192
rect 22738 10180 22744 10192
rect 22683 10152 22744 10180
rect 22738 10140 22744 10152
rect 22796 10140 22802 10192
rect 5796 10016 23000 10112
rect 5997 9979 6055 9985
rect 5997 9976 6009 9979
rect 5736 9948 6009 9976
rect 5997 9945 6009 9948
rect 6043 9945 6055 9979
rect 5997 9939 6055 9945
rect 6181 9979 6239 9985
rect 6181 9945 6193 9979
rect 6227 9976 6239 9979
rect 6454 9976 6460 9988
rect 6227 9948 6460 9976
rect 6227 9945 6239 9948
rect 6181 9939 6239 9945
rect 6454 9936 6460 9948
rect 6512 9976 6518 9988
rect 6733 9979 6791 9985
rect 6733 9976 6745 9979
rect 6512 9948 6745 9976
rect 6512 9936 6518 9948
rect 6733 9945 6745 9948
rect 6779 9945 6791 9979
rect 6733 9939 6791 9945
rect 8846 9936 8852 9988
rect 8904 9976 8910 9988
rect 17313 9979 17371 9985
rect 8904 9948 9076 9976
rect 8904 9936 8910 9948
rect 6825 9911 6883 9917
rect 6825 9908 6837 9911
rect 6012 9880 6224 9908
rect 5905 9843 5963 9849
rect 5905 9809 5917 9843
rect 5951 9840 5963 9843
rect 6012 9840 6040 9880
rect 5951 9812 6040 9840
rect 6196 9840 6224 9880
rect 6564 9880 6837 9908
rect 6564 9849 6592 9880
rect 6825 9877 6837 9880
rect 6871 9877 6883 9911
rect 9048 9908 9076 9948
rect 17313 9945 17325 9979
rect 17359 9976 17371 9979
rect 17494 9976 17500 9988
rect 17359 9948 17500 9976
rect 17359 9945 17371 9948
rect 17313 9939 17371 9945
rect 17494 9936 17500 9948
rect 17552 9936 17558 9988
rect 18046 9976 18052 9988
rect 17991 9948 18052 9976
rect 18046 9936 18052 9948
rect 18104 9936 18110 9988
rect 18230 9976 18236 9988
rect 18156 9948 18236 9976
rect 9309 9911 9367 9917
rect 9309 9908 9321 9911
rect 9048 9880 9321 9908
rect 6825 9871 6883 9877
rect 9309 9877 9321 9880
rect 9355 9877 9367 9911
rect 9309 9871 9367 9877
rect 14918 9868 14924 9920
rect 14976 9908 14982 9920
rect 15473 9911 15531 9917
rect 15473 9908 15485 9911
rect 14976 9880 15485 9908
rect 14976 9868 14982 9880
rect 15473 9877 15485 9880
rect 15519 9877 15531 9911
rect 15473 9871 15531 9877
rect 16194 9911 16252 9917
rect 16194 9877 16206 9911
rect 16240 9908 16252 9911
rect 16390 9908 16396 9920
rect 16240 9880 16396 9908
rect 16240 9877 16252 9880
rect 16194 9871 16252 9877
rect 16390 9868 16396 9880
rect 16448 9868 16454 9920
rect 6549 9843 6607 9849
rect 6549 9840 6561 9843
rect 6196 9812 6561 9840
rect 5951 9809 5963 9812
rect 5905 9803 5963 9809
rect 6549 9809 6561 9812
rect 6595 9809 6607 9843
rect 6549 9803 6607 9809
rect 7009 9843 7067 9849
rect 7009 9809 7021 9843
rect 7055 9840 7067 9843
rect 10686 9840 10692 9852
rect 7055 9812 8064 9840
rect 9062 9812 10692 9840
rect 7055 9809 7067 9812
rect 7009 9803 7067 9809
rect 7837 9775 7895 9781
rect 7837 9741 7849 9775
rect 7883 9772 7895 9775
rect 7883 9744 7972 9772
rect 8036 9758 8064 9812
rect 10686 9800 10692 9812
rect 10744 9840 10750 9852
rect 12618 9849 12624 9852
rect 12606 9843 12624 9849
rect 12606 9840 12618 9843
rect 10744 9812 10902 9840
rect 12563 9812 12618 9840
rect 10744 9800 10750 9812
rect 12606 9809 12618 9812
rect 12606 9803 12624 9809
rect 12618 9800 12624 9803
rect 12676 9800 12682 9852
rect 15286 9840 15292 9852
rect 15231 9812 15292 9840
rect 15286 9800 15292 9812
rect 15344 9800 15350 9852
rect 15562 9840 15568 9852
rect 15507 9812 15568 9840
rect 15562 9800 15568 9812
rect 15620 9800 15626 9852
rect 15657 9843 15715 9849
rect 15657 9809 15669 9843
rect 15703 9809 15715 9843
rect 15657 9803 15715 9809
rect 15933 9843 15991 9849
rect 15933 9809 15945 9843
rect 15979 9840 15991 9843
rect 16022 9840 16028 9852
rect 15979 9812 16028 9840
rect 15979 9809 15991 9812
rect 15933 9803 15991 9809
rect 7883 9741 7895 9744
rect 7837 9735 7895 9741
rect 6365 9639 6423 9645
rect 6365 9636 6377 9639
rect 5736 9608 6377 9636
rect 5736 9296 5764 9608
rect 6365 9605 6377 9608
rect 6411 9605 6423 9639
rect 7944 9636 7972 9744
rect 8294 9732 8300 9784
rect 8352 9732 8358 9784
rect 10042 9732 10048 9784
rect 10100 9772 10106 9784
rect 10137 9775 10195 9781
rect 10137 9772 10149 9775
rect 10100 9744 10149 9772
rect 10100 9732 10106 9744
rect 10137 9741 10149 9744
rect 10183 9741 10195 9775
rect 10137 9735 10195 9741
rect 11330 9732 11336 9784
rect 11388 9732 11394 9784
rect 12342 9772 12348 9784
rect 12287 9744 12348 9772
rect 12342 9732 12348 9744
rect 12400 9732 12406 9784
rect 14274 9732 14280 9784
rect 14332 9772 14338 9784
rect 15672 9772 15700 9803
rect 16022 9800 16028 9812
rect 16080 9800 16086 9852
rect 16758 9800 16764 9852
rect 16816 9840 16822 9852
rect 18156 9840 18184 9948
rect 18230 9936 18236 9948
rect 18288 9936 18294 9988
rect 20622 9936 20628 9988
rect 20680 9976 20686 9988
rect 21453 9979 21511 9985
rect 21453 9976 21465 9979
rect 20680 9948 21465 9976
rect 20680 9936 20686 9948
rect 21453 9945 21465 9948
rect 21499 9945 21511 9979
rect 22462 9976 22468 9988
rect 22407 9948 22468 9976
rect 21453 9939 21511 9945
rect 22462 9936 22468 9948
rect 22520 9936 22526 9988
rect 22005 9911 22063 9917
rect 22005 9877 22017 9911
rect 22051 9908 22063 9911
rect 23753 9911 23811 9917
rect 23753 9908 23765 9911
rect 22051 9880 22508 9908
rect 22051 9877 22063 9880
rect 22005 9871 22063 9877
rect 16816 9812 18184 9840
rect 18328 9852 18380 9858
rect 16816 9800 16822 9812
rect 19334 9800 19340 9852
rect 19392 9840 19398 9852
rect 20073 9843 20131 9849
rect 20073 9840 20085 9843
rect 19392 9812 20085 9840
rect 19392 9800 19398 9812
rect 20073 9809 20085 9812
rect 20119 9809 20131 9843
rect 20073 9803 20131 9809
rect 20162 9800 20168 9852
rect 20220 9840 20226 9852
rect 20334 9843 20392 9849
rect 20334 9840 20346 9843
rect 20220 9812 20346 9840
rect 20220 9800 20226 9812
rect 20334 9809 20346 9812
rect 20380 9809 20392 9843
rect 20334 9803 20392 9809
rect 20806 9800 20812 9852
rect 20864 9840 20870 9852
rect 21821 9843 21879 9849
rect 21821 9840 21833 9843
rect 20864 9812 21833 9840
rect 20864 9800 20870 9812
rect 21821 9809 21833 9812
rect 21867 9840 21879 9843
rect 22186 9840 22192 9852
rect 21867 9812 22192 9840
rect 21867 9809 21879 9812
rect 21821 9803 21879 9809
rect 22186 9800 22192 9812
rect 22244 9840 22250 9852
rect 22281 9843 22339 9849
rect 22281 9840 22293 9843
rect 22244 9812 22293 9840
rect 22244 9800 22250 9812
rect 22281 9809 22293 9812
rect 22327 9809 22339 9843
rect 22480 9840 22508 9880
rect 23032 9880 23765 9908
rect 23032 9840 23060 9880
rect 23753 9877 23765 9880
rect 23799 9877 23811 9911
rect 23753 9871 23811 9877
rect 22480 9812 23060 9840
rect 22281 9803 22339 9809
rect 18328 9794 18380 9800
rect 15746 9772 15752 9784
rect 14332 9744 15752 9772
rect 14332 9732 14338 9744
rect 15746 9732 15752 9744
rect 15804 9732 15810 9784
rect 8202 9713 8208 9716
rect 8182 9707 8208 9713
rect 8182 9704 8194 9707
rect 8147 9676 8194 9704
rect 8182 9673 8194 9676
rect 8182 9667 8208 9673
rect 8202 9664 8208 9667
rect 8260 9664 8266 9716
rect 9953 9707 10011 9713
rect 9953 9704 9965 9707
rect 9600 9676 9965 9704
rect 9600 9670 9628 9676
rect 8404 9642 9628 9670
rect 9953 9673 9965 9676
rect 9999 9673 10011 9707
rect 9953 9667 10011 9673
rect 10689 9707 10747 9713
rect 10689 9673 10701 9707
rect 10735 9704 10747 9707
rect 10870 9704 10876 9716
rect 10735 9676 10876 9704
rect 10735 9673 10747 9676
rect 10689 9667 10747 9673
rect 10870 9664 10876 9676
rect 10928 9664 10934 9716
rect 11054 9664 11060 9716
rect 11112 9704 11118 9716
rect 11724 9707 11782 9713
rect 11724 9704 11736 9707
rect 11112 9676 11736 9704
rect 11112 9664 11118 9676
rect 11724 9673 11736 9676
rect 11770 9673 11782 9707
rect 11724 9667 11782 9673
rect 15841 9707 15899 9713
rect 15841 9673 15853 9707
rect 15887 9704 15899 9707
rect 15930 9704 15936 9716
rect 15887 9676 15936 9704
rect 15887 9673 15899 9676
rect 15841 9667 15899 9673
rect 15930 9664 15936 9676
rect 15988 9664 15994 9716
rect 19150 9704 19156 9716
rect 17604 9676 18184 9704
rect 19095 9676 19156 9704
rect 8404 9636 8432 9642
rect 10318 9636 10324 9648
rect 7944 9608 8432 9636
rect 10263 9608 10324 9636
rect 6365 9599 6423 9605
rect 10318 9596 10324 9608
rect 10376 9596 10382 9648
rect 12046 9639 12104 9645
rect 12046 9605 12058 9639
rect 12092 9636 12104 9639
rect 12986 9636 12992 9648
rect 12092 9608 12992 9636
rect 12092 9605 12104 9608
rect 12046 9599 12104 9605
rect 12986 9596 12992 9608
rect 13044 9596 13050 9648
rect 13725 9639 13783 9645
rect 13725 9605 13737 9639
rect 13771 9636 13783 9639
rect 14274 9636 14280 9648
rect 13771 9608 14280 9636
rect 13771 9605 13783 9608
rect 13725 9599 13783 9605
rect 14274 9596 14280 9608
rect 14332 9596 14338 9648
rect 17034 9596 17040 9648
rect 17092 9636 17098 9648
rect 17402 9636 17408 9648
rect 17092 9608 17408 9636
rect 17092 9596 17098 9608
rect 17402 9596 17408 9608
rect 17460 9636 17466 9648
rect 17604 9636 17632 9676
rect 18156 9670 18184 9676
rect 18156 9642 18920 9670
rect 19150 9664 19156 9676
rect 19208 9664 19214 9716
rect 21634 9704 21640 9716
rect 21579 9676 21640 9704
rect 21634 9664 21640 9676
rect 21692 9664 21698 9716
rect 22097 9707 22155 9713
rect 22097 9673 22109 9707
rect 22143 9704 22155 9707
rect 22186 9704 22192 9716
rect 22143 9676 22192 9704
rect 22143 9673 22155 9676
rect 22097 9667 22155 9673
rect 22186 9664 22192 9676
rect 22244 9664 22250 9716
rect 17460 9608 17632 9636
rect 18892 9636 18920 9642
rect 19429 9639 19487 9645
rect 19429 9636 19441 9639
rect 18892 9608 19441 9636
rect 17460 9596 17466 9608
rect 19429 9605 19441 9608
rect 19475 9605 19487 9639
rect 19429 9599 19487 9605
rect 5796 9472 23000 9568
rect 8294 9432 8300 9444
rect 8239 9404 8300 9432
rect 8294 9392 8300 9404
rect 8352 9392 8358 9444
rect 10686 9432 10692 9444
rect 10631 9404 10692 9432
rect 10686 9392 10692 9404
rect 10744 9392 10750 9444
rect 11330 9392 11336 9444
rect 11388 9432 11394 9444
rect 11517 9435 11575 9441
rect 11517 9432 11529 9435
rect 11388 9404 11529 9432
rect 11388 9392 11394 9404
rect 11517 9401 11529 9404
rect 11563 9401 11575 9435
rect 11517 9395 11575 9401
rect 11606 9392 11612 9444
rect 11664 9432 11670 9444
rect 11664 9404 13124 9432
rect 11664 9392 11670 9404
rect 6457 9367 6515 9373
rect 6457 9364 6469 9367
rect 6288 9336 6469 9364
rect 6288 9296 6316 9336
rect 6457 9333 6469 9336
rect 6503 9333 6515 9367
rect 6457 9327 6515 9333
rect 10318 9324 10324 9376
rect 10376 9324 10382 9376
rect 12986 9364 12992 9376
rect 12931 9336 12992 9364
rect 12986 9324 12992 9336
rect 13044 9324 13050 9376
rect 6638 9296 6644 9308
rect 5736 9268 6316 9296
rect 6583 9268 6644 9296
rect 6638 9256 6644 9268
rect 6696 9256 6702 9308
rect 9122 9256 9128 9308
rect 9180 9296 9186 9308
rect 9309 9299 9367 9305
rect 9309 9296 9321 9299
rect 9180 9268 9321 9296
rect 9180 9256 9186 9268
rect 9309 9265 9321 9268
rect 9355 9265 9367 9299
rect 9309 9259 9367 9265
rect 6917 9231 6975 9237
rect 6917 9197 6929 9231
rect 6963 9228 6975 9231
rect 7190 9228 7196 9240
rect 6963 9200 7196 9228
rect 6963 9197 6975 9200
rect 6917 9191 6975 9197
rect 7190 9188 7196 9200
rect 7248 9188 7254 9240
rect 9570 9231 9628 9237
rect 9570 9197 9582 9231
rect 9616 9228 9628 9231
rect 10336 9228 10364 9324
rect 13096 9308 13124 9404
rect 14550 9392 14556 9444
rect 14608 9432 14614 9444
rect 15013 9435 15071 9441
rect 15013 9432 15025 9435
rect 14608 9404 15025 9432
rect 14608 9392 14614 9404
rect 15013 9401 15025 9404
rect 15059 9401 15071 9435
rect 15013 9395 15071 9401
rect 16114 9392 16120 9444
rect 16172 9432 16178 9444
rect 16209 9435 16267 9441
rect 16209 9432 16221 9435
rect 16172 9404 16221 9432
rect 16172 9392 16178 9404
rect 16209 9401 16221 9404
rect 16255 9401 16267 9435
rect 16209 9395 16267 9401
rect 20162 9392 20168 9444
rect 20220 9432 20226 9444
rect 20257 9435 20315 9441
rect 20257 9432 20269 9435
rect 20220 9404 20269 9432
rect 20220 9392 20226 9404
rect 20257 9401 20269 9404
rect 20303 9401 20315 9435
rect 20257 9395 20315 9401
rect 21545 9435 21603 9441
rect 21545 9401 21557 9435
rect 21591 9432 21603 9435
rect 21634 9432 21640 9444
rect 21591 9404 21640 9432
rect 21591 9401 21603 9404
rect 21545 9395 21603 9401
rect 21634 9392 21640 9404
rect 21692 9392 21698 9444
rect 23382 9432 23388 9444
rect 22020 9404 22416 9432
rect 19978 9324 19984 9376
rect 20036 9364 20042 9376
rect 20036 9336 20668 9364
rect 20036 9324 20042 9336
rect 13078 9256 13084 9308
rect 13136 9296 13142 9308
rect 13173 9299 13231 9305
rect 13173 9296 13185 9299
rect 13136 9268 13185 9296
rect 13136 9256 13142 9268
rect 13173 9265 13185 9268
rect 13219 9265 13231 9299
rect 13173 9259 13231 9265
rect 13446 9256 13452 9308
rect 13504 9296 13510 9308
rect 13633 9299 13691 9305
rect 13633 9296 13645 9299
rect 13504 9268 13645 9296
rect 13504 9256 13510 9268
rect 13633 9265 13645 9268
rect 13679 9265 13691 9299
rect 13633 9259 13691 9265
rect 12897 9231 12955 9237
rect 12897 9228 12909 9231
rect 9616 9200 10364 9228
rect 12544 9200 12909 9228
rect 9616 9197 9628 9200
rect 9570 9191 9628 9197
rect 6825 9163 6883 9169
rect 6825 9129 6837 9163
rect 6871 9160 6883 9163
rect 6871 9154 7236 9160
rect 6871 9132 7190 9154
rect 6871 9129 6883 9132
rect 6825 9123 6883 9129
rect 7178 9120 7190 9132
rect 7224 9120 7236 9154
rect 7178 9114 7236 9120
rect 11716 9132 12296 9160
rect 11517 9095 11575 9101
rect 11517 9061 11529 9095
rect 11563 9092 11575 9095
rect 11716 9092 11744 9132
rect 11563 9064 11744 9092
rect 12268 9092 12296 9132
rect 12434 9120 12440 9172
rect 12492 9160 12498 9172
rect 12544 9160 12572 9200
rect 12897 9197 12909 9200
rect 12943 9197 12955 9231
rect 12897 9191 12955 9197
rect 15838 9188 15844 9240
rect 15896 9228 15902 9240
rect 16393 9231 16451 9237
rect 16393 9228 16405 9231
rect 15896 9200 16405 9228
rect 15896 9188 15902 9200
rect 16393 9197 16405 9200
rect 16439 9197 16451 9231
rect 16758 9228 16764 9240
rect 16703 9200 16764 9228
rect 16393 9191 16451 9197
rect 16758 9188 16764 9200
rect 16816 9188 16822 9240
rect 17678 9188 17684 9240
rect 17736 9228 17742 9240
rect 17972 9231 18030 9237
rect 17972 9228 17984 9231
rect 17736 9200 17984 9228
rect 17736 9188 17742 9200
rect 17972 9197 17984 9200
rect 18018 9197 18030 9231
rect 17972 9191 18030 9197
rect 18690 9188 18696 9240
rect 18748 9228 18754 9240
rect 18785 9231 18843 9237
rect 18785 9228 18797 9231
rect 18748 9200 18797 9228
rect 18748 9188 18754 9200
rect 18785 9197 18797 9200
rect 18831 9197 18843 9231
rect 18785 9191 18843 9197
rect 20346 9188 20352 9240
rect 20404 9228 20410 9240
rect 20640 9237 20668 9336
rect 22020 9305 22048 9404
rect 22388 9364 22416 9404
rect 23032 9404 23388 9432
rect 23032 9364 23060 9404
rect 23382 9392 23388 9404
rect 23440 9392 23446 9444
rect 22388 9336 23060 9364
rect 22005 9299 22063 9305
rect 20824 9268 21312 9296
rect 20441 9231 20499 9237
rect 20441 9228 20453 9231
rect 20404 9200 20453 9228
rect 20404 9188 20410 9200
rect 20441 9197 20453 9200
rect 20487 9197 20499 9231
rect 20441 9191 20499 9197
rect 20625 9231 20683 9237
rect 20625 9197 20637 9231
rect 20671 9197 20683 9231
rect 20625 9191 20683 9197
rect 12492 9132 12572 9160
rect 12636 9163 12694 9169
rect 12492 9120 12498 9132
rect 12636 9129 12648 9163
rect 12682 9160 12694 9163
rect 13357 9163 13415 9169
rect 13357 9160 13369 9163
rect 12682 9132 13369 9160
rect 12682 9129 12694 9132
rect 12636 9123 12694 9129
rect 13357 9129 13369 9132
rect 13403 9129 13415 9163
rect 13894 9163 13952 9169
rect 13894 9160 13906 9163
rect 13357 9123 13415 9129
rect 13464 9132 13906 9160
rect 13464 9092 13492 9132
rect 13894 9129 13906 9132
rect 13940 9129 13952 9163
rect 16482 9160 16488 9172
rect 16427 9132 16488 9160
rect 13894 9123 13952 9129
rect 16482 9120 16488 9132
rect 16540 9120 16546 9172
rect 16577 9163 16635 9169
rect 16577 9129 16589 9163
rect 16623 9160 16635 9163
rect 16623 9132 16896 9160
rect 16623 9129 16635 9132
rect 16577 9123 16635 9129
rect 16868 9101 16896 9132
rect 18506 9120 18512 9172
rect 18564 9160 18570 9172
rect 19046 9163 19104 9169
rect 18564 9132 18644 9160
rect 18564 9120 18570 9132
rect 12268 9064 13492 9092
rect 16853 9095 16911 9101
rect 11563 9061 11575 9064
rect 11517 9055 11575 9061
rect 16853 9061 16865 9095
rect 16899 9061 16911 9095
rect 16853 9055 16911 9061
rect 18325 9095 18383 9101
rect 18325 9061 18337 9095
rect 18371 9092 18383 9095
rect 18616 9092 18644 9132
rect 19046 9129 19058 9163
rect 19092 9160 19104 9163
rect 19794 9160 19800 9172
rect 19092 9132 19800 9160
rect 19092 9129 19104 9132
rect 19046 9123 19104 9129
rect 19794 9120 19800 9132
rect 19852 9160 19858 9172
rect 19978 9160 19984 9172
rect 19852 9132 19984 9160
rect 19852 9120 19858 9132
rect 19978 9120 19984 9132
rect 20036 9120 20042 9172
rect 20533 9163 20591 9169
rect 20533 9160 20545 9163
rect 20180 9132 20545 9160
rect 19334 9092 19340 9104
rect 18371 9064 19340 9092
rect 18371 9061 18383 9064
rect 18325 9055 18383 9061
rect 19334 9052 19340 9064
rect 19392 9052 19398 9104
rect 20180 9101 20208 9132
rect 20533 9129 20545 9132
rect 20579 9160 20591 9163
rect 20824 9160 20852 9268
rect 21284 9228 21312 9268
rect 22005 9265 22017 9299
rect 22051 9265 22063 9299
rect 22005 9259 22063 9265
rect 22094 9256 22100 9308
rect 22152 9296 22158 9308
rect 22189 9299 22247 9305
rect 22189 9296 22201 9299
rect 22152 9268 22201 9296
rect 22152 9256 22158 9268
rect 22189 9265 22201 9268
rect 22235 9265 22247 9299
rect 22189 9259 22247 9265
rect 21284 9200 21864 9228
rect 20579 9132 20852 9160
rect 21836 9160 21864 9200
rect 22002 9160 22008 9172
rect 21836 9132 22008 9160
rect 20579 9129 20591 9132
rect 20533 9123 20591 9129
rect 22002 9120 22008 9132
rect 22060 9120 22066 9172
rect 20165 9095 20223 9101
rect 20165 9061 20177 9095
rect 20211 9061 20223 9095
rect 20165 9055 20223 9061
rect 20901 9095 20959 9101
rect 20901 9061 20913 9095
rect 20947 9092 20959 9095
rect 21174 9092 21180 9104
rect 20947 9064 21180 9092
rect 20947 9061 20959 9064
rect 20901 9055 20959 9061
rect 21174 9052 21180 9064
rect 21232 9052 21238 9104
rect 21818 9052 21824 9104
rect 21876 9092 21882 9104
rect 22373 9095 22431 9101
rect 22373 9092 22385 9095
rect 21876 9064 22385 9092
rect 21876 9052 21882 9064
rect 22373 9061 22385 9064
rect 22419 9061 22431 9095
rect 22373 9055 22431 9061
rect 5796 8928 23000 9024
rect 8113 8891 8171 8897
rect 8113 8857 8125 8891
rect 8159 8888 8171 8891
rect 8846 8888 8852 8900
rect 8159 8860 8852 8888
rect 8159 8857 8171 8860
rect 8113 8851 8171 8857
rect 8846 8848 8852 8860
rect 8904 8848 8910 8900
rect 11054 8888 11060 8900
rect 10796 8860 11060 8888
rect 7285 8823 7343 8829
rect 7285 8820 7297 8823
rect 6840 8792 7297 8820
rect 6454 8712 6460 8764
rect 6512 8752 6518 8764
rect 6549 8755 6607 8761
rect 6549 8752 6561 8755
rect 6512 8724 6561 8752
rect 6512 8712 6518 8724
rect 6549 8721 6561 8724
rect 6595 8752 6607 8755
rect 6840 8752 6868 8792
rect 7285 8789 7297 8792
rect 7331 8789 7343 8823
rect 7285 8783 7343 8789
rect 10505 8823 10563 8829
rect 10505 8789 10517 8823
rect 10551 8820 10563 8823
rect 10796 8820 10824 8860
rect 11054 8848 11060 8860
rect 11112 8848 11118 8900
rect 12618 8848 12624 8900
rect 12676 8888 12682 8900
rect 12989 8891 13047 8897
rect 12989 8888 13001 8891
rect 12676 8860 13001 8888
rect 12676 8848 12682 8860
rect 12989 8857 13001 8860
rect 13035 8857 13047 8891
rect 12989 8851 13047 8857
rect 13173 8891 13231 8897
rect 13173 8857 13185 8891
rect 13219 8888 13231 8891
rect 13262 8888 13268 8900
rect 13219 8860 13268 8888
rect 13219 8857 13231 8860
rect 13173 8851 13231 8857
rect 13262 8848 13268 8860
rect 13320 8848 13326 8900
rect 14737 8891 14795 8897
rect 14737 8857 14749 8891
rect 14783 8888 14795 8891
rect 15378 8888 15384 8900
rect 14783 8860 15384 8888
rect 14783 8857 14795 8860
rect 14737 8851 14795 8857
rect 15378 8848 15384 8860
rect 15436 8848 15442 8900
rect 16482 8848 16488 8900
rect 16540 8888 16546 8900
rect 16853 8891 16911 8897
rect 16853 8888 16865 8891
rect 16540 8860 16865 8888
rect 16540 8848 16546 8860
rect 16853 8857 16865 8860
rect 16899 8857 16911 8891
rect 16853 8851 16911 8857
rect 17497 8891 17555 8897
rect 17497 8857 17509 8891
rect 17543 8888 17555 8891
rect 17543 8860 19564 8888
rect 17543 8857 17555 8860
rect 17497 8851 17555 8857
rect 13618 8823 13676 8829
rect 13618 8820 13630 8823
rect 10551 8792 10824 8820
rect 11808 8792 12572 8820
rect 10551 8789 10563 8792
rect 10505 8783 10563 8789
rect 6595 8724 6868 8752
rect 6917 8755 6975 8761
rect 6595 8721 6607 8724
rect 6549 8715 6607 8721
rect 6917 8721 6929 8755
rect 6963 8752 6975 8755
rect 7377 8755 7435 8761
rect 7377 8752 7389 8755
rect 6963 8724 7389 8752
rect 6963 8721 6975 8724
rect 6917 8715 6975 8721
rect 7377 8721 7389 8724
rect 7423 8752 7435 8755
rect 7834 8752 7840 8764
rect 7423 8724 7840 8752
rect 7423 8721 7435 8724
rect 7377 8715 7435 8721
rect 7834 8712 7840 8724
rect 7892 8712 7898 8764
rect 10686 8752 10692 8764
rect 9338 8724 10692 8752
rect 10686 8712 10692 8724
rect 10744 8752 10750 8764
rect 10744 8724 10810 8752
rect 10744 8712 10750 8724
rect 11808 8670 11836 8792
rect 12544 8786 12572 8792
rect 13004 8792 13630 8820
rect 13004 8786 13032 8792
rect 12544 8758 13032 8786
rect 13618 8789 13630 8792
rect 13664 8820 13676 8823
rect 14274 8820 14280 8832
rect 13664 8792 14280 8820
rect 13664 8789 13676 8792
rect 13618 8783 13676 8789
rect 14274 8780 14280 8792
rect 14332 8780 14338 8832
rect 16942 8780 16948 8832
rect 17000 8820 17006 8832
rect 19536 8820 19564 8860
rect 20162 8848 20168 8900
rect 20220 8888 20226 8900
rect 21545 8891 21603 8897
rect 21545 8888 21557 8891
rect 20220 8860 21557 8888
rect 20220 8848 20226 8860
rect 21545 8857 21557 8860
rect 21591 8857 21603 8891
rect 21545 8851 21603 8857
rect 20073 8823 20131 8829
rect 20073 8820 20085 8823
rect 17000 8792 17448 8820
rect 17000 8780 17006 8792
rect 17420 8786 17448 8792
rect 18156 8792 19012 8820
rect 19536 8792 20085 8820
rect 18156 8786 18184 8792
rect 13262 8752 13268 8764
rect 13207 8724 13268 8752
rect 13262 8712 13268 8724
rect 13320 8712 13326 8764
rect 13357 8755 13415 8761
rect 13357 8721 13369 8755
rect 13403 8752 13415 8755
rect 13446 8752 13452 8764
rect 13403 8724 13452 8752
rect 13403 8721 13415 8724
rect 13357 8715 13415 8721
rect 13446 8712 13452 8724
rect 13504 8712 13510 8764
rect 15470 8752 15476 8764
rect 15415 8724 15476 8752
rect 15470 8712 15476 8724
rect 15528 8712 15534 8764
rect 15734 8755 15792 8761
rect 15734 8721 15746 8755
rect 15780 8752 15792 8755
rect 16206 8752 16212 8764
rect 15780 8724 16212 8752
rect 15780 8721 15792 8724
rect 15734 8715 15792 8721
rect 16206 8712 16212 8724
rect 16264 8712 16270 8764
rect 17420 8758 18184 8786
rect 18322 8712 18328 8764
rect 18380 8752 18386 8764
rect 18984 8752 19012 8792
rect 20073 8789 20085 8792
rect 20119 8789 20131 8823
rect 20073 8783 20131 8789
rect 19797 8755 19855 8761
rect 19797 8752 19809 8755
rect 18380 8724 18722 8752
rect 18984 8724 19809 8752
rect 18380 8712 18386 8724
rect 19797 8721 19809 8724
rect 19843 8721 19855 8755
rect 19797 8715 19855 8721
rect 19996 8724 20378 8752
rect 12805 8687 12863 8693
rect 7208 8588 8156 8616
rect 6365 8551 6423 8557
rect 6365 8548 6377 8551
rect 5736 8520 6377 8548
rect 5736 8344 5764 8520
rect 6365 8517 6377 8520
rect 6411 8517 6423 8551
rect 6365 8511 6423 8517
rect 6733 8551 6791 8557
rect 6733 8517 6745 8551
rect 6779 8548 6791 8551
rect 7009 8551 7067 8557
rect 7009 8548 7021 8551
rect 6779 8520 7021 8548
rect 6779 8517 6791 8520
rect 6733 8511 6791 8517
rect 7009 8517 7021 8520
rect 7055 8548 7067 8551
rect 7208 8548 7236 8588
rect 7055 8520 7236 8548
rect 8128 8548 8156 8588
rect 8312 8560 8340 8670
rect 12805 8653 12817 8687
rect 12851 8684 12863 8687
rect 13078 8684 13084 8696
rect 12851 8656 13084 8684
rect 12851 8653 12863 8656
rect 12805 8647 12863 8653
rect 13078 8644 13084 8656
rect 13136 8644 13142 8696
rect 14476 8656 15240 8684
rect 8466 8619 8524 8625
rect 8466 8585 8478 8619
rect 8512 8616 8524 8619
rect 10410 8616 10416 8628
rect 8512 8588 10416 8616
rect 8512 8585 8524 8588
rect 8466 8579 8524 8585
rect 10410 8576 10416 8588
rect 10468 8576 10474 8628
rect 11632 8619 11690 8625
rect 11632 8585 11644 8619
rect 11678 8616 11690 8619
rect 11678 8588 12756 8616
rect 11678 8585 11690 8588
rect 11632 8579 11690 8585
rect 12728 8582 12756 8588
rect 8294 8548 8300 8560
rect 8128 8520 8300 8548
rect 7055 8517 7067 8520
rect 7009 8511 7067 8517
rect 8294 8508 8300 8520
rect 8352 8508 8358 8560
rect 8662 8508 8668 8560
rect 8720 8548 8726 8560
rect 9493 8551 9551 8557
rect 12728 8554 13400 8582
rect 9493 8548 9505 8551
rect 8720 8520 9505 8548
rect 8720 8508 8726 8520
rect 9493 8517 9505 8520
rect 9539 8517 9551 8551
rect 13372 8548 13400 8554
rect 14476 8548 14504 8656
rect 13372 8520 14504 8548
rect 15212 8548 15240 8656
rect 16776 8656 18828 8684
rect 16666 8576 16672 8628
rect 16724 8616 16730 8628
rect 16776 8616 16804 8656
rect 18506 8616 18512 8628
rect 16724 8588 16804 8616
rect 18451 8588 18512 8616
rect 16724 8576 16730 8588
rect 18506 8576 18512 8588
rect 18564 8576 18570 8628
rect 18800 8616 18828 8656
rect 19613 8619 19671 8625
rect 19613 8616 19625 8619
rect 18800 8588 19625 8616
rect 19613 8585 19625 8588
rect 19659 8585 19671 8619
rect 19613 8579 19671 8585
rect 17497 8551 17555 8557
rect 17497 8548 17509 8551
rect 15212 8520 17509 8548
rect 9493 8511 9551 8517
rect 17497 8517 17509 8520
rect 17543 8517 17555 8551
rect 17497 8511 17555 8517
rect 17586 8508 17592 8560
rect 17644 8548 17650 8560
rect 19996 8548 20024 8724
rect 20254 8644 20260 8696
rect 20312 8684 20318 8696
rect 20312 8656 20470 8684
rect 20312 8644 20318 8656
rect 20162 8576 20168 8628
rect 20220 8616 20226 8628
rect 21200 8619 21258 8625
rect 21200 8616 21212 8619
rect 20220 8588 20392 8616
rect 20220 8576 20226 8588
rect 20364 8582 20392 8588
rect 21008 8588 21212 8616
rect 21008 8582 21036 8588
rect 20364 8554 21036 8582
rect 21200 8585 21212 8588
rect 21246 8585 21258 8619
rect 21200 8579 21258 8585
rect 17644 8520 20024 8548
rect 17644 8508 17650 8520
rect 5796 8384 23000 8480
rect 6273 8347 6331 8353
rect 6273 8344 6285 8347
rect 5736 8316 6285 8344
rect 6273 8313 6285 8316
rect 6319 8313 6331 8347
rect 8294 8344 8300 8356
rect 8239 8316 8300 8344
rect 6273 8307 6331 8313
rect 8294 8304 8300 8316
rect 8352 8304 8358 8356
rect 10686 8344 10692 8356
rect 10631 8316 10692 8344
rect 10686 8304 10692 8316
rect 10744 8304 10750 8356
rect 13173 8347 13231 8353
rect 13173 8313 13185 8347
rect 13219 8344 13231 8347
rect 13262 8344 13268 8356
rect 13219 8316 13268 8344
rect 13219 8313 13231 8316
rect 13173 8307 13231 8313
rect 13262 8304 13268 8316
rect 13320 8304 13326 8356
rect 17218 8344 17224 8356
rect 16316 8316 16896 8344
rect 17163 8316 17224 8344
rect 16316 8310 16344 8316
rect 12437 8279 12495 8285
rect 12437 8245 12449 8279
rect 12483 8276 12495 8279
rect 13832 8282 16344 8310
rect 13832 8276 13860 8282
rect 16758 8276 16764 8288
rect 12483 8248 13860 8276
rect 16500 8248 16764 8276
rect 12483 8245 12495 8248
rect 12437 8239 12495 8245
rect 10686 8168 10692 8220
rect 10744 8208 10750 8220
rect 11057 8211 11115 8217
rect 11057 8208 11069 8211
rect 10744 8180 11069 8208
rect 10744 8168 10750 8180
rect 11057 8177 11069 8180
rect 11103 8177 11115 8211
rect 11057 8171 11115 8177
rect 13725 8211 13783 8217
rect 13725 8177 13737 8211
rect 13771 8208 13783 8211
rect 16500 8208 16528 8248
rect 16758 8236 16764 8248
rect 16816 8236 16822 8288
rect 13771 8180 16528 8208
rect 16868 8208 16896 8316
rect 17218 8304 17224 8316
rect 17276 8304 17282 8356
rect 18230 8304 18236 8356
rect 18288 8344 18294 8356
rect 18288 8316 18644 8344
rect 18288 8304 18294 8316
rect 17586 8276 17592 8288
rect 17328 8248 17592 8276
rect 17328 8208 17356 8248
rect 17586 8236 17592 8248
rect 17644 8236 17650 8288
rect 18616 8217 18644 8316
rect 18966 8304 18972 8356
rect 19024 8344 19030 8356
rect 20257 8347 20315 8353
rect 20257 8344 20269 8347
rect 19024 8316 20269 8344
rect 19024 8304 19030 8316
rect 20257 8313 20269 8316
rect 20303 8313 20315 8347
rect 20257 8307 20315 8313
rect 20901 8347 20959 8353
rect 20901 8313 20913 8347
rect 20947 8344 20959 8347
rect 21174 8344 21180 8356
rect 20947 8316 21180 8344
rect 20947 8313 20959 8316
rect 20901 8307 20959 8313
rect 21174 8304 21180 8316
rect 21232 8304 21238 8356
rect 22741 8347 22799 8353
rect 22741 8313 22753 8347
rect 22787 8344 22799 8347
rect 23198 8344 23204 8356
rect 22787 8316 23204 8344
rect 22787 8313 22799 8316
rect 22741 8307 22799 8313
rect 23198 8304 23204 8316
rect 23256 8304 23262 8356
rect 16868 8180 17356 8208
rect 18601 8211 18659 8217
rect 13771 8177 13783 8180
rect 13725 8171 13783 8177
rect 6549 8143 6607 8149
rect 6549 8109 6561 8143
rect 6595 8140 6607 8143
rect 6638 8140 6644 8152
rect 6595 8112 6644 8140
rect 6595 8109 6607 8112
rect 6549 8103 6607 8109
rect 6638 8100 6644 8112
rect 6696 8100 6702 8152
rect 6917 8143 6975 8149
rect 6917 8109 6929 8143
rect 6963 8140 6975 8143
rect 7190 8140 7196 8152
rect 6963 8112 7196 8140
rect 6963 8109 6975 8112
rect 6917 8103 6975 8109
rect 7190 8100 7196 8112
rect 7248 8100 7254 8152
rect 9122 8100 9128 8152
rect 9180 8140 9186 8152
rect 9309 8143 9367 8149
rect 9309 8140 9321 8143
rect 9180 8112 9321 8140
rect 9180 8100 9186 8112
rect 9309 8109 9321 8112
rect 9355 8109 9367 8143
rect 9309 8103 9367 8109
rect 11790 8100 11796 8152
rect 11848 8140 11854 8152
rect 13081 8143 13139 8149
rect 13081 8140 13093 8143
rect 11848 8112 13093 8140
rect 11848 8100 11854 8112
rect 13081 8109 13093 8112
rect 13127 8109 13139 8143
rect 14274 8140 14280 8152
rect 14219 8112 14280 8140
rect 13081 8103 13139 8109
rect 14274 8100 14280 8112
rect 14332 8100 14338 8152
rect 15010 8100 15016 8152
rect 15068 8140 15074 8152
rect 15304 8149 15332 8180
rect 18601 8177 18613 8211
rect 18647 8177 18659 8211
rect 18601 8171 18659 8177
rect 15105 8143 15163 8149
rect 15105 8140 15117 8143
rect 15068 8112 15117 8140
rect 15068 8100 15074 8112
rect 15105 8109 15117 8112
rect 15151 8109 15163 8143
rect 15105 8103 15163 8109
rect 15289 8143 15347 8149
rect 15289 8109 15301 8143
rect 15335 8109 15347 8143
rect 15289 8103 15347 8109
rect 18046 8100 18052 8152
rect 18104 8140 18110 8152
rect 18340 8143 18398 8149
rect 18340 8140 18352 8143
rect 18104 8112 18352 8140
rect 18104 8100 18110 8112
rect 18340 8109 18352 8112
rect 18386 8109 18398 8143
rect 18340 8103 18398 8109
rect 18506 8100 18512 8152
rect 18564 8140 18570 8152
rect 19058 8149 19064 8152
rect 18785 8143 18843 8149
rect 18785 8140 18797 8143
rect 18564 8112 18797 8140
rect 18564 8100 18570 8112
rect 18785 8109 18797 8112
rect 18831 8109 18843 8143
rect 19046 8143 19064 8149
rect 19046 8140 19058 8143
rect 19003 8112 19058 8140
rect 18785 8103 18843 8109
rect 19046 8109 19058 8112
rect 19046 8103 19064 8109
rect 19058 8100 19064 8103
rect 19116 8100 19122 8152
rect 20346 8100 20352 8152
rect 20404 8140 20410 8152
rect 20441 8143 20499 8149
rect 20441 8140 20453 8143
rect 20404 8112 20453 8140
rect 20404 8100 20410 8112
rect 20441 8109 20453 8112
rect 20487 8109 20499 8143
rect 20441 8103 20499 8109
rect 20530 8100 20536 8152
rect 20588 8140 20594 8152
rect 21361 8143 21419 8149
rect 20588 8112 20649 8140
rect 20588 8100 20594 8112
rect 21361 8109 21373 8143
rect 21407 8140 21419 8143
rect 21450 8140 21456 8152
rect 21407 8112 21456 8140
rect 21407 8109 21419 8112
rect 21361 8103 21419 8109
rect 21450 8100 21456 8112
rect 21508 8100 21514 8152
rect 6733 8075 6791 8081
rect 6733 8041 6745 8075
rect 6779 8072 6791 8075
rect 6779 8066 7231 8072
rect 6779 8044 7185 8066
rect 6779 8041 6791 8044
rect 6733 8035 6791 8041
rect 7173 8032 7185 8044
rect 7219 8032 7231 8066
rect 9398 8032 9404 8084
rect 9456 8072 9462 8084
rect 11330 8081 11336 8084
rect 9570 8075 9628 8081
rect 9570 8072 9582 8075
rect 9456 8044 9582 8072
rect 9456 8032 9462 8044
rect 9570 8041 9582 8044
rect 9616 8041 9628 8075
rect 9570 8035 9628 8041
rect 11318 8075 11336 8081
rect 11318 8041 11330 8075
rect 11388 8072 11394 8084
rect 11388 8044 11437 8072
rect 11318 8035 11336 8041
rect 11330 8032 11336 8035
rect 11388 8032 11394 8044
rect 14826 8032 14832 8084
rect 14884 8072 14890 8084
rect 14921 8075 14979 8081
rect 14921 8072 14933 8075
rect 14884 8044 14933 8072
rect 14884 8032 14890 8044
rect 14921 8041 14933 8044
rect 14967 8041 14979 8075
rect 14921 8035 14979 8041
rect 15194 8032 15200 8084
rect 15252 8072 15258 8084
rect 19978 8072 19984 8084
rect 15252 8044 19984 8072
rect 15252 8032 15258 8044
rect 19978 8032 19984 8044
rect 20036 8032 20042 8084
rect 20625 8075 20683 8081
rect 20625 8041 20637 8075
rect 20671 8041 20683 8075
rect 20625 8035 20683 8041
rect 7173 8026 7231 8032
rect 11974 7964 11980 8016
rect 12032 8004 12038 8016
rect 12437 8007 12495 8013
rect 12437 8004 12449 8007
rect 12032 7976 12449 8004
rect 12032 7964 12038 7976
rect 12437 7973 12449 7976
rect 12483 7973 12495 8007
rect 13446 8004 13452 8016
rect 13391 7976 13452 8004
rect 12437 7967 12495 7973
rect 13446 7964 13452 7976
rect 13504 7964 13510 8016
rect 14458 7964 14464 8016
rect 14516 8004 14522 8016
rect 15105 8007 15163 8013
rect 15105 8004 15117 8007
rect 14516 7976 15117 8004
rect 14516 7964 14522 7976
rect 15105 7973 15117 7976
rect 15151 7973 15163 8007
rect 15105 7967 15163 7973
rect 20165 8007 20223 8013
rect 20165 7973 20177 8007
rect 20211 8004 20223 8007
rect 20640 8004 20668 8035
rect 20714 8032 20720 8084
rect 20772 8072 20778 8084
rect 21634 8081 21640 8084
rect 21622 8075 21640 8081
rect 21622 8072 21634 8075
rect 20772 8044 21634 8072
rect 20772 8032 20778 8044
rect 21622 8041 21634 8044
rect 21622 8035 21640 8041
rect 21634 8032 21640 8035
rect 21692 8032 21698 8084
rect 20211 7976 20668 8004
rect 20211 7973 20223 7976
rect 20165 7967 20223 7973
rect 5796 7840 23000 7936
rect 6917 7803 6975 7809
rect 6917 7769 6929 7803
rect 6963 7800 6975 7803
rect 9217 7803 9275 7809
rect 6963 7772 7497 7800
rect 6963 7769 6975 7772
rect 6917 7763 6975 7769
rect 7469 7741 7497 7772
rect 9217 7769 9229 7803
rect 9263 7800 9275 7803
rect 9398 7800 9404 7812
rect 9263 7772 9404 7800
rect 9263 7769 9275 7772
rect 9217 7763 9275 7769
rect 9398 7760 9404 7772
rect 9456 7760 9462 7812
rect 10042 7760 10048 7812
rect 10100 7800 10106 7812
rect 11241 7803 11299 7809
rect 10100 7772 11008 7800
rect 10100 7760 10106 7772
rect 7454 7735 7512 7741
rect 7116 7704 7420 7732
rect 6638 7664 6644 7676
rect 6583 7636 6644 7664
rect 6638 7624 6644 7636
rect 6696 7664 6702 7676
rect 7116 7664 7144 7704
rect 6696 7636 7144 7664
rect 7193 7667 7251 7673
rect 6696 7624 6702 7636
rect 7193 7633 7205 7667
rect 7239 7664 7251 7667
rect 7282 7664 7288 7676
rect 7239 7636 7288 7664
rect 7239 7633 7251 7636
rect 7193 7627 7251 7633
rect 7282 7624 7288 7636
rect 7340 7624 7346 7676
rect 7392 7664 7420 7704
rect 7454 7701 7466 7735
rect 7500 7701 7512 7735
rect 10980 7732 11008 7772
rect 11241 7769 11253 7803
rect 11287 7800 11299 7803
rect 11330 7800 11336 7812
rect 11287 7772 11336 7800
rect 11287 7769 11299 7772
rect 11241 7763 11299 7769
rect 11330 7760 11336 7772
rect 11388 7760 11394 7812
rect 13725 7803 13783 7809
rect 13725 7769 13737 7803
rect 13771 7800 13783 7803
rect 15194 7800 15200 7812
rect 13771 7772 13952 7800
rect 13771 7769 13783 7772
rect 13725 7763 13783 7769
rect 13924 7766 13952 7772
rect 14568 7772 15200 7800
rect 14568 7766 14596 7772
rect 11701 7735 11759 7741
rect 7454 7695 7512 7701
rect 7576 7704 10088 7732
rect 10980 7704 11468 7732
rect 7576 7664 7604 7704
rect 10060 7698 10088 7704
rect 10060 7670 10732 7698
rect 7392 7636 7604 7664
rect 10704 7664 10732 7670
rect 10870 7664 10876 7676
rect 10928 7673 10934 7676
rect 11440 7673 11468 7704
rect 11701 7701 11713 7735
rect 11747 7732 11759 7735
rect 12606 7735 12664 7741
rect 12606 7732 12618 7735
rect 11747 7704 12618 7732
rect 11747 7701 11759 7704
rect 11701 7695 11759 7701
rect 12606 7701 12618 7704
rect 12652 7701 12664 7735
rect 12606 7695 12664 7701
rect 13262 7692 13268 7744
rect 13320 7732 13326 7744
rect 13924 7738 14596 7766
rect 15194 7760 15200 7772
rect 15252 7760 15258 7812
rect 16022 7800 16028 7812
rect 15967 7772 16028 7800
rect 16022 7760 16028 7772
rect 16080 7760 16086 7812
rect 18966 7760 18972 7812
rect 19024 7800 19030 7812
rect 21545 7803 21603 7809
rect 21545 7800 21557 7803
rect 19024 7772 19196 7800
rect 19024 7760 19030 7772
rect 19168 7732 19196 7772
rect 19812 7772 21557 7800
rect 19812 7732 19840 7772
rect 21545 7769 21557 7772
rect 21591 7769 21603 7803
rect 21545 7763 21603 7769
rect 13320 7704 13400 7732
rect 19168 7704 19840 7732
rect 20073 7735 20131 7741
rect 13320 7692 13326 7704
rect 10928 7667 10946 7673
rect 10704 7636 10876 7664
rect 10870 7624 10876 7636
rect 10934 7633 10946 7667
rect 10928 7627 10946 7633
rect 11425 7667 11483 7673
rect 11425 7633 11437 7667
rect 11471 7664 11483 7667
rect 11885 7667 11943 7673
rect 11885 7664 11897 7667
rect 11471 7636 11897 7664
rect 11471 7633 11483 7636
rect 11425 7627 11483 7633
rect 11885 7633 11897 7636
rect 11931 7664 11943 7667
rect 12894 7664 12900 7676
rect 11931 7636 12900 7664
rect 11931 7633 11943 7636
rect 11885 7627 11943 7633
rect 10928 7624 10934 7627
rect 12894 7624 12900 7636
rect 12952 7624 12958 7676
rect 8846 7596 8852 7608
rect 8791 7568 8852 7596
rect 8846 7556 8852 7568
rect 8904 7556 8910 7608
rect 9033 7599 9091 7605
rect 9033 7565 9045 7599
rect 9079 7596 9091 7599
rect 10042 7596 10048 7608
rect 9079 7568 10048 7596
rect 9079 7565 9091 7568
rect 9033 7559 9091 7565
rect 5902 7488 5908 7540
rect 5960 7488 5966 7540
rect 6362 7488 6368 7540
rect 6420 7528 6426 7540
rect 9784 7537 9812 7568
rect 10042 7556 10048 7568
rect 10100 7556 10106 7608
rect 11149 7599 11207 7605
rect 11149 7565 11161 7599
rect 11195 7596 11207 7599
rect 12342 7596 12348 7608
rect 11195 7568 12348 7596
rect 11195 7565 11207 7568
rect 11149 7559 11207 7565
rect 12342 7556 12348 7568
rect 12400 7556 12406 7608
rect 13372 7596 13400 7704
rect 20073 7701 20085 7735
rect 20119 7732 20131 7735
rect 20162 7732 20168 7744
rect 20119 7704 20168 7732
rect 20119 7701 20131 7704
rect 20073 7695 20131 7701
rect 20162 7692 20168 7704
rect 20220 7692 20226 7744
rect 22281 7735 22339 7741
rect 22281 7701 22293 7735
rect 22327 7732 22339 7735
rect 23477 7735 23535 7741
rect 23477 7732 23489 7735
rect 22327 7704 22600 7732
rect 22327 7701 22339 7704
rect 22281 7695 22339 7701
rect 13998 7624 14004 7676
rect 14056 7664 14062 7676
rect 14093 7667 14151 7673
rect 14093 7664 14105 7667
rect 14056 7636 14105 7664
rect 14056 7624 14062 7636
rect 14093 7633 14105 7636
rect 14139 7633 14151 7667
rect 14093 7627 14151 7633
rect 14185 7667 14243 7673
rect 14185 7633 14197 7667
rect 14231 7664 14243 7667
rect 14458 7664 14464 7676
rect 14231 7636 14464 7664
rect 14231 7633 14243 7636
rect 14185 7627 14243 7633
rect 14458 7624 14464 7636
rect 14516 7624 14522 7676
rect 14734 7624 14740 7676
rect 14792 7664 14798 7676
rect 18322 7664 18328 7676
rect 14792 7636 18328 7664
rect 14792 7624 14798 7636
rect 18322 7624 18328 7636
rect 18380 7624 18386 7676
rect 18598 7624 18604 7676
rect 18656 7664 18662 7676
rect 18877 7667 18935 7673
rect 18877 7664 18889 7667
rect 18656 7636 18889 7664
rect 18656 7624 18662 7636
rect 18877 7633 18889 7636
rect 18923 7633 18935 7667
rect 18877 7627 18935 7633
rect 19978 7624 19984 7676
rect 20036 7664 20042 7676
rect 20036 7636 20378 7664
rect 20036 7624 20042 7636
rect 22370 7624 22376 7676
rect 22428 7624 22434 7676
rect 22572 7664 22600 7704
rect 23032 7704 23489 7732
rect 23032 7664 23060 7704
rect 23477 7701 23489 7704
rect 23523 7701 23535 7735
rect 23477 7695 23535 7701
rect 22572 7636 23060 7664
rect 14369 7599 14427 7605
rect 14369 7596 14381 7599
rect 13372 7568 14381 7596
rect 14369 7565 14381 7568
rect 14415 7565 14427 7599
rect 14369 7559 14427 7565
rect 17126 7556 17132 7608
rect 17184 7596 17190 7608
rect 17313 7599 17371 7605
rect 17184 7568 17245 7596
rect 17184 7556 17190 7568
rect 17313 7565 17325 7599
rect 17359 7596 17371 7599
rect 17402 7596 17408 7608
rect 17359 7568 17408 7596
rect 17359 7565 17371 7568
rect 17313 7559 17371 7565
rect 17402 7556 17408 7568
rect 17460 7556 17466 7608
rect 18046 7556 18052 7608
rect 18104 7596 18110 7608
rect 20254 7596 20260 7608
rect 18104 7568 20260 7596
rect 18104 7556 18110 7568
rect 20254 7556 20260 7568
rect 20312 7596 20318 7608
rect 20312 7568 20470 7596
rect 20312 7556 20318 7568
rect 21542 7556 21548 7608
rect 21600 7596 21606 7608
rect 22097 7599 22155 7605
rect 22097 7596 22109 7599
rect 21600 7568 22109 7596
rect 21600 7556 21606 7568
rect 22097 7565 22109 7568
rect 22143 7596 22155 7599
rect 22388 7596 22416 7624
rect 22143 7568 22416 7596
rect 22143 7565 22155 7568
rect 22097 7559 22155 7565
rect 6457 7531 6515 7537
rect 6457 7528 6469 7531
rect 6420 7500 6469 7528
rect 6420 7488 6426 7500
rect 6457 7497 6469 7500
rect 6503 7497 6515 7531
rect 6457 7491 6515 7497
rect 9769 7531 9827 7537
rect 9769 7497 9781 7531
rect 9815 7497 9827 7531
rect 11606 7528 11612 7540
rect 11551 7500 11612 7528
rect 9769 7491 9827 7497
rect 11606 7488 11612 7500
rect 11664 7488 11670 7540
rect 14277 7531 14335 7537
rect 14277 7497 14289 7531
rect 14323 7528 14335 7531
rect 16574 7528 16580 7540
rect 14323 7500 16580 7528
rect 14323 7497 14335 7500
rect 14277 7491 14335 7497
rect 16574 7488 16580 7500
rect 16632 7488 16638 7540
rect 5721 7463 5779 7469
rect 5721 7429 5733 7463
rect 5767 7460 5779 7463
rect 5920 7460 5948 7488
rect 5767 7432 5948 7460
rect 5767 7429 5779 7432
rect 5721 7423 5779 7429
rect 5736 7120 5764 7423
rect 6086 7420 6092 7472
rect 6144 7460 6150 7472
rect 8573 7463 8631 7469
rect 8573 7460 8585 7463
rect 6144 7432 8585 7460
rect 6144 7420 6150 7432
rect 8573 7429 8585 7432
rect 8619 7460 8631 7463
rect 9122 7460 9128 7472
rect 8619 7432 9128 7460
rect 8619 7429 8631 7432
rect 8573 7423 8631 7429
rect 9122 7420 9128 7432
rect 9180 7420 9186 7472
rect 12161 7463 12219 7469
rect 12161 7429 12173 7463
rect 12207 7460 12219 7463
rect 12526 7460 12532 7472
rect 12207 7432 12532 7460
rect 12207 7429 12219 7432
rect 12161 7423 12219 7429
rect 12526 7420 12532 7432
rect 12584 7420 12590 7472
rect 13078 7420 13084 7472
rect 13136 7460 13142 7472
rect 13725 7463 13783 7469
rect 13725 7460 13737 7463
rect 13136 7432 13737 7460
rect 13136 7420 13142 7432
rect 13725 7429 13737 7432
rect 13771 7429 13783 7463
rect 13725 7423 13783 7429
rect 18138 7420 18144 7472
rect 18196 7460 18202 7472
rect 18340 7466 19656 7494
rect 19794 7488 19800 7540
rect 19852 7528 19858 7540
rect 19889 7531 19947 7537
rect 19889 7528 19901 7531
rect 19852 7500 19901 7528
rect 19852 7488 19858 7500
rect 19889 7497 19901 7500
rect 19935 7497 19947 7531
rect 21200 7531 21258 7537
rect 21200 7528 21212 7531
rect 19889 7491 19947 7497
rect 21008 7500 21212 7528
rect 21008 7494 21036 7500
rect 18340 7460 18368 7466
rect 18196 7432 18368 7460
rect 19628 7460 19656 7466
rect 20364 7466 21036 7494
rect 21200 7497 21212 7500
rect 21246 7497 21258 7531
rect 21200 7491 21258 7497
rect 21913 7531 21971 7537
rect 21913 7497 21925 7531
rect 21959 7528 21971 7531
rect 22002 7528 22008 7540
rect 21959 7500 22008 7528
rect 21959 7497 21971 7500
rect 21913 7491 21971 7497
rect 22002 7488 22008 7500
rect 22060 7488 22066 7540
rect 20364 7460 20392 7466
rect 19628 7432 20392 7460
rect 18196 7420 18202 7432
rect 5796 7296 23000 7392
rect 5997 7259 6055 7265
rect 5997 7225 6009 7259
rect 6043 7256 6055 7259
rect 6086 7256 6092 7268
rect 6043 7228 6092 7256
rect 6043 7225 6055 7228
rect 5997 7219 6055 7225
rect 6086 7216 6092 7228
rect 6144 7216 6150 7268
rect 6362 7256 6368 7268
rect 6307 7228 6368 7256
rect 6362 7216 6368 7228
rect 6420 7216 6426 7268
rect 13170 7216 13176 7268
rect 13228 7256 13234 7268
rect 13228 7228 14688 7256
rect 13228 7216 13234 7228
rect 12158 7188 12164 7200
rect 12216 7197 12222 7200
rect 12216 7191 12242 7197
rect 12123 7160 12164 7188
rect 12158 7148 12164 7160
rect 12230 7157 12242 7191
rect 12216 7151 12242 7157
rect 12216 7148 12222 7151
rect 5905 7123 5963 7129
rect 5905 7120 5917 7123
rect 5552 7092 5917 7120
rect 5552 7061 5580 7092
rect 5905 7089 5917 7092
rect 5951 7089 5963 7123
rect 6914 7120 6920 7132
rect 6859 7092 6920 7120
rect 5905 7083 5963 7089
rect 6914 7080 6920 7092
rect 6972 7080 6978 7132
rect 12526 7120 12532 7132
rect 10980 7092 11454 7120
rect 12471 7092 12532 7120
rect 9312 7064 9364 7070
rect 5537 7055 5595 7061
rect 5537 7021 5549 7055
rect 5583 7021 5595 7055
rect 5537 7015 5595 7021
rect 6181 7055 6239 7061
rect 6181 7021 6193 7055
rect 6227 7021 6239 7055
rect 9309 7052 9312 7061
rect 9248 7024 9312 7052
rect 6181 7015 6239 7021
rect 9309 7015 9312 7024
rect 5629 6919 5687 6925
rect 5629 6885 5641 6919
rect 5675 6916 5687 6919
rect 6196 6916 6224 7015
rect 9364 7015 9367 7061
rect 9312 7006 9364 7012
rect 7006 6944 7012 6996
rect 7064 6984 7070 6996
rect 7178 6987 7236 6993
rect 7178 6984 7190 6987
rect 7064 6956 7190 6984
rect 7064 6944 7070 6956
rect 7178 6953 7190 6956
rect 7224 6953 7236 6987
rect 10226 6984 10232 6996
rect 7178 6947 7236 6953
rect 7668 6956 8156 6984
rect 6457 6919 6515 6925
rect 6457 6916 6469 6919
rect 5675 6888 6469 6916
rect 5675 6885 5687 6888
rect 5629 6879 5687 6885
rect 6457 6885 6469 6888
rect 6503 6885 6515 6919
rect 6457 6879 6515 6885
rect 6549 6919 6607 6925
rect 6549 6885 6561 6919
rect 6595 6916 6607 6919
rect 6822 6916 6828 6928
rect 6595 6888 6828 6916
rect 6595 6885 6607 6888
rect 6549 6879 6607 6885
rect 6822 6876 6828 6888
rect 6880 6876 6886 6928
rect 7466 6876 7472 6928
rect 7524 6916 7530 6928
rect 7668 6916 7696 6956
rect 7524 6888 7696 6916
rect 8128 6916 8156 6956
rect 8496 6956 9076 6984
rect 10171 6956 10232 6984
rect 8297 6919 8355 6925
rect 8297 6916 8309 6919
rect 8128 6888 8309 6916
rect 7524 6876 7530 6888
rect 8297 6885 8309 6888
rect 8343 6916 8355 6919
rect 8496 6916 8524 6956
rect 8343 6888 8524 6916
rect 9048 6916 9076 6956
rect 10226 6944 10232 6956
rect 10284 6944 10290 6996
rect 10980 6984 11008 7092
rect 12526 7080 12532 7092
rect 12584 7080 12590 7132
rect 13078 7052 13084 7064
rect 12282 7024 13084 7052
rect 13078 7012 13084 7024
rect 13136 7012 13142 7064
rect 13630 7052 13636 7064
rect 13575 7024 13636 7052
rect 13630 7012 13636 7024
rect 13688 7012 13694 7064
rect 14660 7052 14688 7228
rect 14734 7216 14740 7268
rect 14792 7256 14798 7268
rect 15013 7259 15071 7265
rect 15013 7256 15025 7259
rect 14792 7228 15025 7256
rect 14792 7216 14798 7228
rect 15013 7225 15025 7228
rect 15059 7225 15071 7259
rect 15013 7219 15071 7225
rect 16942 7216 16948 7268
rect 17000 7256 17006 7268
rect 17589 7259 17647 7265
rect 17589 7256 17601 7259
rect 17000 7228 17601 7256
rect 17000 7216 17006 7228
rect 17589 7225 17601 7228
rect 17635 7225 17647 7259
rect 17862 7256 17868 7268
rect 17807 7228 17868 7256
rect 17589 7219 17647 7225
rect 17862 7216 17868 7228
rect 17920 7216 17926 7268
rect 18966 7256 18972 7268
rect 18800 7228 18972 7256
rect 15197 7191 15255 7197
rect 15197 7157 15209 7191
rect 15243 7188 15255 7191
rect 15654 7188 15660 7200
rect 15243 7160 15660 7188
rect 15243 7157 15255 7160
rect 15197 7151 15255 7157
rect 15654 7148 15660 7160
rect 15712 7148 15718 7200
rect 18800 7197 18828 7228
rect 18966 7216 18972 7228
rect 19024 7216 19030 7268
rect 20254 7216 20260 7268
rect 20312 7256 20318 7268
rect 20625 7259 20683 7265
rect 20625 7256 20637 7259
rect 20312 7228 20637 7256
rect 20312 7216 20318 7228
rect 20625 7225 20637 7228
rect 20671 7225 20683 7259
rect 21542 7256 21548 7268
rect 20625 7219 20683 7225
rect 21192 7228 21548 7256
rect 18785 7191 18843 7197
rect 18785 7157 18797 7191
rect 18831 7157 18843 7191
rect 18785 7151 18843 7157
rect 16206 7120 16212 7132
rect 16151 7092 16212 7120
rect 16206 7080 16212 7092
rect 16264 7080 16270 7132
rect 19242 7120 19248 7132
rect 19187 7092 19248 7120
rect 19242 7080 19248 7092
rect 19300 7080 19306 7132
rect 20714 7120 20720 7132
rect 20659 7092 20720 7120
rect 20714 7080 20720 7092
rect 20772 7080 20778 7132
rect 20901 7123 20959 7129
rect 20901 7089 20913 7123
rect 20947 7120 20959 7123
rect 21192 7120 21220 7228
rect 21542 7216 21548 7228
rect 21600 7216 21606 7268
rect 21358 7120 21364 7132
rect 20947 7092 21220 7120
rect 21303 7092 21364 7120
rect 20947 7089 20959 7092
rect 20901 7083 20959 7089
rect 21358 7080 21364 7092
rect 21416 7080 21422 7132
rect 15381 7055 15439 7061
rect 15381 7052 15393 7055
rect 14660 7024 15393 7052
rect 15381 7021 15393 7024
rect 15427 7052 15439 7055
rect 17770 7052 17776 7064
rect 15427 7024 16712 7052
rect 15427 7021 15439 7024
rect 15381 7015 15439 7021
rect 10428 6956 11008 6984
rect 11057 6987 11115 6993
rect 10428 6916 10456 6956
rect 11057 6953 11069 6987
rect 11103 6984 11115 6987
rect 11238 6984 11244 6996
rect 11103 6956 11244 6984
rect 11103 6953 11115 6956
rect 11057 6947 11115 6953
rect 11238 6944 11244 6956
rect 11296 6944 11302 6996
rect 13894 6987 13952 6993
rect 13894 6984 13906 6987
rect 13280 6956 13906 6984
rect 13280 6928 13308 6956
rect 13894 6953 13906 6956
rect 13940 6984 13952 6987
rect 13998 6984 14004 6996
rect 13940 6956 14004 6984
rect 13940 6953 13952 6956
rect 13894 6947 13952 6953
rect 13998 6944 14004 6956
rect 14056 6944 14062 6996
rect 15749 6987 15807 6993
rect 15749 6953 15761 6987
rect 15795 6984 15807 6987
rect 16470 6987 16528 6993
rect 16470 6984 16482 6987
rect 15795 6956 16482 6984
rect 15795 6953 15807 6956
rect 15749 6947 15807 6953
rect 16470 6953 16482 6956
rect 16516 6953 16528 6987
rect 16684 6984 16712 7024
rect 17236 7024 17776 7052
rect 17236 6984 17264 7024
rect 17770 7012 17776 7024
rect 17828 7052 17834 7064
rect 18049 7055 18107 7061
rect 18049 7052 18061 7055
rect 17828 7024 18061 7052
rect 17828 7012 17834 7024
rect 18049 7021 18061 7024
rect 18095 7052 18107 7055
rect 18969 7055 19027 7061
rect 18969 7052 18981 7055
rect 18095 7024 18981 7052
rect 18095 7021 18107 7024
rect 18049 7015 18107 7021
rect 18969 7021 18981 7024
rect 19015 7021 19027 7055
rect 18969 7015 19027 7021
rect 21177 7055 21235 7061
rect 21177 7021 21189 7055
rect 21223 7052 21235 7055
rect 23845 7055 23903 7061
rect 23845 7052 23857 7055
rect 21223 7024 23857 7052
rect 21223 7021 21235 7024
rect 21177 7015 21235 7021
rect 23845 7021 23857 7024
rect 23891 7021 23903 7055
rect 23845 7015 23903 7021
rect 21634 6993 21640 6996
rect 16684 6956 17264 6984
rect 19153 6987 19211 6993
rect 16470 6947 16528 6953
rect 19153 6953 19165 6987
rect 19199 6984 19211 6987
rect 19506 6987 19564 6993
rect 19506 6984 19518 6987
rect 19199 6956 19518 6984
rect 19199 6953 19211 6956
rect 19153 6947 19211 6953
rect 19506 6953 19518 6956
rect 19552 6953 19564 6987
rect 21622 6987 21640 6993
rect 21622 6984 21634 6987
rect 21579 6956 21634 6984
rect 19506 6947 19564 6953
rect 21622 6953 21634 6956
rect 21622 6947 21640 6953
rect 21634 6944 21640 6947
rect 21692 6944 21698 6996
rect 9048 6888 10456 6916
rect 8343 6885 8355 6888
rect 8297 6879 8355 6885
rect 13262 6876 13268 6928
rect 13320 6876 13326 6928
rect 18325 6919 18383 6925
rect 18325 6885 18337 6919
rect 18371 6916 18383 6919
rect 18966 6916 18972 6928
rect 18371 6888 18972 6916
rect 18371 6885 18383 6888
rect 18325 6879 18383 6885
rect 18966 6876 18972 6888
rect 19024 6876 19030 6928
rect 22462 6876 22468 6928
rect 22520 6916 22526 6928
rect 22741 6919 22799 6925
rect 22741 6916 22753 6919
rect 22520 6888 22753 6916
rect 22520 6876 22526 6888
rect 22741 6885 22753 6888
rect 22787 6885 22799 6919
rect 22741 6879 22799 6885
rect 5796 6752 23000 6848
rect 6181 6715 6239 6721
rect 6181 6681 6193 6715
rect 6227 6712 6239 6715
rect 6227 6684 6776 6712
rect 6227 6681 6239 6684
rect 6181 6675 6239 6681
rect 6086 6644 6092 6656
rect 6031 6616 6092 6644
rect 6086 6604 6092 6616
rect 6144 6604 6150 6656
rect 6748 6644 6776 6684
rect 7668 6684 8156 6712
rect 7668 6656 7696 6684
rect 7469 6647 7527 6653
rect 7469 6644 7481 6647
rect 6748 6616 7481 6644
rect 6748 6585 6776 6616
rect 7469 6613 7481 6616
rect 7515 6613 7527 6647
rect 7650 6644 7656 6656
rect 7595 6616 7656 6644
rect 7469 6607 7527 6613
rect 7650 6604 7656 6616
rect 7708 6604 7714 6656
rect 7834 6644 7840 6656
rect 7779 6616 7840 6644
rect 7834 6604 7840 6616
rect 7892 6604 7898 6656
rect 8128 6593 8156 6684
rect 11606 6672 11612 6724
rect 11664 6712 11670 6724
rect 12069 6715 12127 6721
rect 12069 6712 12081 6715
rect 11664 6684 12081 6712
rect 11664 6672 11670 6684
rect 12069 6681 12081 6684
rect 12115 6681 12127 6715
rect 12069 6675 12127 6681
rect 13262 6672 13268 6724
rect 13320 6712 13326 6724
rect 13725 6715 13783 6721
rect 13725 6712 13737 6715
rect 13320 6684 13737 6712
rect 13320 6672 13326 6684
rect 13725 6681 13737 6684
rect 13771 6681 13783 6715
rect 13725 6675 13783 6681
rect 20165 6715 20223 6721
rect 20165 6681 20177 6715
rect 20211 6712 20223 6715
rect 20714 6712 20720 6724
rect 20211 6684 20720 6712
rect 20211 6681 20223 6684
rect 20165 6675 20223 6681
rect 20714 6672 20720 6684
rect 20772 6672 20778 6724
rect 22281 6715 22339 6721
rect 22281 6681 22293 6715
rect 22327 6712 22339 6715
rect 23661 6715 23719 6721
rect 23661 6712 23673 6715
rect 22327 6684 23673 6712
rect 22327 6681 22339 6684
rect 22281 6675 22339 6681
rect 23661 6681 23673 6684
rect 23707 6681 23719 6715
rect 23661 6675 23719 6681
rect 10410 6604 10416 6656
rect 10468 6644 10474 6656
rect 10597 6647 10655 6653
rect 10597 6644 10609 6647
rect 10468 6616 10609 6644
rect 10468 6604 10474 6616
rect 10597 6613 10609 6616
rect 10643 6613 10655 6647
rect 10597 6607 10655 6613
rect 13814 6604 13820 6656
rect 13872 6644 13878 6656
rect 15182 6647 15240 6653
rect 15182 6644 15194 6647
rect 13872 6616 14044 6644
rect 13872 6604 13878 6616
rect 6733 6579 6791 6585
rect 6733 6545 6745 6579
rect 6779 6545 6791 6579
rect 6733 6539 6791 6545
rect 6822 6536 6828 6588
rect 6880 6576 6886 6588
rect 8113 6587 8171 6593
rect 7009 6579 7067 6585
rect 7009 6576 7021 6579
rect 6880 6548 7021 6576
rect 6880 6536 6886 6548
rect 7009 6545 7021 6548
rect 7055 6545 7067 6579
rect 7009 6539 7067 6545
rect 7561 6579 7619 6585
rect 7561 6545 7573 6579
rect 7607 6576 7619 6579
rect 7929 6579 7987 6585
rect 7929 6576 7941 6579
rect 7607 6548 7941 6576
rect 7607 6545 7619 6548
rect 7561 6539 7619 6545
rect 7929 6545 7941 6548
rect 7975 6545 7987 6579
rect 8113 6553 8125 6587
rect 8159 6553 8171 6587
rect 8478 6585 8484 6588
rect 8466 6579 8484 6585
rect 8466 6576 8478 6579
rect 8113 6547 8171 6553
rect 8423 6548 8478 6576
rect 7929 6539 7987 6545
rect 8466 6545 8478 6548
rect 8466 6539 8484 6545
rect 8478 6536 8484 6539
rect 8536 6536 8542 6588
rect 11974 6576 11980 6588
rect 11822 6548 11980 6576
rect 11974 6536 11980 6548
rect 12032 6536 12038 6588
rect 12342 6576 12348 6588
rect 12287 6548 12348 6576
rect 12342 6536 12348 6548
rect 12400 6536 12406 6588
rect 12606 6579 12664 6585
rect 12606 6576 12618 6579
rect 12452 6548 12618 6576
rect 6365 6511 6423 6517
rect 6365 6477 6377 6511
rect 6411 6508 6423 6511
rect 6917 6511 6975 6517
rect 6917 6508 6929 6511
rect 6411 6480 6929 6508
rect 6411 6477 6423 6480
rect 6365 6471 6423 6477
rect 6917 6477 6929 6480
rect 6963 6508 6975 6511
rect 7466 6508 7472 6520
rect 6963 6480 7472 6508
rect 6963 6477 6975 6480
rect 6917 6471 6975 6477
rect 7466 6468 7472 6480
rect 7524 6468 7530 6520
rect 7834 6468 7840 6520
rect 7892 6508 7898 6520
rect 8021 6511 8079 6517
rect 8021 6508 8033 6511
rect 7892 6480 8033 6508
rect 7892 6468 7898 6480
rect 8021 6477 8033 6480
rect 8067 6477 8079 6511
rect 8021 6471 8079 6477
rect 8202 6468 8208 6520
rect 8260 6508 8266 6520
rect 10318 6508 10324 6520
rect 8260 6480 8321 6508
rect 9876 6480 10324 6508
rect 8260 6468 8266 6480
rect 9585 6443 9643 6449
rect 9585 6409 9597 6443
rect 9631 6440 9643 6443
rect 9876 6440 9904 6480
rect 10318 6468 10324 6480
rect 10376 6508 10382 6520
rect 12452 6508 12480 6548
rect 12606 6545 12618 6548
rect 12652 6545 12664 6579
rect 14016 6576 14044 6616
rect 14476 6616 15194 6644
rect 14476 6576 14504 6616
rect 15182 6613 15194 6616
rect 15228 6613 15240 6647
rect 22922 6644 22928 6656
rect 15182 6607 15240 6613
rect 21744 6616 22232 6644
rect 14016 6548 14504 6576
rect 12606 6539 12664 6545
rect 14642 6536 14648 6588
rect 14700 6576 14706 6588
rect 14921 6579 14979 6585
rect 14921 6576 14933 6579
rect 14700 6548 14933 6576
rect 14700 6536 14706 6548
rect 14921 6545 14933 6548
rect 14967 6545 14979 6579
rect 18322 6576 18328 6588
rect 18267 6548 18328 6576
rect 14921 6539 14979 6545
rect 18322 6536 18328 6548
rect 18380 6536 18386 6588
rect 20809 6579 20867 6585
rect 20809 6545 20821 6579
rect 20855 6576 20867 6579
rect 20990 6576 20996 6588
rect 20855 6548 20996 6576
rect 20855 6545 20867 6548
rect 20809 6539 20867 6545
rect 20990 6536 20996 6548
rect 21048 6536 21054 6588
rect 21637 6579 21695 6585
rect 21637 6545 21649 6579
rect 21683 6576 21695 6579
rect 21744 6576 21772 6616
rect 21683 6548 21772 6576
rect 21683 6545 21695 6548
rect 21637 6539 21695 6545
rect 21818 6536 21824 6588
rect 21876 6576 21882 6588
rect 21913 6579 21971 6585
rect 21913 6576 21925 6579
rect 21876 6548 21925 6576
rect 21876 6536 21882 6548
rect 21913 6545 21925 6548
rect 21959 6545 21971 6579
rect 22204 6576 22232 6616
rect 22756 6616 22928 6644
rect 22756 6576 22784 6616
rect 22922 6604 22928 6616
rect 22980 6604 22986 6656
rect 22204 6548 22784 6576
rect 21913 6539 21971 6545
rect 18598 6508 18604 6520
rect 10376 6480 10994 6508
rect 11992 6480 12480 6508
rect 18543 6480 18604 6508
rect 10376 6468 10382 6480
rect 9631 6412 9904 6440
rect 9631 6409 9643 6412
rect 9585 6403 9643 6409
rect 6546 6372 6552 6384
rect 6491 6344 6552 6372
rect 6546 6332 6552 6344
rect 6604 6332 6610 6384
rect 7742 6332 7748 6384
rect 7800 6372 7806 6384
rect 7837 6375 7895 6381
rect 7837 6372 7849 6375
rect 7800 6344 7849 6372
rect 7800 6332 7806 6344
rect 7837 6341 7849 6344
rect 7883 6341 7895 6375
rect 7837 6335 7895 6341
rect 9950 6332 9956 6384
rect 10008 6372 10014 6384
rect 10152 6378 11100 6406
rect 11238 6400 11244 6452
rect 11296 6440 11302 6452
rect 11724 6443 11782 6449
rect 11724 6440 11736 6443
rect 11296 6412 11736 6440
rect 11296 6400 11302 6412
rect 11724 6409 11736 6412
rect 11770 6409 11782 6443
rect 11724 6403 11782 6409
rect 10152 6372 10180 6378
rect 10008 6344 10180 6372
rect 11072 6372 11100 6378
rect 11992 6372 12020 6480
rect 18598 6468 18604 6480
rect 18656 6468 18662 6520
rect 19794 6468 19800 6520
rect 19852 6508 19858 6520
rect 20533 6511 20591 6517
rect 20533 6508 20545 6511
rect 19852 6480 20545 6508
rect 19852 6468 19858 6480
rect 20533 6477 20545 6480
rect 20579 6477 20591 6511
rect 20533 6471 20591 6477
rect 20993 6443 21051 6449
rect 20993 6409 21005 6443
rect 21039 6440 21051 6443
rect 21192 6446 21956 6474
rect 21192 6440 21220 6446
rect 21039 6412 21220 6440
rect 21928 6440 21956 6446
rect 24029 6443 24087 6449
rect 24029 6440 24041 6443
rect 21928 6412 24041 6440
rect 21039 6409 21051 6412
rect 20993 6403 21051 6409
rect 24029 6409 24041 6412
rect 24075 6409 24087 6443
rect 24029 6403 24087 6409
rect 11072 6344 12020 6372
rect 10008 6332 10014 6344
rect 16206 6332 16212 6384
rect 16264 6372 16270 6384
rect 16301 6375 16359 6381
rect 16301 6372 16313 6375
rect 16264 6344 16313 6372
rect 16264 6332 16270 6344
rect 16301 6341 16313 6344
rect 16347 6341 16359 6375
rect 16301 6335 16359 6341
rect 21453 6375 21511 6381
rect 21453 6341 21465 6375
rect 21499 6372 21511 6375
rect 21818 6372 21824 6384
rect 21499 6344 21824 6372
rect 21499 6341 21511 6344
rect 21453 6335 21511 6341
rect 21818 6332 21824 6344
rect 21876 6332 21882 6384
rect 5796 6208 23000 6304
rect 6917 6171 6975 6177
rect 6917 6137 6929 6171
rect 6963 6168 6975 6171
rect 7006 6168 7012 6180
rect 6963 6140 7012 6168
rect 6963 6137 6975 6140
rect 6917 6131 6975 6137
rect 7006 6128 7012 6140
rect 7064 6128 7070 6180
rect 7742 6168 7748 6180
rect 7687 6140 7748 6168
rect 7742 6128 7748 6140
rect 7800 6128 7806 6180
rect 8205 6171 8263 6177
rect 8205 6137 8217 6171
rect 8251 6168 8263 6171
rect 8386 6168 8392 6180
rect 8251 6140 8392 6168
rect 8251 6137 8263 6140
rect 8205 6131 8263 6137
rect 8386 6128 8392 6140
rect 8444 6128 8450 6180
rect 9122 6128 9128 6180
rect 9180 6128 9186 6180
rect 10318 6128 10324 6180
rect 10376 6168 10382 6180
rect 10413 6171 10471 6177
rect 10413 6168 10425 6171
rect 10376 6140 10425 6168
rect 10376 6128 10382 6140
rect 10413 6137 10425 6140
rect 10459 6137 10471 6171
rect 10413 6131 10471 6137
rect 12250 6128 12256 6180
rect 12308 6168 12314 6180
rect 12345 6171 12403 6177
rect 12345 6168 12357 6171
rect 12308 6140 12357 6168
rect 12308 6128 12314 6140
rect 12345 6137 12357 6140
rect 12391 6137 12403 6171
rect 12345 6131 12403 6137
rect 13173 6171 13231 6177
rect 13173 6137 13185 6171
rect 13219 6168 13231 6171
rect 13814 6168 13820 6180
rect 13219 6140 13820 6168
rect 13219 6137 13231 6140
rect 13173 6131 13231 6137
rect 13814 6128 13820 6140
rect 13872 6128 13878 6180
rect 18049 6171 18107 6177
rect 18049 6137 18061 6171
rect 18095 6168 18107 6171
rect 18782 6168 18788 6180
rect 18095 6140 18788 6168
rect 18095 6137 18107 6140
rect 18049 6131 18107 6137
rect 18782 6128 18788 6140
rect 18840 6128 18846 6180
rect 18966 6168 18972 6180
rect 18911 6140 18972 6168
rect 18966 6128 18972 6140
rect 19024 6128 19030 6180
rect 19794 6168 19800 6180
rect 19739 6140 19800 6168
rect 19794 6128 19800 6140
rect 19852 6128 19858 6180
rect 21085 6171 21143 6177
rect 21085 6137 21097 6171
rect 21131 6168 21143 6171
rect 21131 6140 21956 6168
rect 21131 6137 21143 6140
rect 21085 6131 21143 6137
rect 9140 6100 9168 6128
rect 16206 6100 16212 6112
rect 9140 6072 10272 6100
rect 10244 6066 10272 6072
rect 12360 6072 13492 6100
rect 6546 6032 6552 6044
rect 6491 6004 6552 6032
rect 6546 5992 6552 6004
rect 6604 5992 6610 6044
rect 7650 5992 7656 6044
rect 7708 6032 7714 6044
rect 10244 6038 10824 6066
rect 10796 6032 10824 6038
rect 12360 6032 12388 6072
rect 12544 6041 12572 6072
rect 7708 6004 8156 6032
rect 10796 6004 12388 6032
rect 12529 6035 12587 6041
rect 7708 5992 7714 6004
rect 6730 5924 6736 5976
rect 6788 5964 6794 5976
rect 8021 5967 8079 5973
rect 8021 5964 8033 5967
rect 6788 5936 8033 5964
rect 6788 5924 6794 5936
rect 8021 5933 8033 5936
rect 8067 5933 8079 5967
rect 8128 5964 8156 6004
rect 12529 6001 12541 6035
rect 12575 6001 12587 6035
rect 12529 5995 12587 6001
rect 12713 6035 12771 6041
rect 12713 6001 12725 6035
rect 12759 6001 12771 6035
rect 12713 5995 12771 6001
rect 12805 6035 12863 6041
rect 12805 6001 12817 6035
rect 12851 6032 12863 6035
rect 13357 6035 13415 6041
rect 13357 6032 13369 6035
rect 12851 6004 13369 6032
rect 12851 6001 12863 6004
rect 12805 5995 12863 6001
rect 13357 6001 13369 6004
rect 13403 6001 13415 6035
rect 13357 5995 13415 6001
rect 10597 5967 10655 5973
rect 10597 5964 10609 5967
rect 8128 5936 10609 5964
rect 8021 5927 8079 5933
rect 10597 5933 10609 5936
rect 10643 5933 10655 5967
rect 10597 5927 10655 5933
rect 12728 5896 12756 5995
rect 12894 5924 12900 5976
rect 12952 5964 12958 5976
rect 12989 5967 13047 5973
rect 12989 5964 13001 5967
rect 12952 5936 13001 5964
rect 12952 5924 12958 5936
rect 12989 5933 13001 5936
rect 13035 5933 13047 5967
rect 13262 5964 13268 5976
rect 13207 5936 13268 5964
rect 12989 5927 13047 5933
rect 13262 5924 13268 5936
rect 13320 5924 13326 5976
rect 13464 5964 13492 6072
rect 13924 6072 14504 6100
rect 13924 5973 13952 6072
rect 14274 6032 14280 6044
rect 14219 6004 14280 6032
rect 14274 5992 14280 6004
rect 14332 5992 14338 6044
rect 14476 6032 14504 6072
rect 16040 6072 16212 6100
rect 16040 6032 16068 6072
rect 16206 6060 16212 6072
rect 16264 6100 16270 6112
rect 16393 6103 16451 6109
rect 16264 6072 16344 6100
rect 16264 6060 16270 6072
rect 14476 6004 16068 6032
rect 16316 6032 16344 6072
rect 16393 6069 16405 6103
rect 16439 6100 16451 6103
rect 20257 6103 20315 6109
rect 20257 6100 20269 6103
rect 16439 6072 16712 6100
rect 16439 6069 16451 6072
rect 16393 6063 16451 6069
rect 16577 6035 16635 6041
rect 16577 6032 16589 6035
rect 16316 6004 16589 6032
rect 16577 6001 16589 6004
rect 16623 6001 16635 6035
rect 16684 6032 16712 6072
rect 19536 6072 20269 6100
rect 18138 6032 18144 6044
rect 16684 6004 18144 6032
rect 16577 5995 16635 6001
rect 18138 5992 18144 6004
rect 18196 5992 18202 6044
rect 19536 6041 19564 6072
rect 20257 6069 20269 6072
rect 20303 6069 20315 6103
rect 21545 6103 21603 6109
rect 21545 6100 21557 6103
rect 20257 6063 20315 6069
rect 20732 6072 21557 6100
rect 19521 6035 19579 6041
rect 19521 6001 19533 6035
rect 19567 6001 19579 6035
rect 19521 5995 19579 6001
rect 20070 5992 20076 6044
rect 20128 6032 20134 6044
rect 20732 6041 20760 6072
rect 21545 6069 21557 6072
rect 21591 6069 21603 6103
rect 21928 6100 21956 6140
rect 22002 6128 22008 6180
rect 22060 6168 22066 6180
rect 22373 6171 22431 6177
rect 22373 6168 22385 6171
rect 22060 6140 22385 6168
rect 22060 6128 22066 6140
rect 22373 6137 22385 6140
rect 22419 6137 22431 6171
rect 22373 6131 22431 6137
rect 22186 6100 22192 6112
rect 21928 6072 22192 6100
rect 21545 6063 21603 6069
rect 22186 6060 22192 6072
rect 22244 6060 22250 6112
rect 20441 6035 20499 6041
rect 20441 6032 20453 6035
rect 20128 6004 20453 6032
rect 20128 5992 20134 6004
rect 20441 6001 20453 6004
rect 20487 6001 20499 6035
rect 20441 5995 20499 6001
rect 20717 6035 20775 6041
rect 20717 6001 20729 6035
rect 20763 6001 20775 6035
rect 20717 5995 20775 6001
rect 21266 5992 21272 6044
rect 21324 6032 21330 6044
rect 21729 6035 21787 6041
rect 21729 6032 21741 6035
rect 21324 6004 21741 6032
rect 21324 5992 21330 6004
rect 21729 6001 21741 6004
rect 21775 6001 21787 6035
rect 21729 5995 21787 6001
rect 21818 5992 21824 6044
rect 21876 6032 21882 6044
rect 21876 6004 21937 6032
rect 21876 5992 21882 6004
rect 13725 5967 13783 5973
rect 13725 5964 13737 5967
rect 13464 5936 13737 5964
rect 13725 5933 13737 5936
rect 13771 5933 13783 5967
rect 13909 5967 13967 5973
rect 13909 5964 13921 5967
rect 13725 5927 13783 5933
rect 13832 5936 13921 5964
rect 13832 5896 13860 5936
rect 13909 5933 13921 5936
rect 13955 5933 13967 5967
rect 13909 5927 13967 5933
rect 14090 5967 14154 5973
rect 14090 5933 14105 5967
rect 14139 5933 14154 5967
rect 16850 5964 16856 5976
rect 16795 5936 16856 5964
rect 12728 5868 12940 5896
rect 12912 5862 12940 5868
rect 13648 5868 13860 5896
rect 14090 5908 14154 5933
rect 16850 5924 16856 5936
rect 16908 5924 16914 5976
rect 17770 5964 17776 5976
rect 17715 5936 17776 5964
rect 17770 5924 17776 5936
rect 17828 5924 17834 5976
rect 19613 5967 19671 5973
rect 19613 5933 19625 5967
rect 19659 5964 19671 5967
rect 20346 5964 20352 5976
rect 19659 5936 20352 5964
rect 19659 5933 19671 5936
rect 19613 5927 19671 5933
rect 20346 5924 20352 5936
rect 20404 5924 20410 5976
rect 13648 5862 13676 5868
rect 12912 5834 13676 5862
rect 14090 5856 14096 5908
rect 14148 5856 14154 5908
rect 5796 5664 23000 5760
rect 10870 4156 10876 4208
rect 10928 4196 10934 4208
rect 10928 4168 19196 4196
rect 10928 4156 10934 4168
rect 19168 4140 19196 4168
rect 19150 4088 19156 4140
rect 19208 4088 19214 4140
rect 14 144 20 196
rect 72 184 78 196
rect 72 156 2636 184
rect 72 144 78 156
rect 2608 116 2636 156
rect 13446 144 13452 196
rect 13504 144 13510 196
rect 13464 116 13492 144
rect 2608 88 13492 116
<< via1 >>
rect 15936 21768 15988 21820
rect 10324 21743 10376 21752
rect 10324 21709 10333 21743
rect 10333 21709 10367 21743
rect 10367 21709 10376 21743
rect 10324 21700 10376 21709
rect 14280 21700 14332 21752
rect 16488 21700 16540 21752
rect 18236 21768 18288 21820
rect 19616 21700 19668 21752
rect 10140 21675 10192 21684
rect 10140 21641 10149 21675
rect 10149 21641 10183 21675
rect 10183 21641 10192 21675
rect 10140 21632 10192 21641
rect 10508 21607 10560 21616
rect 10508 21573 10517 21607
rect 10517 21573 10551 21607
rect 10551 21573 10560 21607
rect 10508 21564 10560 21573
rect 15476 21564 15528 21616
rect 18420 21632 18472 21684
rect 21272 21768 21324 21820
rect 22744 21768 22796 21820
rect 20352 21700 20404 21752
rect 21088 21700 21140 21752
rect 22008 21743 22060 21752
rect 22008 21709 22017 21743
rect 22017 21709 22051 21743
rect 22051 21709 22060 21743
rect 22008 21700 22060 21709
rect 17408 21564 17460 21616
rect 19156 21607 19208 21616
rect 19156 21573 19165 21607
rect 19165 21573 19199 21607
rect 19199 21573 19208 21607
rect 19156 21564 19208 21573
rect 19892 21607 19944 21616
rect 19892 21573 19901 21607
rect 19901 21573 19935 21607
rect 19935 21573 19944 21607
rect 19892 21564 19944 21573
rect 19984 21564 20036 21616
rect 21640 21564 21692 21616
rect 22376 21607 22428 21616
rect 22376 21573 22385 21607
rect 22385 21573 22419 21607
rect 22419 21573 22428 21607
rect 22376 21564 22428 21573
rect 10140 21403 10192 21412
rect 10140 21369 10149 21403
rect 10149 21369 10183 21403
rect 10183 21369 10192 21403
rect 10140 21360 10192 21369
rect 15936 21403 15988 21412
rect 15936 21369 15945 21403
rect 15945 21369 15979 21403
rect 15979 21369 15988 21403
rect 15936 21360 15988 21369
rect 18236 21360 18288 21412
rect 17132 21292 17184 21344
rect 19156 21292 19208 21344
rect 19984 21360 20036 21412
rect 22008 21360 22060 21412
rect 22192 21292 22244 21344
rect 10968 21156 11020 21208
rect 13084 21156 13136 21208
rect 13360 21156 13412 21208
rect 14464 21156 14516 21208
rect 15108 21156 15160 21208
rect 16488 21224 16540 21276
rect 17408 21267 17460 21276
rect 17408 21233 17417 21267
rect 17417 21233 17451 21267
rect 17451 21233 17460 21267
rect 17408 21224 17460 21233
rect 15936 21156 15988 21208
rect 19616 21224 19668 21276
rect 21456 21224 21508 21276
rect 14280 21088 14332 21140
rect 16120 21088 16172 21140
rect 20076 21156 20128 21208
rect 21272 21199 21324 21208
rect 21272 21165 21281 21199
rect 21281 21165 21315 21199
rect 21315 21165 21324 21199
rect 21272 21156 21324 21165
rect 18420 21088 18472 21140
rect 9956 21020 10008 21072
rect 12624 21020 12676 21072
rect 14372 21063 14424 21072
rect 14372 21029 14381 21063
rect 14381 21029 14415 21063
rect 14415 21029 14424 21063
rect 14372 21020 14424 21029
rect 14740 21020 14792 21072
rect 16212 21063 16264 21072
rect 16212 21029 16221 21063
rect 16221 21029 16255 21063
rect 16255 21029 16264 21063
rect 16212 21020 16264 21029
rect 17684 21020 17736 21072
rect 18880 21063 18932 21072
rect 18880 21029 18889 21063
rect 18889 21029 18923 21063
rect 18923 21029 18932 21063
rect 18880 21020 18932 21029
rect 10891 20816 10943 20868
rect 12609 20816 12661 20868
rect 14280 20859 14332 20868
rect 14280 20825 14289 20859
rect 14289 20825 14323 20859
rect 14323 20825 14332 20859
rect 14280 20816 14332 20825
rect 15476 20816 15528 20868
rect 20444 20816 20496 20868
rect 13084 20748 13136 20800
rect 16212 20791 16264 20800
rect 7564 20723 7616 20732
rect 7564 20689 7592 20723
rect 7592 20689 7616 20723
rect 7564 20680 7616 20689
rect 10876 20680 10928 20732
rect 12624 20680 12676 20732
rect 16212 20757 16240 20791
rect 16240 20757 16264 20791
rect 16212 20748 16264 20757
rect 18880 20791 18932 20800
rect 18880 20757 18904 20791
rect 18904 20757 18932 20791
rect 18880 20748 18932 20757
rect 19892 20748 19944 20800
rect 15108 20723 15160 20732
rect 7288 20655 7340 20664
rect 7288 20621 7297 20655
rect 7297 20621 7331 20655
rect 7331 20621 7340 20655
rect 7288 20612 7340 20621
rect 11520 20544 11572 20596
rect 14464 20612 14516 20664
rect 9128 20476 9180 20528
rect 9956 20476 10008 20528
rect 13360 20476 13412 20528
rect 15108 20689 15117 20723
rect 15117 20689 15151 20723
rect 15151 20689 15160 20723
rect 15108 20680 15160 20689
rect 22560 20680 22612 20732
rect 15936 20655 15988 20664
rect 15936 20621 15945 20655
rect 15945 20621 15979 20655
rect 15979 20621 15988 20655
rect 15936 20612 15988 20621
rect 19156 20655 19208 20664
rect 19156 20621 19165 20655
rect 19165 20621 19199 20655
rect 19199 20621 19208 20655
rect 19156 20612 19208 20621
rect 20076 20655 20128 20664
rect 20076 20621 20085 20655
rect 20085 20621 20119 20655
rect 20119 20621 20128 20655
rect 20076 20612 20128 20621
rect 22008 20612 22060 20664
rect 15476 20476 15528 20528
rect 17132 20476 17184 20528
rect 17684 20476 17736 20528
rect 10324 20272 10376 20324
rect 6828 20179 6880 20188
rect 6828 20145 6837 20179
rect 6837 20145 6871 20179
rect 6871 20145 6880 20179
rect 6828 20136 6880 20145
rect 10692 20136 10744 20188
rect 22928 20179 22980 20188
rect 22928 20145 22937 20179
rect 22937 20145 22971 20179
rect 22971 20145 22980 20179
rect 22928 20136 22980 20145
rect 12624 20068 12676 20120
rect 15936 20068 15988 20120
rect 20076 20068 20128 20120
rect 6920 20000 6972 20052
rect 10232 20043 10284 20052
rect 6736 19932 6788 19984
rect 10232 20009 10256 20043
rect 10256 20009 10284 20043
rect 10232 20000 10284 20009
rect 12348 20000 12400 20052
rect 15476 20000 15528 20052
rect 16304 20000 16356 20052
rect 8760 19932 8812 19984
rect 8944 19932 8996 19984
rect 13452 19932 13504 19984
rect 14740 19932 14792 19984
rect 16028 19932 16080 19984
rect 17868 19932 17920 19984
rect 18880 20000 18932 20052
rect 20168 19932 20220 19984
rect 22928 20000 22980 20052
rect 7564 19728 7616 19780
rect 8944 19728 8996 19780
rect 9128 19771 9180 19780
rect 9128 19737 9137 19771
rect 9137 19737 9171 19771
rect 9171 19737 9180 19771
rect 9128 19728 9180 19737
rect 10232 19728 10284 19780
rect 16120 19728 16172 19780
rect 16304 19771 16356 19780
rect 16304 19737 16313 19771
rect 16313 19737 16347 19771
rect 16347 19737 16356 19771
rect 16304 19728 16356 19737
rect 8760 19660 8812 19712
rect 18880 19728 18932 19780
rect 22008 19728 22060 19780
rect 7012 19592 7064 19644
rect 10508 19635 10560 19644
rect 10508 19601 10517 19635
rect 10517 19601 10551 19635
rect 10551 19601 10560 19635
rect 10508 19592 10560 19601
rect 12164 19592 12216 19644
rect 12348 19592 12400 19644
rect 12624 19592 12676 19644
rect 7932 19456 7984 19508
rect 12716 19524 12768 19576
rect 16856 19592 16908 19644
rect 17684 19592 17736 19644
rect 10324 19456 10376 19508
rect 11980 19456 12032 19508
rect 17868 19524 17920 19576
rect 22744 19524 22796 19576
rect 8760 19388 8812 19440
rect 9956 19388 10008 19440
rect 11796 19388 11848 19440
rect 13176 19388 13228 19440
rect 14188 19431 14240 19440
rect 14188 19397 14197 19431
rect 14197 19397 14231 19431
rect 14231 19397 14240 19431
rect 14188 19388 14240 19397
rect 14556 19388 14608 19440
rect 17592 19388 17644 19440
rect 19248 19388 19300 19440
rect 6920 19227 6972 19236
rect 6920 19193 6929 19227
rect 6929 19193 6963 19227
rect 6963 19193 6972 19227
rect 6920 19184 6972 19193
rect 10324 19227 10376 19236
rect 10324 19193 10333 19227
rect 10333 19193 10367 19227
rect 10367 19193 10376 19227
rect 10324 19184 10376 19193
rect 12072 19116 12124 19168
rect 12992 19116 13044 19168
rect 14188 19116 14240 19168
rect 14832 19116 14884 19168
rect 17592 19184 17644 19236
rect 19248 19116 19300 19168
rect 22192 19184 22244 19236
rect 8944 19048 8996 19100
rect 9956 19091 10008 19100
rect 9956 19057 9965 19091
rect 9965 19057 9999 19091
rect 9999 19057 10008 19091
rect 9956 19048 10008 19057
rect 6920 18980 6972 19032
rect 10232 18980 10284 19032
rect 10968 18980 11020 19032
rect 11520 19048 11572 19100
rect 11980 19091 12032 19100
rect 11980 19057 11989 19091
rect 11989 19057 12023 19091
rect 12023 19057 12032 19091
rect 11980 19048 12032 19057
rect 14556 19091 14608 19100
rect 14556 19057 14565 19091
rect 14565 19057 14599 19091
rect 14599 19057 14608 19091
rect 14556 19048 14608 19057
rect 16120 19048 16172 19100
rect 20168 19048 20220 19100
rect 11612 19023 11664 19032
rect 11612 18989 11621 19023
rect 11621 18989 11655 19023
rect 11655 18989 11664 19023
rect 11612 18980 11664 18989
rect 11796 19023 11848 19032
rect 11796 18989 11805 19023
rect 11805 18989 11839 19023
rect 11839 18989 11848 19023
rect 11796 18980 11848 18989
rect 13360 18980 13412 19032
rect 17132 18980 17184 19032
rect 17316 18980 17368 19032
rect 17868 18980 17920 19032
rect 20352 18980 20404 19032
rect 22744 18980 22796 19032
rect 9956 18844 10008 18896
rect 10968 18844 11020 18896
rect 17776 18844 17828 18896
rect 18604 18887 18656 18896
rect 18604 18853 18613 18887
rect 18613 18853 18647 18887
rect 18647 18853 18656 18887
rect 18604 18844 18656 18853
rect 20904 18844 20956 18896
rect 21272 18844 21324 18896
rect 8760 18640 8812 18692
rect 12164 18640 12216 18692
rect 13176 18640 13228 18692
rect 20076 18640 20128 18692
rect 20904 18640 20956 18692
rect 22928 18640 22980 18692
rect 6736 18547 6788 18556
rect 6736 18513 6745 18547
rect 6745 18513 6779 18547
rect 6779 18513 6788 18547
rect 6736 18504 6788 18513
rect 14832 18572 14884 18624
rect 16120 18572 16172 18624
rect 17592 18572 17644 18624
rect 17776 18615 17828 18624
rect 17776 18581 17785 18615
rect 17785 18581 17819 18615
rect 17819 18581 17828 18615
rect 17776 18572 17828 18581
rect 20168 18572 20220 18624
rect 9128 18504 9180 18556
rect 10968 18547 11020 18556
rect 10968 18513 10996 18547
rect 10996 18513 11020 18547
rect 10968 18504 11020 18513
rect 13452 18504 13504 18556
rect 15568 18504 15620 18556
rect 17868 18547 17920 18556
rect 17868 18513 17877 18547
rect 17877 18513 17911 18547
rect 17911 18513 17920 18547
rect 17868 18504 17920 18513
rect 21640 18572 21692 18624
rect 22192 18504 22244 18556
rect 22928 18504 22980 18556
rect 8668 18436 8720 18488
rect 9036 18479 9088 18488
rect 9036 18445 9045 18479
rect 9045 18445 9079 18479
rect 9079 18445 9088 18479
rect 9036 18436 9088 18445
rect 10692 18479 10744 18488
rect 10692 18445 10701 18479
rect 10701 18445 10735 18479
rect 10735 18445 10744 18479
rect 10692 18436 10744 18445
rect 14556 18436 14608 18488
rect 17316 18479 17368 18488
rect 17316 18445 17325 18479
rect 17325 18445 17359 18479
rect 17359 18445 17368 18479
rect 17316 18436 17368 18445
rect 17684 18436 17736 18488
rect 12992 18368 13044 18420
rect 6552 18300 6604 18352
rect 8852 18300 8904 18352
rect 15752 18300 15804 18352
rect 18420 18300 18472 18352
rect 18880 18300 18932 18352
rect 19892 18436 19944 18488
rect 20352 18300 20404 18352
rect 21824 18300 21876 18352
rect 7472 18028 7524 18080
rect 8852 18096 8904 18148
rect 9036 18096 9088 18148
rect 11980 18028 12032 18080
rect 13268 18096 13320 18148
rect 26424 18096 26476 18148
rect 16488 18028 16540 18080
rect 17684 18071 17736 18080
rect 17684 18037 17693 18071
rect 17693 18037 17727 18071
rect 17727 18037 17736 18071
rect 17684 18028 17736 18037
rect 9956 18003 10008 18012
rect 9956 17969 9965 18003
rect 9965 17969 9999 18003
rect 9999 17969 10008 18003
rect 9956 17960 10008 17969
rect 6920 17892 6972 17944
rect 9588 17892 9640 17944
rect 9772 17892 9824 17944
rect 10232 17892 10284 17944
rect 11336 17960 11388 18012
rect 12072 17960 12124 18012
rect 12256 17960 12308 18012
rect 22744 18003 22796 18012
rect 22744 17969 22753 18003
rect 22753 17969 22787 18003
rect 22787 17969 22796 18003
rect 12164 17892 12216 17944
rect 14280 17867 14332 17876
rect 14280 17833 14308 17867
rect 14308 17833 14332 17867
rect 14280 17824 14332 17833
rect 15568 17892 15620 17944
rect 15752 17935 15804 17944
rect 15752 17901 15761 17935
rect 15761 17901 15795 17935
rect 15795 17901 15804 17935
rect 15752 17892 15804 17901
rect 15844 17935 15896 17944
rect 15844 17901 15853 17935
rect 15853 17901 15887 17935
rect 15887 17901 15896 17935
rect 15844 17892 15896 17901
rect 16028 17892 16080 17944
rect 22744 17960 22796 17969
rect 17316 17892 17368 17944
rect 19800 17935 19852 17944
rect 19800 17901 19809 17935
rect 19809 17901 19843 17935
rect 19843 17901 19852 17935
rect 19800 17892 19852 17901
rect 14464 17824 14516 17876
rect 16304 17824 16356 17876
rect 21456 17892 21508 17944
rect 22468 17935 22520 17944
rect 22468 17901 22492 17935
rect 22492 17901 22520 17935
rect 22468 17892 22520 17901
rect 7104 17756 7156 17808
rect 10324 17756 10376 17808
rect 10968 17756 11020 17808
rect 13360 17799 13412 17808
rect 13360 17765 13369 17799
rect 13369 17765 13403 17799
rect 13403 17765 13412 17799
rect 13360 17756 13412 17765
rect 14832 17756 14884 17808
rect 21456 17756 21508 17808
rect 9588 17552 9640 17604
rect 9772 17484 9824 17536
rect 7288 17416 7340 17468
rect 7472 17459 7524 17468
rect 7472 17425 7500 17459
rect 7500 17425 7524 17459
rect 7472 17416 7524 17425
rect 8852 17416 8904 17468
rect 6552 17391 6604 17400
rect 6552 17357 6561 17391
rect 6561 17357 6595 17391
rect 6595 17357 6604 17391
rect 6552 17348 6604 17357
rect 10140 17416 10192 17468
rect 12256 17552 12308 17604
rect 10692 17416 10744 17468
rect 14096 17484 14148 17536
rect 6828 17255 6880 17264
rect 6828 17221 6837 17255
rect 6837 17221 6871 17255
rect 6871 17221 6880 17255
rect 6828 17212 6880 17221
rect 10324 17348 10376 17400
rect 12992 17416 13044 17468
rect 14464 17416 14516 17468
rect 13360 17280 13412 17332
rect 9036 17212 9088 17264
rect 10324 17212 10376 17264
rect 14740 17212 14792 17264
rect 15660 17459 15712 17468
rect 15660 17425 15669 17459
rect 15669 17425 15703 17459
rect 15703 17425 15712 17459
rect 15660 17416 15712 17425
rect 17684 17416 17736 17468
rect 17132 17348 17184 17400
rect 19708 17527 19760 17536
rect 19708 17493 19717 17527
rect 19717 17493 19751 17527
rect 19751 17493 19760 17527
rect 19708 17484 19760 17493
rect 19524 17459 19576 17468
rect 19524 17425 19533 17459
rect 19533 17425 19567 17459
rect 19567 17425 19576 17459
rect 19524 17416 19576 17425
rect 21824 17552 21876 17604
rect 22192 17459 22244 17468
rect 22192 17425 22216 17459
rect 22216 17425 22244 17459
rect 22192 17416 22244 17425
rect 22744 17416 22796 17468
rect 15844 17212 15896 17264
rect 16856 17212 16908 17264
rect 19064 17280 19116 17332
rect 21088 17323 21140 17332
rect 21088 17289 21097 17323
rect 21097 17289 21131 17323
rect 21131 17289 21140 17323
rect 21088 17280 21140 17289
rect 17868 17212 17920 17264
rect 18604 17212 18656 17264
rect 20168 17212 20220 17264
rect 10140 17008 10192 17060
rect 11336 17051 11388 17060
rect 11336 17017 11345 17051
rect 11345 17017 11379 17051
rect 11379 17017 11388 17051
rect 11336 17008 11388 17017
rect 11980 17051 12032 17060
rect 11980 17017 11989 17051
rect 11989 17017 12023 17051
rect 12023 17017 12032 17051
rect 11980 17008 12032 17017
rect 15292 17008 15344 17060
rect 16304 17008 16356 17060
rect 19708 17008 19760 17060
rect 12072 16940 12124 16992
rect 10876 16915 10928 16924
rect 10876 16881 10885 16915
rect 10885 16881 10919 16915
rect 10919 16881 10928 16915
rect 10876 16872 10928 16881
rect 12900 16872 12952 16924
rect 10324 16804 10376 16856
rect 11612 16804 11664 16856
rect 11796 16847 11848 16856
rect 11796 16813 11805 16847
rect 11805 16813 11839 16847
rect 11839 16813 11848 16847
rect 11796 16804 11848 16813
rect 11888 16804 11940 16856
rect 13268 16804 13320 16856
rect 14280 16872 14332 16924
rect 18144 16915 18196 16924
rect 18144 16881 18153 16915
rect 18153 16881 18187 16915
rect 18187 16881 18196 16915
rect 18144 16872 18196 16881
rect 20076 16872 20128 16924
rect 23480 16872 23532 16924
rect 14096 16847 14148 16856
rect 14096 16813 14105 16847
rect 14105 16813 14139 16847
rect 14139 16813 14148 16847
rect 14096 16804 14148 16813
rect 14464 16804 14516 16856
rect 14648 16847 14700 16856
rect 14648 16813 14676 16847
rect 14676 16813 14700 16847
rect 14648 16804 14700 16813
rect 15568 16804 15620 16856
rect 18420 16804 18472 16856
rect 20904 16847 20956 16856
rect 20904 16813 20913 16847
rect 20913 16813 20947 16847
rect 20947 16813 20956 16847
rect 20904 16804 20956 16813
rect 16672 16736 16724 16788
rect 17776 16736 17828 16788
rect 20720 16779 20772 16788
rect 20720 16745 20729 16779
rect 20729 16745 20763 16779
rect 20763 16745 20772 16779
rect 20720 16736 20772 16745
rect 21456 16736 21508 16788
rect 13084 16668 13136 16720
rect 20076 16668 20128 16720
rect 20168 16668 20220 16720
rect 20996 16668 21048 16720
rect 8852 16464 8904 16516
rect 11612 16464 11664 16516
rect 13084 16464 13136 16516
rect 13268 16464 13320 16516
rect 15752 16464 15804 16516
rect 7932 16396 7984 16448
rect 6184 16371 6236 16380
rect 6184 16337 6193 16371
rect 6193 16337 6227 16371
rect 6227 16337 6236 16371
rect 6184 16328 6236 16337
rect 6920 16328 6972 16380
rect 7288 16328 7340 16380
rect 9036 16371 9088 16380
rect 9036 16337 9045 16371
rect 9045 16337 9079 16371
rect 9079 16337 9088 16371
rect 9036 16328 9088 16337
rect 10968 16396 11020 16448
rect 12808 16396 12860 16448
rect 14832 16396 14884 16448
rect 15384 16439 15436 16448
rect 15384 16405 15412 16439
rect 15412 16405 15436 16439
rect 15384 16396 15436 16405
rect 10600 16328 10652 16380
rect 11612 16328 11664 16380
rect 11980 16328 12032 16380
rect 13360 16328 13412 16380
rect 15936 16328 15988 16380
rect 16672 16464 16724 16516
rect 17776 16464 17828 16516
rect 20720 16464 20772 16516
rect 21640 16464 21692 16516
rect 22192 16464 22244 16516
rect 22376 16464 22428 16516
rect 18604 16396 18656 16448
rect 20352 16439 20404 16448
rect 20352 16405 20380 16439
rect 20380 16405 20404 16439
rect 20352 16396 20404 16405
rect 16672 16371 16724 16380
rect 16672 16337 16681 16371
rect 16681 16337 16715 16371
rect 16715 16337 16724 16371
rect 16672 16328 16724 16337
rect 19892 16328 19944 16380
rect 8852 16303 8904 16312
rect 8852 16269 8861 16303
rect 8861 16269 8895 16303
rect 8895 16269 8904 16303
rect 8852 16260 8904 16269
rect 9864 16260 9916 16312
rect 16856 16260 16908 16312
rect 17960 16260 18012 16312
rect 22284 16260 22336 16312
rect 22928 16260 22980 16312
rect 9220 16235 9272 16244
rect 9220 16201 9229 16235
rect 9229 16201 9263 16235
rect 9263 16201 9272 16235
rect 9220 16192 9272 16201
rect 10232 16192 10284 16244
rect 11888 16192 11940 16244
rect 9036 16124 9088 16176
rect 10048 16124 10100 16176
rect 10968 16124 11020 16176
rect 12716 16167 12768 16176
rect 12716 16133 12725 16167
rect 12725 16133 12759 16167
rect 12759 16133 12768 16167
rect 12716 16124 12768 16133
rect 21272 16124 21324 16176
rect 6920 15920 6972 15972
rect 8852 15920 8904 15972
rect 11152 15920 11204 15972
rect 11796 15963 11848 15972
rect 11796 15929 11805 15963
rect 11805 15929 11839 15963
rect 11839 15929 11848 15963
rect 11796 15920 11848 15929
rect 12992 15920 13044 15972
rect 9036 15895 9088 15904
rect 7196 15716 7248 15768
rect 7472 15716 7524 15768
rect 7932 15716 7984 15768
rect 9036 15861 9045 15895
rect 9045 15861 9079 15895
rect 9079 15861 9088 15895
rect 9036 15852 9088 15861
rect 8944 15716 8996 15768
rect 9496 15759 9548 15768
rect 9496 15725 9505 15759
rect 9505 15725 9539 15759
rect 9539 15725 9548 15759
rect 9496 15716 9548 15725
rect 10048 15716 10100 15768
rect 10784 15716 10836 15768
rect 10416 15648 10468 15700
rect 11612 15716 11664 15768
rect 12348 15716 12400 15768
rect 12440 15648 12492 15700
rect 16856 15852 16908 15904
rect 16672 15827 16724 15836
rect 16672 15793 16681 15827
rect 16681 15793 16715 15827
rect 16715 15793 16724 15827
rect 16672 15784 16724 15793
rect 14464 15716 14516 15768
rect 16948 15716 17000 15768
rect 8760 15623 8812 15632
rect 8760 15589 8769 15623
rect 8769 15589 8803 15623
rect 8803 15589 8812 15623
rect 8760 15580 8812 15589
rect 10232 15580 10284 15632
rect 14280 15580 14332 15632
rect 17316 15648 17368 15700
rect 18604 15716 18656 15768
rect 20076 15784 20128 15836
rect 22744 15827 22796 15836
rect 22744 15793 22753 15827
rect 22753 15793 22787 15827
rect 22787 15793 22796 15827
rect 22744 15784 22796 15793
rect 17776 15623 17828 15632
rect 17776 15589 17785 15623
rect 17785 15589 17819 15623
rect 17819 15589 17828 15623
rect 17776 15580 17828 15589
rect 19064 15759 19116 15768
rect 19064 15725 19073 15759
rect 19073 15725 19107 15759
rect 19107 15725 19116 15759
rect 19064 15716 19116 15725
rect 20996 15716 21048 15768
rect 21456 15716 21508 15768
rect 21916 15648 21968 15700
rect 19064 15580 19116 15632
rect 21732 15580 21784 15632
rect 6184 15376 6236 15428
rect 9220 15376 9272 15428
rect 12072 15308 12124 15360
rect 6828 15240 6880 15292
rect 7932 15240 7984 15292
rect 8668 15240 8720 15292
rect 8944 15240 8996 15292
rect 10232 15240 10284 15292
rect 10784 15240 10836 15292
rect 11888 15240 11940 15292
rect 12624 15240 12676 15292
rect 16948 15376 17000 15428
rect 18972 15376 19024 15428
rect 21088 15308 21140 15360
rect 14740 15240 14792 15292
rect 15660 15240 15712 15292
rect 10416 15215 10468 15224
rect 10416 15181 10425 15215
rect 10425 15181 10459 15215
rect 10459 15181 10468 15215
rect 10692 15215 10744 15224
rect 10416 15172 10468 15181
rect 10692 15181 10701 15215
rect 10701 15181 10735 15215
rect 10735 15181 10744 15215
rect 10692 15172 10744 15181
rect 11796 15172 11848 15224
rect 13176 15215 13228 15224
rect 13176 15181 13185 15215
rect 13185 15181 13219 15215
rect 13219 15181 13228 15215
rect 13176 15172 13228 15181
rect 16028 15172 16080 15224
rect 16856 15240 16908 15292
rect 18604 15240 18656 15292
rect 17960 15172 18012 15224
rect 21456 15215 21508 15224
rect 21456 15181 21465 15215
rect 21465 15181 21499 15215
rect 21499 15181 21508 15215
rect 21456 15172 21508 15181
rect 22284 15215 22336 15224
rect 22284 15181 22293 15215
rect 22293 15181 22327 15215
rect 22327 15181 22336 15215
rect 22284 15172 22336 15181
rect 11336 15036 11388 15088
rect 12808 15036 12860 15088
rect 14464 15147 14516 15156
rect 14464 15113 14473 15147
rect 14473 15113 14507 15147
rect 14507 15113 14516 15147
rect 14464 15104 14516 15113
rect 19800 15104 19852 15156
rect 15936 15036 15988 15088
rect 16304 15036 16356 15088
rect 17316 15036 17368 15088
rect 19984 15036 20036 15088
rect 22468 15079 22520 15088
rect 22468 15045 22477 15079
rect 22477 15045 22511 15079
rect 22511 15045 22520 15079
rect 22468 15036 22520 15045
rect 10140 14832 10192 14884
rect 10416 14832 10468 14884
rect 10692 14832 10744 14884
rect 9036 14764 9088 14816
rect 17408 14832 17460 14884
rect 20996 14832 21048 14884
rect 20352 14764 20404 14816
rect 6920 14739 6972 14748
rect 6920 14705 6929 14739
rect 6929 14705 6963 14739
rect 6963 14705 6972 14739
rect 6920 14696 6972 14705
rect 6736 14628 6788 14680
rect 18236 14696 18288 14748
rect 18788 14739 18840 14748
rect 18788 14705 18797 14739
rect 18797 14705 18831 14739
rect 18831 14705 18840 14739
rect 18788 14696 18840 14705
rect 20444 14696 20496 14748
rect 22744 14739 22796 14748
rect 10876 14671 10928 14680
rect 10876 14637 10885 14671
rect 10885 14637 10919 14671
rect 10919 14637 10928 14671
rect 10876 14628 10928 14637
rect 10968 14628 11020 14680
rect 12348 14628 12400 14680
rect 13360 14628 13412 14680
rect 14464 14671 14516 14680
rect 14464 14637 14473 14671
rect 14473 14637 14507 14671
rect 14507 14637 14516 14671
rect 14464 14628 14516 14637
rect 16212 14671 16264 14680
rect 16212 14637 16221 14671
rect 16221 14637 16255 14671
rect 16255 14637 16264 14671
rect 16212 14628 16264 14637
rect 16488 14671 16540 14680
rect 16488 14637 16516 14671
rect 16516 14637 16540 14671
rect 16488 14628 16540 14637
rect 6552 14492 6604 14544
rect 15200 14560 15252 14612
rect 18512 14671 18564 14680
rect 18512 14637 18521 14671
rect 18521 14637 18555 14671
rect 18555 14637 18564 14671
rect 18512 14628 18564 14637
rect 20076 14628 20128 14680
rect 20352 14628 20404 14680
rect 22744 14705 22753 14739
rect 22753 14705 22787 14739
rect 22787 14705 22796 14739
rect 22744 14696 22796 14705
rect 22468 14671 22520 14680
rect 22468 14637 22492 14671
rect 22492 14637 22520 14671
rect 22468 14628 22520 14637
rect 13452 14492 13504 14544
rect 14556 14492 14608 14544
rect 15844 14535 15896 14544
rect 15844 14501 15853 14535
rect 15853 14501 15887 14535
rect 15887 14501 15896 14535
rect 15844 14492 15896 14501
rect 18604 14560 18656 14612
rect 18972 14560 19024 14612
rect 19984 14560 20036 14612
rect 20168 14535 20220 14544
rect 20168 14501 20177 14535
rect 20177 14501 20211 14535
rect 20211 14501 20220 14535
rect 20168 14492 20220 14501
rect 20628 14492 20680 14544
rect 10600 14288 10652 14340
rect 11796 14288 11848 14340
rect 14556 14288 14608 14340
rect 17132 14288 17184 14340
rect 18972 14331 19024 14340
rect 18972 14297 18981 14331
rect 18981 14297 19015 14331
rect 19015 14297 19024 14331
rect 18972 14288 19024 14297
rect 21916 14288 21968 14340
rect 13452 14220 13504 14272
rect 14280 14220 14332 14272
rect 6552 14195 6604 14204
rect 6552 14161 6561 14195
rect 6561 14161 6595 14195
rect 6595 14161 6604 14195
rect 6552 14152 6604 14161
rect 7288 14152 7340 14204
rect 7932 14152 7984 14204
rect 11152 14152 11204 14204
rect 12808 14152 12860 14204
rect 14372 14195 14424 14204
rect 6920 14084 6972 14136
rect 12348 14084 12400 14136
rect 14372 14161 14381 14195
rect 14381 14161 14415 14195
rect 14415 14161 14424 14195
rect 14372 14152 14424 14161
rect 14556 14195 14608 14204
rect 14556 14161 14565 14195
rect 14565 14161 14599 14195
rect 14599 14161 14608 14195
rect 14556 14152 14608 14161
rect 15200 14152 15252 14204
rect 15752 14152 15804 14204
rect 16948 14152 17000 14204
rect 18604 14195 18656 14204
rect 18604 14161 18628 14195
rect 18628 14161 18656 14195
rect 18604 14152 18656 14161
rect 18788 14152 18840 14204
rect 19064 14152 19116 14204
rect 15568 14084 15620 14136
rect 16580 14127 16632 14136
rect 16580 14093 16589 14127
rect 16589 14093 16623 14127
rect 16623 14093 16632 14127
rect 16580 14084 16632 14093
rect 15476 14059 15528 14068
rect 15476 14025 15485 14059
rect 15485 14025 15519 14059
rect 15519 14025 15528 14059
rect 15476 14016 15528 14025
rect 9128 13948 9180 14000
rect 11796 13948 11848 14000
rect 20352 14152 20404 14204
rect 21272 14195 21324 14204
rect 21272 14161 21296 14195
rect 21296 14161 21324 14195
rect 21272 14152 21324 14161
rect 21456 14152 21508 14204
rect 22284 14152 22336 14204
rect 19892 14084 19944 14136
rect 22928 13948 22980 14000
rect 6736 13744 6788 13796
rect 7932 13744 7984 13796
rect 9036 13744 9088 13796
rect 11336 13744 11388 13796
rect 14372 13744 14424 13796
rect 10232 13676 10284 13728
rect 10784 13676 10836 13728
rect 6368 13608 6420 13660
rect 9128 13608 9180 13660
rect 12532 13608 12584 13660
rect 12716 13608 12768 13660
rect 18328 13787 18380 13796
rect 18328 13753 18337 13787
rect 18337 13753 18371 13787
rect 18371 13753 18380 13787
rect 18328 13744 18380 13753
rect 21732 13744 21784 13796
rect 17960 13608 18012 13660
rect 18788 13651 18840 13660
rect 18788 13617 18797 13651
rect 18797 13617 18831 13651
rect 18831 13617 18840 13651
rect 18788 13608 18840 13617
rect 6184 13404 6236 13456
rect 6736 13472 6788 13524
rect 6920 13540 6972 13592
rect 9496 13540 9548 13592
rect 10968 13540 11020 13592
rect 10692 13447 10744 13456
rect 10692 13413 10701 13447
rect 10701 13413 10735 13447
rect 10735 13413 10744 13447
rect 10692 13404 10744 13413
rect 11612 13404 11664 13456
rect 13360 13540 13412 13592
rect 17776 13540 17828 13592
rect 17132 13472 17184 13524
rect 19892 13608 19944 13660
rect 22744 13651 22796 13660
rect 22744 13617 22753 13651
rect 22753 13617 22787 13651
rect 22787 13617 22796 13651
rect 22744 13608 22796 13617
rect 20444 13583 20496 13592
rect 20444 13549 20453 13583
rect 20453 13549 20487 13583
rect 20487 13549 20496 13583
rect 20444 13540 20496 13549
rect 20720 13540 20772 13592
rect 22468 13583 22520 13592
rect 22468 13549 22492 13583
rect 22492 13549 22520 13583
rect 22468 13540 22520 13549
rect 20536 13515 20588 13524
rect 20536 13481 20545 13515
rect 20545 13481 20579 13515
rect 20579 13481 20588 13515
rect 20536 13472 20588 13481
rect 12992 13404 13044 13456
rect 13452 13404 13504 13456
rect 20168 13404 20220 13456
rect 6920 13200 6972 13252
rect 9496 13200 9548 13252
rect 6368 13064 6420 13116
rect 6736 13107 6788 13116
rect 6736 13073 6745 13107
rect 6745 13073 6779 13107
rect 6779 13073 6788 13107
rect 6736 13064 6788 13073
rect 10784 13132 10836 13184
rect 7288 13039 7340 13048
rect 7288 13005 7297 13039
rect 7297 13005 7331 13039
rect 7331 13005 7340 13039
rect 7288 12996 7340 13005
rect 12532 13200 12584 13252
rect 16028 13200 16080 13252
rect 17316 13200 17368 13252
rect 12716 13132 12768 13184
rect 13452 13132 13504 13184
rect 14556 13132 14608 13184
rect 16120 13132 16172 13184
rect 20536 13200 20588 13252
rect 21732 13200 21784 13252
rect 21640 13132 21692 13184
rect 13360 13064 13412 13116
rect 15292 13107 15344 13116
rect 10692 12996 10744 13048
rect 11980 12996 12032 13048
rect 12348 12996 12400 13048
rect 15292 13073 15301 13107
rect 15301 13073 15335 13107
rect 15335 13073 15344 13107
rect 15292 13064 15344 13073
rect 15568 13064 15620 13116
rect 17224 13064 17276 13116
rect 17500 13064 17552 13116
rect 18788 13064 18840 13116
rect 20444 13064 20496 13116
rect 21824 13107 21876 13116
rect 21824 13073 21833 13107
rect 21833 13073 21867 13107
rect 21867 13073 21876 13107
rect 21824 13064 21876 13073
rect 22008 13064 22060 13116
rect 21456 13039 21508 13048
rect 10048 12928 10100 12980
rect 10784 12928 10836 12980
rect 21456 13005 21465 13039
rect 21465 13005 21499 13039
rect 21499 13005 21508 13039
rect 21456 12996 21508 13005
rect 15660 12860 15712 12912
rect 17040 12860 17092 12912
rect 17500 12903 17552 12912
rect 17500 12869 17509 12903
rect 17509 12869 17543 12903
rect 17543 12869 17552 12903
rect 17500 12860 17552 12869
rect 20168 12860 20220 12912
rect 10232 12656 10284 12708
rect 11980 12656 12032 12708
rect 10416 12588 10468 12640
rect 6552 12495 6604 12504
rect 6552 12461 6561 12495
rect 6561 12461 6595 12495
rect 6595 12461 6604 12495
rect 6552 12452 6604 12461
rect 7932 12520 7984 12572
rect 13268 12563 13320 12572
rect 13268 12529 13277 12563
rect 13277 12529 13311 12563
rect 13311 12529 13320 12563
rect 13268 12520 13320 12529
rect 16764 12656 16816 12708
rect 17132 12699 17184 12708
rect 8852 12452 8904 12504
rect 12992 12495 13044 12504
rect 12992 12461 13016 12495
rect 13016 12461 13044 12495
rect 12992 12452 13044 12461
rect 13452 12452 13504 12504
rect 15844 12520 15896 12572
rect 15568 12452 15620 12504
rect 16764 12495 16816 12504
rect 16764 12461 16773 12495
rect 16773 12461 16807 12495
rect 16807 12461 16816 12495
rect 16764 12452 16816 12461
rect 17132 12665 17141 12699
rect 17141 12665 17175 12699
rect 17175 12665 17184 12699
rect 17132 12656 17184 12665
rect 21640 12656 21692 12708
rect 22928 12656 22980 12708
rect 18788 12520 18840 12572
rect 17132 12452 17184 12504
rect 20168 12495 20220 12504
rect 6736 12384 6788 12436
rect 6368 12316 6420 12368
rect 10232 12316 10284 12368
rect 18972 12384 19024 12436
rect 16764 12316 16816 12368
rect 17960 12316 18012 12368
rect 20168 12461 20177 12495
rect 20177 12461 20211 12495
rect 20211 12461 20220 12495
rect 20168 12452 20220 12461
rect 21088 12495 21140 12504
rect 21088 12461 21097 12495
rect 21097 12461 21131 12495
rect 21131 12461 21140 12495
rect 21088 12452 21140 12461
rect 21640 12427 21692 12436
rect 21640 12393 21668 12427
rect 21668 12393 21692 12427
rect 21640 12384 21692 12393
rect 28724 12316 28776 12368
rect 6736 12112 6788 12164
rect 8852 12155 8904 12164
rect 8852 12121 8861 12155
rect 8861 12121 8895 12155
rect 8895 12121 8904 12155
rect 8852 12112 8904 12121
rect 6552 11976 6604 12028
rect 10784 12044 10836 12096
rect 7288 11908 7340 11960
rect 14556 12112 14608 12164
rect 16764 12112 16816 12164
rect 10048 11951 10100 11960
rect 10048 11917 10057 11951
rect 10057 11917 10091 11951
rect 10091 11917 10100 11951
rect 10048 11908 10100 11917
rect 10232 11951 10284 11960
rect 10232 11917 10241 11951
rect 10241 11917 10275 11951
rect 10275 11917 10284 11951
rect 10232 11908 10284 11917
rect 13268 12044 13320 12096
rect 15660 12044 15712 12096
rect 21640 12112 21692 12164
rect 17500 12044 17552 12096
rect 17960 12087 18012 12096
rect 17960 12053 17969 12087
rect 17969 12053 18003 12087
rect 18003 12053 18012 12087
rect 17960 12044 18012 12053
rect 20076 12044 20128 12096
rect 13452 11976 13504 12028
rect 15476 11976 15528 12028
rect 15568 11976 15620 12028
rect 11980 11908 12032 11960
rect 10600 11840 10652 11892
rect 6368 11815 6420 11824
rect 6368 11781 6377 11815
rect 6377 11781 6411 11815
rect 6411 11781 6420 11815
rect 6368 11772 6420 11781
rect 17132 12019 17184 12028
rect 17132 11985 17141 12019
rect 17141 11985 17175 12019
rect 17175 11985 17184 12019
rect 17132 11976 17184 11985
rect 21180 12019 21232 12028
rect 17316 11883 17368 11892
rect 17316 11849 17325 11883
rect 17325 11849 17359 11883
rect 17359 11849 17368 11883
rect 17316 11840 17368 11849
rect 21180 11985 21204 12019
rect 21204 11985 21232 12019
rect 21180 11976 21232 11985
rect 18512 11951 18564 11960
rect 18512 11917 18521 11951
rect 18521 11917 18555 11951
rect 18555 11917 18564 11951
rect 18512 11908 18564 11917
rect 21456 11951 21508 11960
rect 21456 11917 21465 11951
rect 21465 11917 21499 11951
rect 21499 11917 21508 11951
rect 21456 11908 21508 11917
rect 22192 11908 22244 11960
rect 18236 11840 18288 11892
rect 17592 11815 17644 11824
rect 17592 11781 17601 11815
rect 17601 11781 17635 11815
rect 17635 11781 17644 11815
rect 17592 11772 17644 11781
rect 19984 11772 20036 11824
rect 21732 11772 21784 11824
rect 7932 11568 7984 11620
rect 10416 11568 10468 11620
rect 13268 11568 13320 11620
rect 6368 11500 6420 11552
rect 8852 11500 8904 11552
rect 11980 11500 12032 11552
rect 21640 11500 21692 11552
rect 14004 11475 14056 11484
rect 6184 11364 6236 11416
rect 6644 11407 6696 11416
rect 6644 11373 6653 11407
rect 6653 11373 6687 11407
rect 6687 11373 6696 11407
rect 6644 11364 6696 11373
rect 7196 11364 7248 11416
rect 8668 11364 8720 11416
rect 14004 11441 14013 11475
rect 14013 11441 14047 11475
rect 14047 11441 14056 11475
rect 14004 11432 14056 11441
rect 22744 11475 22796 11484
rect 22744 11441 22753 11475
rect 22753 11441 22787 11475
rect 22787 11441 22796 11475
rect 22744 11432 22796 11441
rect 10508 11364 10560 11416
rect 11612 11407 11664 11416
rect 11612 11373 11621 11407
rect 11621 11373 11655 11407
rect 11655 11373 11664 11407
rect 11612 11364 11664 11373
rect 12348 11364 12400 11416
rect 14556 11364 14608 11416
rect 15476 11407 15528 11416
rect 15476 11373 15485 11407
rect 15485 11373 15519 11407
rect 15519 11373 15528 11407
rect 15476 11364 15528 11373
rect 15844 11407 15896 11416
rect 15844 11373 15853 11407
rect 15853 11373 15887 11407
rect 15887 11373 15896 11407
rect 15844 11364 15896 11373
rect 16856 11407 16908 11416
rect 16856 11373 16865 11407
rect 16865 11373 16899 11407
rect 16899 11373 16908 11407
rect 16856 11364 16908 11373
rect 17592 11364 17644 11416
rect 18788 11407 18840 11416
rect 9036 11228 9088 11280
rect 15752 11339 15804 11348
rect 15752 11305 15761 11339
rect 15761 11305 15795 11339
rect 15795 11305 15804 11339
rect 18788 11373 18797 11407
rect 18797 11373 18831 11407
rect 18831 11373 18840 11407
rect 18788 11364 18840 11373
rect 21180 11364 21232 11416
rect 15752 11296 15804 11305
rect 19156 11296 19208 11348
rect 20444 11296 20496 11348
rect 20536 11296 20588 11348
rect 20812 11339 20864 11348
rect 20812 11305 20821 11339
rect 20821 11305 20855 11339
rect 20855 11305 20864 11339
rect 20812 11296 20864 11305
rect 17316 11228 17368 11280
rect 17868 11228 17920 11280
rect 18052 11228 18104 11280
rect 21364 11271 21416 11280
rect 21364 11237 21373 11271
rect 21373 11237 21407 11271
rect 21407 11237 21416 11271
rect 21364 11228 21416 11237
rect 11336 11024 11388 11076
rect 10600 10956 10652 11008
rect 6644 10888 6696 10940
rect 10048 10888 10100 10940
rect 10508 10888 10560 10940
rect 15752 11024 15804 11076
rect 20812 11024 20864 11076
rect 13452 10888 13504 10940
rect 15936 10888 15988 10940
rect 18420 10888 18472 10940
rect 21088 10956 21140 11008
rect 21364 10956 21416 11008
rect 20168 10888 20220 10940
rect 7288 10863 7340 10872
rect 7288 10829 7297 10863
rect 7297 10829 7331 10863
rect 7331 10829 7340 10863
rect 7288 10820 7340 10829
rect 9036 10820 9088 10872
rect 13268 10820 13320 10872
rect 16856 10820 16908 10872
rect 21456 10863 21508 10872
rect 21456 10829 21465 10863
rect 21465 10829 21499 10863
rect 21499 10829 21508 10863
rect 21456 10820 21508 10829
rect 21916 10820 21968 10872
rect 10876 10752 10928 10804
rect 8668 10727 8720 10736
rect 8668 10693 8677 10727
rect 8677 10693 8711 10727
rect 8711 10693 8720 10727
rect 8668 10684 8720 10693
rect 9036 10684 9088 10736
rect 14464 10684 14516 10736
rect 20536 10684 20588 10736
rect 26240 10684 26292 10736
rect 10508 10480 10560 10532
rect 13268 10480 13320 10532
rect 14556 10480 14608 10532
rect 16120 10480 16172 10532
rect 18236 10480 18288 10532
rect 8668 10412 8720 10464
rect 11336 10455 11388 10464
rect 11336 10421 11345 10455
rect 11345 10421 11379 10455
rect 11379 10421 11388 10455
rect 11336 10412 11388 10421
rect 17684 10455 17736 10464
rect 17684 10421 17693 10455
rect 17693 10421 17727 10455
rect 17727 10421 17736 10455
rect 17684 10412 17736 10421
rect 20260 10523 20312 10532
rect 20260 10489 20269 10523
rect 20269 10489 20303 10523
rect 20303 10489 20312 10523
rect 20260 10480 20312 10489
rect 6828 10319 6880 10328
rect 6828 10285 6837 10319
rect 6837 10285 6871 10319
rect 6871 10285 6880 10319
rect 6828 10276 6880 10285
rect 11612 10344 11664 10396
rect 17960 10344 18012 10396
rect 18788 10387 18840 10396
rect 18788 10353 18797 10387
rect 18797 10353 18831 10387
rect 18831 10353 18840 10387
rect 18788 10344 18840 10353
rect 21272 10344 21324 10396
rect 9128 10276 9180 10328
rect 12348 10276 12400 10328
rect 13268 10276 13320 10328
rect 14188 10319 14240 10328
rect 14188 10285 14197 10319
rect 14197 10285 14231 10319
rect 14231 10285 14240 10319
rect 14188 10276 14240 10285
rect 14464 10276 14516 10328
rect 15292 10276 15344 10328
rect 16856 10276 16908 10328
rect 18052 10319 18104 10328
rect 18052 10285 18061 10319
rect 18061 10285 18095 10319
rect 18095 10285 18104 10319
rect 18052 10276 18104 10285
rect 20352 10276 20404 10328
rect 20628 10319 20680 10328
rect 20628 10285 20637 10319
rect 20637 10285 20671 10319
rect 20671 10285 20680 10319
rect 20628 10276 20680 10285
rect 21456 10276 21508 10328
rect 9036 10208 9088 10260
rect 16120 10208 16172 10260
rect 17316 10251 17368 10260
rect 17316 10217 17340 10251
rect 17340 10217 17368 10251
rect 17316 10208 17368 10217
rect 14556 10140 14608 10192
rect 14924 10140 14976 10192
rect 17224 10140 17276 10192
rect 18144 10140 18196 10192
rect 23204 10276 23256 10328
rect 21916 10208 21968 10260
rect 20812 10140 20864 10192
rect 22744 10183 22796 10192
rect 22744 10149 22753 10183
rect 22753 10149 22787 10183
rect 22787 10149 22796 10183
rect 22744 10140 22796 10149
rect 6460 9936 6512 9988
rect 8852 9936 8904 9988
rect 17500 9936 17552 9988
rect 18052 9979 18104 9988
rect 18052 9945 18061 9979
rect 18061 9945 18095 9979
rect 18095 9945 18104 9979
rect 18052 9936 18104 9945
rect 14924 9868 14976 9920
rect 16396 9868 16448 9920
rect 10692 9800 10744 9852
rect 12624 9843 12676 9852
rect 12624 9809 12652 9843
rect 12652 9809 12676 9843
rect 12624 9800 12676 9809
rect 15292 9843 15344 9852
rect 15292 9809 15301 9843
rect 15301 9809 15335 9843
rect 15335 9809 15344 9843
rect 15292 9800 15344 9809
rect 15568 9843 15620 9852
rect 15568 9809 15577 9843
rect 15577 9809 15611 9843
rect 15611 9809 15620 9843
rect 15568 9800 15620 9809
rect 8300 9732 8352 9784
rect 10048 9732 10100 9784
rect 11336 9732 11388 9784
rect 12348 9775 12400 9784
rect 12348 9741 12357 9775
rect 12357 9741 12391 9775
rect 12391 9741 12400 9775
rect 12348 9732 12400 9741
rect 14280 9732 14332 9784
rect 16028 9800 16080 9852
rect 16764 9800 16816 9852
rect 18236 9936 18288 9988
rect 20628 9936 20680 9988
rect 22468 9979 22520 9988
rect 22468 9945 22477 9979
rect 22477 9945 22511 9979
rect 22511 9945 22520 9979
rect 22468 9936 22520 9945
rect 18328 9800 18380 9852
rect 19340 9800 19392 9852
rect 20168 9800 20220 9852
rect 20812 9800 20864 9852
rect 22192 9800 22244 9852
rect 15752 9732 15804 9784
rect 8208 9707 8260 9716
rect 8208 9673 8228 9707
rect 8228 9673 8260 9707
rect 8208 9664 8260 9673
rect 10876 9664 10928 9716
rect 11060 9664 11112 9716
rect 15936 9664 15988 9716
rect 19156 9707 19208 9716
rect 10324 9639 10376 9648
rect 10324 9605 10333 9639
rect 10333 9605 10367 9639
rect 10367 9605 10376 9639
rect 10324 9596 10376 9605
rect 12992 9596 13044 9648
rect 14280 9596 14332 9648
rect 17040 9596 17092 9648
rect 17408 9596 17460 9648
rect 19156 9673 19165 9707
rect 19165 9673 19199 9707
rect 19199 9673 19208 9707
rect 19156 9664 19208 9673
rect 21640 9707 21692 9716
rect 21640 9673 21649 9707
rect 21649 9673 21683 9707
rect 21683 9673 21692 9707
rect 21640 9664 21692 9673
rect 22192 9664 22244 9716
rect 8300 9435 8352 9444
rect 8300 9401 8309 9435
rect 8309 9401 8343 9435
rect 8343 9401 8352 9435
rect 8300 9392 8352 9401
rect 10692 9435 10744 9444
rect 10692 9401 10701 9435
rect 10701 9401 10735 9435
rect 10735 9401 10744 9435
rect 10692 9392 10744 9401
rect 11336 9392 11388 9444
rect 11612 9392 11664 9444
rect 10324 9324 10376 9376
rect 12992 9367 13044 9376
rect 12992 9333 13001 9367
rect 13001 9333 13035 9367
rect 13035 9333 13044 9367
rect 12992 9324 13044 9333
rect 6644 9299 6696 9308
rect 6644 9265 6653 9299
rect 6653 9265 6687 9299
rect 6687 9265 6696 9299
rect 6644 9256 6696 9265
rect 9128 9256 9180 9308
rect 7196 9188 7248 9240
rect 14556 9392 14608 9444
rect 16120 9392 16172 9444
rect 20168 9392 20220 9444
rect 21640 9392 21692 9444
rect 19984 9324 20036 9376
rect 13084 9256 13136 9308
rect 13452 9256 13504 9308
rect 12440 9120 12492 9172
rect 15844 9188 15896 9240
rect 16764 9231 16816 9240
rect 16764 9197 16773 9231
rect 16773 9197 16807 9231
rect 16807 9197 16816 9231
rect 16764 9188 16816 9197
rect 17684 9188 17736 9240
rect 18696 9188 18748 9240
rect 20352 9188 20404 9240
rect 23388 9392 23440 9444
rect 16488 9163 16540 9172
rect 16488 9129 16497 9163
rect 16497 9129 16531 9163
rect 16531 9129 16540 9163
rect 16488 9120 16540 9129
rect 18512 9120 18564 9172
rect 19800 9120 19852 9172
rect 19984 9120 20036 9172
rect 19340 9052 19392 9104
rect 22100 9256 22152 9308
rect 22008 9120 22060 9172
rect 21180 9052 21232 9104
rect 21824 9052 21876 9104
rect 8852 8848 8904 8900
rect 6460 8712 6512 8764
rect 11060 8848 11112 8900
rect 12624 8848 12676 8900
rect 13268 8848 13320 8900
rect 15384 8848 15436 8900
rect 16488 8848 16540 8900
rect 7840 8712 7892 8764
rect 10692 8712 10744 8764
rect 14280 8780 14332 8832
rect 16948 8780 17000 8832
rect 20168 8848 20220 8900
rect 13268 8755 13320 8764
rect 13268 8721 13277 8755
rect 13277 8721 13311 8755
rect 13311 8721 13320 8755
rect 13268 8712 13320 8721
rect 13452 8712 13504 8764
rect 15476 8755 15528 8764
rect 15476 8721 15485 8755
rect 15485 8721 15519 8755
rect 15519 8721 15528 8755
rect 15476 8712 15528 8721
rect 16212 8712 16264 8764
rect 18328 8712 18380 8764
rect 13084 8644 13136 8696
rect 10416 8576 10468 8628
rect 8300 8508 8352 8560
rect 8668 8508 8720 8560
rect 16672 8576 16724 8628
rect 18512 8619 18564 8628
rect 18512 8585 18521 8619
rect 18521 8585 18555 8619
rect 18555 8585 18564 8619
rect 18512 8576 18564 8585
rect 17592 8508 17644 8560
rect 20260 8644 20312 8696
rect 20168 8576 20220 8628
rect 8300 8347 8352 8356
rect 8300 8313 8309 8347
rect 8309 8313 8343 8347
rect 8343 8313 8352 8347
rect 8300 8304 8352 8313
rect 10692 8347 10744 8356
rect 10692 8313 10701 8347
rect 10701 8313 10735 8347
rect 10735 8313 10744 8347
rect 10692 8304 10744 8313
rect 13268 8304 13320 8356
rect 17224 8347 17276 8356
rect 10692 8168 10744 8220
rect 16764 8236 16816 8288
rect 17224 8313 17233 8347
rect 17233 8313 17267 8347
rect 17267 8313 17276 8347
rect 17224 8304 17276 8313
rect 18236 8304 18288 8356
rect 17592 8236 17644 8288
rect 18972 8304 19024 8356
rect 21180 8304 21232 8356
rect 23204 8304 23256 8356
rect 6644 8100 6696 8152
rect 7196 8100 7248 8152
rect 9128 8100 9180 8152
rect 11796 8100 11848 8152
rect 14280 8143 14332 8152
rect 14280 8109 14289 8143
rect 14289 8109 14323 8143
rect 14323 8109 14332 8143
rect 14280 8100 14332 8109
rect 15016 8100 15068 8152
rect 18052 8100 18104 8152
rect 18512 8100 18564 8152
rect 19064 8143 19116 8152
rect 19064 8109 19092 8143
rect 19092 8109 19116 8143
rect 19064 8100 19116 8109
rect 20352 8100 20404 8152
rect 20536 8143 20588 8152
rect 20536 8109 20545 8143
rect 20545 8109 20579 8143
rect 20579 8109 20588 8143
rect 20536 8100 20588 8109
rect 21456 8100 21508 8152
rect 9404 8032 9456 8084
rect 11336 8075 11388 8084
rect 11336 8041 11364 8075
rect 11364 8041 11388 8075
rect 11336 8032 11388 8041
rect 14832 8032 14884 8084
rect 15200 8032 15252 8084
rect 19984 8032 20036 8084
rect 11980 7964 12032 8016
rect 13452 8007 13504 8016
rect 13452 7973 13461 8007
rect 13461 7973 13495 8007
rect 13495 7973 13504 8007
rect 13452 7964 13504 7973
rect 14464 7964 14516 8016
rect 20720 8032 20772 8084
rect 21640 8075 21692 8084
rect 21640 8041 21668 8075
rect 21668 8041 21692 8075
rect 21640 8032 21692 8041
rect 9404 7760 9456 7812
rect 10048 7760 10100 7812
rect 6644 7667 6696 7676
rect 6644 7633 6653 7667
rect 6653 7633 6687 7667
rect 6687 7633 6696 7667
rect 6644 7624 6696 7633
rect 7288 7624 7340 7676
rect 11336 7760 11388 7812
rect 10876 7667 10928 7676
rect 13268 7692 13320 7744
rect 15200 7760 15252 7812
rect 16028 7803 16080 7812
rect 16028 7769 16037 7803
rect 16037 7769 16071 7803
rect 16071 7769 16080 7803
rect 16028 7760 16080 7769
rect 18972 7760 19024 7812
rect 10876 7633 10900 7667
rect 10900 7633 10928 7667
rect 10876 7624 10928 7633
rect 12900 7624 12952 7676
rect 8852 7599 8904 7608
rect 8852 7565 8861 7599
rect 8861 7565 8895 7599
rect 8895 7565 8904 7599
rect 8852 7556 8904 7565
rect 5908 7488 5960 7540
rect 6368 7488 6420 7540
rect 10048 7556 10100 7608
rect 12348 7599 12400 7608
rect 12348 7565 12357 7599
rect 12357 7565 12391 7599
rect 12391 7565 12400 7599
rect 12348 7556 12400 7565
rect 20168 7692 20220 7744
rect 14004 7624 14056 7676
rect 14464 7624 14516 7676
rect 14740 7624 14792 7676
rect 18328 7624 18380 7676
rect 18604 7624 18656 7676
rect 19984 7624 20036 7676
rect 22376 7624 22428 7676
rect 17132 7599 17184 7608
rect 17132 7565 17141 7599
rect 17141 7565 17175 7599
rect 17175 7565 17184 7599
rect 17132 7556 17184 7565
rect 17408 7556 17460 7608
rect 18052 7556 18104 7608
rect 20260 7556 20312 7608
rect 21548 7556 21600 7608
rect 11612 7531 11664 7540
rect 11612 7497 11621 7531
rect 11621 7497 11655 7531
rect 11655 7497 11664 7531
rect 11612 7488 11664 7497
rect 16580 7488 16632 7540
rect 6092 7463 6144 7472
rect 6092 7429 6101 7463
rect 6101 7429 6135 7463
rect 6135 7429 6144 7463
rect 6092 7420 6144 7429
rect 9128 7420 9180 7472
rect 12532 7420 12584 7472
rect 13084 7420 13136 7472
rect 18144 7420 18196 7472
rect 19800 7488 19852 7540
rect 22008 7488 22060 7540
rect 6092 7216 6144 7268
rect 6368 7259 6420 7268
rect 6368 7225 6377 7259
rect 6377 7225 6411 7259
rect 6411 7225 6420 7259
rect 6368 7216 6420 7225
rect 13176 7216 13228 7268
rect 12164 7191 12216 7200
rect 12164 7157 12196 7191
rect 12196 7157 12216 7191
rect 12164 7148 12216 7157
rect 6920 7123 6972 7132
rect 6920 7089 6929 7123
rect 6929 7089 6963 7123
rect 6963 7089 6972 7123
rect 6920 7080 6972 7089
rect 12532 7123 12584 7132
rect 9312 7055 9364 7064
rect 9312 7021 9321 7055
rect 9321 7021 9355 7055
rect 9355 7021 9364 7055
rect 9312 7012 9364 7021
rect 7012 6944 7064 6996
rect 10232 6987 10284 6996
rect 6828 6876 6880 6928
rect 7472 6876 7524 6928
rect 10232 6953 10241 6987
rect 10241 6953 10275 6987
rect 10275 6953 10284 6987
rect 10232 6944 10284 6953
rect 12532 7089 12541 7123
rect 12541 7089 12575 7123
rect 12575 7089 12584 7123
rect 12532 7080 12584 7089
rect 13084 7012 13136 7064
rect 13636 7055 13688 7064
rect 13636 7021 13645 7055
rect 13645 7021 13679 7055
rect 13679 7021 13688 7055
rect 13636 7012 13688 7021
rect 14740 7216 14792 7268
rect 16948 7216 17000 7268
rect 17868 7259 17920 7268
rect 17868 7225 17877 7259
rect 17877 7225 17911 7259
rect 17911 7225 17920 7259
rect 17868 7216 17920 7225
rect 15660 7148 15712 7200
rect 18972 7216 19024 7268
rect 20260 7216 20312 7268
rect 16212 7123 16264 7132
rect 16212 7089 16221 7123
rect 16221 7089 16255 7123
rect 16255 7089 16264 7123
rect 16212 7080 16264 7089
rect 19248 7123 19300 7132
rect 19248 7089 19257 7123
rect 19257 7089 19291 7123
rect 19291 7089 19300 7123
rect 19248 7080 19300 7089
rect 20720 7123 20772 7132
rect 20720 7089 20729 7123
rect 20729 7089 20763 7123
rect 20763 7089 20772 7123
rect 20720 7080 20772 7089
rect 21548 7216 21600 7268
rect 21364 7123 21416 7132
rect 21364 7089 21373 7123
rect 21373 7089 21407 7123
rect 21407 7089 21416 7123
rect 21364 7080 21416 7089
rect 11244 6944 11296 6996
rect 14004 6944 14056 6996
rect 17776 7012 17828 7064
rect 21640 6987 21692 6996
rect 21640 6953 21668 6987
rect 21668 6953 21692 6987
rect 21640 6944 21692 6953
rect 13268 6876 13320 6928
rect 18972 6876 19024 6928
rect 22468 6876 22520 6928
rect 6092 6647 6144 6656
rect 6092 6613 6101 6647
rect 6101 6613 6135 6647
rect 6135 6613 6144 6647
rect 6092 6604 6144 6613
rect 7656 6647 7708 6656
rect 7656 6613 7665 6647
rect 7665 6613 7699 6647
rect 7699 6613 7708 6647
rect 7656 6604 7708 6613
rect 7840 6647 7892 6656
rect 7840 6613 7849 6647
rect 7849 6613 7883 6647
rect 7883 6613 7892 6647
rect 7840 6604 7892 6613
rect 11612 6672 11664 6724
rect 13268 6672 13320 6724
rect 20720 6672 20772 6724
rect 10416 6604 10468 6656
rect 13820 6604 13872 6656
rect 6828 6536 6880 6588
rect 8484 6579 8536 6588
rect 8484 6545 8512 6579
rect 8512 6545 8536 6579
rect 8484 6536 8536 6545
rect 11980 6536 12032 6588
rect 12348 6579 12400 6588
rect 12348 6545 12357 6579
rect 12357 6545 12391 6579
rect 12391 6545 12400 6579
rect 12348 6536 12400 6545
rect 7472 6468 7524 6520
rect 7840 6468 7892 6520
rect 8208 6511 8260 6520
rect 8208 6477 8217 6511
rect 8217 6477 8251 6511
rect 8251 6477 8260 6511
rect 8208 6468 8260 6477
rect 10324 6468 10376 6520
rect 14648 6536 14700 6588
rect 18328 6579 18380 6588
rect 18328 6545 18337 6579
rect 18337 6545 18371 6579
rect 18371 6545 18380 6579
rect 18328 6536 18380 6545
rect 20996 6536 21048 6588
rect 21824 6536 21876 6588
rect 22928 6604 22980 6656
rect 18604 6511 18656 6520
rect 6552 6375 6604 6384
rect 6552 6341 6561 6375
rect 6561 6341 6595 6375
rect 6595 6341 6604 6375
rect 6552 6332 6604 6341
rect 7748 6332 7800 6384
rect 9956 6332 10008 6384
rect 11244 6400 11296 6452
rect 18604 6477 18613 6511
rect 18613 6477 18647 6511
rect 18647 6477 18656 6511
rect 18604 6468 18656 6477
rect 19800 6468 19852 6520
rect 16212 6332 16264 6384
rect 21824 6332 21876 6384
rect 7012 6128 7064 6180
rect 7748 6171 7800 6180
rect 7748 6137 7757 6171
rect 7757 6137 7791 6171
rect 7791 6137 7800 6171
rect 7748 6128 7800 6137
rect 8392 6128 8444 6180
rect 9128 6128 9180 6180
rect 10324 6128 10376 6180
rect 12256 6128 12308 6180
rect 13820 6128 13872 6180
rect 18788 6128 18840 6180
rect 18972 6171 19024 6180
rect 18972 6137 18981 6171
rect 18981 6137 19015 6171
rect 19015 6137 19024 6171
rect 18972 6128 19024 6137
rect 19800 6171 19852 6180
rect 19800 6137 19809 6171
rect 19809 6137 19843 6171
rect 19843 6137 19852 6171
rect 19800 6128 19852 6137
rect 6552 6035 6604 6044
rect 6552 6001 6561 6035
rect 6561 6001 6595 6035
rect 6595 6001 6604 6035
rect 6552 5992 6604 6001
rect 7656 5992 7708 6044
rect 6736 5967 6788 5976
rect 6736 5933 6745 5967
rect 6745 5933 6779 5967
rect 6779 5933 6788 5967
rect 6736 5924 6788 5933
rect 12900 5924 12952 5976
rect 13268 5967 13320 5976
rect 13268 5933 13277 5967
rect 13277 5933 13311 5967
rect 13311 5933 13320 5967
rect 13268 5924 13320 5933
rect 14280 6035 14332 6044
rect 14280 6001 14289 6035
rect 14289 6001 14323 6035
rect 14323 6001 14332 6035
rect 14280 5992 14332 6001
rect 16212 6060 16264 6112
rect 18144 5992 18196 6044
rect 20076 5992 20128 6044
rect 22008 6128 22060 6180
rect 22192 6060 22244 6112
rect 21272 5992 21324 6044
rect 21824 6035 21876 6044
rect 21824 6001 21833 6035
rect 21833 6001 21867 6035
rect 21867 6001 21876 6035
rect 21824 5992 21876 6001
rect 16856 5967 16908 5976
rect 16856 5933 16865 5967
rect 16865 5933 16899 5967
rect 16899 5933 16908 5967
rect 16856 5924 16908 5933
rect 17776 5967 17828 5976
rect 17776 5933 17785 5967
rect 17785 5933 17819 5967
rect 17819 5933 17828 5967
rect 17776 5924 17828 5933
rect 20352 5924 20404 5976
rect 14096 5856 14148 5908
rect 10876 4156 10928 4208
rect 19156 4088 19208 4140
rect 20 144 72 196
rect 13452 144 13504 196
<< metal2 >>
rect 32 14811 60 27744
rect 18602 27734 18658 27743
rect 18602 27669 18658 27678
rect 8000 22060 8620 22080
rect 8000 22004 8042 22060
rect 8098 22004 8122 22060
rect 8178 22004 8202 22060
rect 8258 22004 8282 22060
rect 8338 22004 8362 22060
rect 8418 22004 8442 22060
rect 8498 22004 8522 22060
rect 8578 22004 8620 22060
rect 8000 21984 8620 22004
rect 13600 22060 14220 22080
rect 13600 22004 13642 22060
rect 13698 22004 13722 22060
rect 13778 22004 13802 22060
rect 13858 22004 13882 22060
rect 13938 22004 13962 22060
rect 14018 22004 14042 22060
rect 14098 22004 14122 22060
rect 14178 22004 14220 22060
rect 13600 21984 14220 22004
rect 15936 21820 15988 21826
rect 15936 21762 15988 21768
rect 18236 21820 18288 21826
rect 18616 21808 18644 27669
rect 21822 25294 21878 25303
rect 21822 25229 21878 25238
rect 19200 22060 19820 22080
rect 19200 22004 19242 22060
rect 19298 22004 19322 22060
rect 19378 22004 19402 22060
rect 19458 22004 19482 22060
rect 19538 22004 19562 22060
rect 19618 22004 19642 22060
rect 19698 22004 19722 22060
rect 19778 22004 19820 22060
rect 19200 21984 19820 22004
rect 20350 21878 20406 21887
rect 20350 21813 20406 21822
rect 21272 21820 21324 21826
rect 18616 21780 18736 21808
rect 18236 21762 18288 21768
rect 10324 21752 10376 21758
rect 10324 21694 10376 21700
rect 14280 21752 14332 21758
rect 14280 21694 14332 21700
rect 10140 21684 10192 21690
rect 10140 21626 10192 21632
rect 9240 21516 9860 21536
rect 9240 21460 9282 21516
rect 9338 21460 9362 21516
rect 9418 21460 9442 21516
rect 9498 21460 9522 21516
rect 9578 21460 9602 21516
rect 9658 21460 9682 21516
rect 9738 21460 9762 21516
rect 9818 21460 9860 21516
rect 9240 21440 9860 21460
rect 10152 21418 10180 21626
rect 10140 21412 10192 21418
rect 10140 21354 10192 21360
rect 9956 21072 10008 21078
rect 9956 21014 10008 21020
rect 8000 20972 8620 20992
rect 8000 20916 8042 20972
rect 8098 20916 8122 20972
rect 8178 20916 8202 20972
rect 8258 20916 8282 20972
rect 8338 20916 8362 20972
rect 8418 20916 8442 20972
rect 8498 20916 8522 20972
rect 8578 20916 8620 20972
rect 8000 20896 8620 20916
rect 7564 20732 7616 20738
rect 7564 20674 7616 20680
rect 7288 20664 7340 20670
rect 7288 20606 7340 20612
rect 6828 20188 6880 20194
rect 7300 20176 7328 20606
rect 6880 20148 7328 20176
rect 6828 20130 6880 20136
rect 6920 20052 6972 20058
rect 6920 19994 6972 20000
rect 6736 19984 6788 19990
rect 6736 19926 6788 19932
rect 6748 19768 6776 19926
rect 6656 19740 6776 19768
rect 6656 18748 6684 19740
rect 6932 19242 6960 19994
rect 7012 19644 7064 19650
rect 7012 19586 7064 19592
rect 6920 19236 6972 19242
rect 6920 19178 6972 19184
rect 6920 19032 6972 19038
rect 6920 18974 6972 18980
rect 6932 18816 6960 18974
rect 7024 18816 7052 19586
rect 6932 18788 7052 18816
rect 6656 18720 6776 18748
rect 6748 18562 6776 18720
rect 6736 18556 6788 18562
rect 6736 18498 6788 18504
rect 6552 18352 6604 18358
rect 6552 18294 6604 18300
rect 6564 17406 6592 18294
rect 6932 17950 6960 18788
rect 6920 17944 6972 17950
rect 6920 17886 6972 17892
rect 6552 17400 6604 17406
rect 6552 17342 6604 17348
rect 6828 17264 6880 17270
rect 6828 17206 6880 17212
rect 6840 17048 6868 17206
rect 6656 17020 6868 17048
rect 6184 16380 6236 16386
rect 6184 16322 6236 16328
rect 6196 15434 6224 16322
rect 6656 15824 6684 17020
rect 6932 16386 6960 17886
rect 7104 17808 7156 17814
rect 7104 17750 7156 17756
rect 6920 16380 6972 16386
rect 6920 16322 6972 16328
rect 6932 15978 6960 16322
rect 7116 16031 7144 17750
rect 7300 17474 7328 20148
rect 7576 19786 7604 20674
rect 9968 20534 9996 21014
rect 9128 20528 9180 20534
rect 9128 20470 9180 20476
rect 9956 20528 10008 20534
rect 9956 20470 10008 20476
rect 8760 19984 8812 19990
rect 8760 19926 8812 19932
rect 8944 19984 8996 19990
rect 8944 19926 8996 19932
rect 8000 19884 8620 19904
rect 8000 19828 8042 19884
rect 8098 19828 8122 19884
rect 8178 19828 8202 19884
rect 8258 19828 8282 19884
rect 8338 19828 8362 19884
rect 8418 19828 8442 19884
rect 8498 19828 8522 19884
rect 8578 19828 8620 19884
rect 8000 19808 8620 19828
rect 7564 19780 7616 19786
rect 7564 19722 7616 19728
rect 8772 19718 8800 19926
rect 8956 19786 8984 19926
rect 9140 19786 9168 20470
rect 9240 20428 9860 20448
rect 9240 20372 9282 20428
rect 9338 20372 9362 20428
rect 9418 20372 9442 20428
rect 9498 20372 9522 20428
rect 9578 20372 9602 20428
rect 9658 20372 9682 20428
rect 9738 20372 9762 20428
rect 9818 20372 9860 20428
rect 9240 20352 9860 20372
rect 8944 19780 8996 19786
rect 8944 19722 8996 19728
rect 9128 19780 9180 19786
rect 9128 19722 9180 19728
rect 8760 19712 8812 19718
rect 8760 19654 8812 19660
rect 7932 19508 7984 19514
rect 7932 19450 7984 19456
rect 7472 18080 7524 18086
rect 7472 18022 7524 18028
rect 7484 17474 7512 18022
rect 7288 17468 7340 17474
rect 7288 17410 7340 17416
rect 7472 17468 7524 17474
rect 7472 17410 7524 17416
rect 7300 16386 7328 17410
rect 7944 16454 7972 19450
rect 8760 19440 8812 19446
rect 8760 19382 8812 19388
rect 8000 18796 8620 18816
rect 8000 18740 8042 18796
rect 8098 18740 8122 18796
rect 8178 18740 8202 18796
rect 8258 18740 8282 18796
rect 8338 18740 8362 18796
rect 8418 18740 8442 18796
rect 8498 18740 8522 18796
rect 8578 18740 8620 18796
rect 8000 18720 8620 18740
rect 8772 18698 8800 19382
rect 8956 19106 8984 19722
rect 8944 19100 8996 19106
rect 8944 19042 8996 19048
rect 8760 18692 8812 18698
rect 8760 18634 8812 18640
rect 9140 18562 9168 19722
rect 9968 19446 9996 20470
rect 10336 20330 10364 21694
rect 10508 21616 10560 21622
rect 10508 21558 10560 21564
rect 10520 20856 10548 21558
rect 10968 21208 11020 21214
rect 10968 21150 11020 21156
rect 13084 21208 13136 21214
rect 13084 21150 13136 21156
rect 13360 21208 13412 21214
rect 13360 21150 13412 21156
rect 10891 20868 10943 20874
rect 10520 20828 10891 20856
rect 10891 20810 10943 20816
rect 10876 20732 10928 20738
rect 10704 20692 10876 20720
rect 10324 20324 10376 20330
rect 10324 20266 10376 20272
rect 10336 20176 10364 20266
rect 10704 20188 10732 20692
rect 10876 20674 10928 20680
rect 10336 20148 10548 20176
rect 10232 20052 10284 20058
rect 10232 19994 10284 20000
rect 10244 19786 10272 19994
rect 10232 19780 10284 19786
rect 10232 19722 10284 19728
rect 10520 19650 10548 20148
rect 10686 20136 10692 20188
rect 10744 20136 10750 20188
rect 10508 19644 10560 19650
rect 10508 19586 10560 19592
rect 10324 19508 10376 19514
rect 10324 19450 10376 19456
rect 9956 19440 10008 19446
rect 9956 19382 10008 19388
rect 9240 19340 9860 19360
rect 9240 19284 9282 19340
rect 9338 19284 9362 19340
rect 9418 19284 9442 19340
rect 9498 19284 9522 19340
rect 9578 19284 9602 19340
rect 9658 19284 9682 19340
rect 9738 19284 9762 19340
rect 9818 19284 9860 19340
rect 9240 19264 9860 19284
rect 9968 19106 9996 19382
rect 10336 19242 10364 19450
rect 10324 19236 10376 19242
rect 10324 19178 10376 19184
rect 9956 19100 10008 19106
rect 9956 19042 10008 19048
rect 10232 19032 10284 19038
rect 10232 18974 10284 18980
rect 9956 18896 10008 18902
rect 9956 18838 10008 18844
rect 9128 18556 9180 18562
rect 9128 18498 9180 18504
rect 8668 18488 8720 18494
rect 8668 18430 8720 18436
rect 9036 18488 9088 18494
rect 9036 18430 9088 18436
rect 8000 17708 8620 17728
rect 8000 17652 8042 17708
rect 8098 17652 8122 17708
rect 8178 17652 8202 17708
rect 8258 17652 8282 17708
rect 8338 17652 8362 17708
rect 8418 17652 8442 17708
rect 8498 17652 8522 17708
rect 8578 17652 8620 17708
rect 8000 17632 8620 17652
rect 8680 17524 8708 18430
rect 8852 18352 8904 18358
rect 8852 18294 8904 18300
rect 8864 18154 8892 18294
rect 9048 18154 9076 18430
rect 9240 18252 9860 18272
rect 9240 18196 9282 18252
rect 9338 18196 9362 18252
rect 9418 18196 9442 18252
rect 9498 18196 9522 18252
rect 9578 18196 9602 18252
rect 9658 18196 9682 18252
rect 9738 18196 9762 18252
rect 9818 18196 9860 18252
rect 9240 18176 9860 18196
rect 8852 18148 8904 18154
rect 8852 18090 8904 18096
rect 9036 18148 9088 18154
rect 9036 18090 9088 18096
rect 9968 18018 9996 18838
rect 9956 18012 10008 18018
rect 9956 17954 10008 17960
rect 9588 17944 9640 17950
rect 9588 17886 9640 17892
rect 9772 17944 9824 17950
rect 10244 17944 10272 18974
rect 10704 18494 10732 20136
rect 10980 19038 11008 21150
rect 12624 21072 12676 21078
rect 12624 21014 12676 21020
rect 12636 20874 12664 21014
rect 12609 20868 12664 20874
rect 12661 20828 12664 20868
rect 12609 20810 12661 20816
rect 13096 20806 13124 21150
rect 13084 20800 13136 20806
rect 13084 20742 13136 20748
rect 12624 20732 12676 20738
rect 12624 20674 12676 20680
rect 11520 20596 11572 20602
rect 11520 20538 11572 20544
rect 11532 19106 11560 20538
rect 12636 20126 12664 20674
rect 13372 20534 13400 21150
rect 14292 21146 14320 21694
rect 15470 21564 15476 21616
rect 15528 21564 15534 21616
rect 14840 21516 15460 21536
rect 14840 21460 14882 21516
rect 14938 21460 14962 21516
rect 15018 21460 15042 21516
rect 15098 21460 15122 21516
rect 15178 21460 15202 21516
rect 15258 21460 15282 21516
rect 15338 21460 15362 21516
rect 15418 21460 15460 21516
rect 14840 21440 15460 21460
rect 14464 21208 14516 21214
rect 14464 21150 14516 21156
rect 15108 21208 15160 21214
rect 15108 21150 15160 21156
rect 14280 21140 14332 21146
rect 14280 21082 14332 21088
rect 13600 20972 14220 20992
rect 13600 20916 13642 20972
rect 13698 20916 13722 20972
rect 13778 20916 13802 20972
rect 13858 20916 13882 20972
rect 13938 20916 13962 20972
rect 14018 20916 14042 20972
rect 14098 20916 14122 20972
rect 14178 20916 14220 20972
rect 13600 20896 14220 20916
rect 14292 20874 14320 21082
rect 14372 21072 14424 21078
rect 14372 21014 14424 21020
rect 14280 20868 14332 20874
rect 14280 20810 14332 20816
rect 13360 20528 13412 20534
rect 13360 20470 13412 20476
rect 12624 20120 12676 20126
rect 13372 20108 13400 20470
rect 12624 20062 12676 20068
rect 13280 20080 13400 20108
rect 12348 20052 12400 20058
rect 12348 19994 12400 20000
rect 12360 19650 12388 19994
rect 12636 19650 12664 20062
rect 12164 19644 12216 19650
rect 12164 19586 12216 19592
rect 12348 19644 12400 19650
rect 12348 19586 12400 19592
rect 12624 19644 12676 19650
rect 13280 19632 13308 20080
rect 13452 19984 13504 19990
rect 13452 19926 13504 19932
rect 13464 19768 13492 19926
rect 13600 19884 14220 19904
rect 13600 19828 13642 19884
rect 13698 19828 13722 19884
rect 13778 19828 13802 19884
rect 13858 19828 13882 19884
rect 13938 19828 13962 19884
rect 14018 19828 14042 19884
rect 14098 19828 14122 19884
rect 14178 19828 14220 19884
rect 13600 19808 14220 19828
rect 13464 19740 13584 19768
rect 13556 19632 13584 19740
rect 13280 19604 13400 19632
rect 13556 19604 13676 19632
rect 12624 19586 12676 19592
rect 11980 19508 12032 19514
rect 11980 19450 12032 19456
rect 11796 19440 11848 19446
rect 11796 19382 11848 19388
rect 11520 19100 11572 19106
rect 11520 19042 11572 19048
rect 11808 19038 11836 19382
rect 11992 19106 12020 19450
rect 12176 19428 12204 19586
rect 12716 19576 12768 19582
rect 12716 19518 12768 19524
rect 12176 19400 12296 19428
rect 12072 19168 12124 19174
rect 12072 19110 12124 19116
rect 11980 19100 12032 19106
rect 11980 19042 12032 19048
rect 10968 19032 11020 19038
rect 10968 18974 11020 18980
rect 11612 19032 11664 19038
rect 11612 18974 11664 18980
rect 11796 19032 11848 19038
rect 11796 18974 11848 18980
rect 10968 18896 11020 18902
rect 10968 18838 11020 18844
rect 10980 18562 11008 18838
rect 10968 18556 11020 18562
rect 10968 18498 11020 18504
rect 10692 18488 10744 18494
rect 10692 18430 10744 18436
rect 10226 17892 10232 17944
rect 10284 17892 10290 17944
rect 9772 17886 9824 17892
rect 9600 17610 9628 17886
rect 9588 17604 9640 17610
rect 9588 17546 9640 17552
rect 9784 17542 9812 17886
rect 10244 17864 10272 17892
rect 9968 17836 10272 17864
rect 8588 17496 8708 17524
rect 9772 17536 9824 17542
rect 8588 16776 8616 17496
rect 9772 17478 9824 17484
rect 8852 17468 8904 17474
rect 8852 17410 8904 17416
rect 8588 16748 8708 16776
rect 8000 16620 8620 16640
rect 8000 16564 8042 16620
rect 8098 16564 8122 16620
rect 8178 16564 8202 16620
rect 8258 16564 8282 16620
rect 8338 16564 8362 16620
rect 8418 16564 8442 16620
rect 8498 16564 8522 16620
rect 8578 16564 8620 16620
rect 8000 16544 8620 16564
rect 7932 16448 7984 16454
rect 7932 16390 7984 16396
rect 7288 16380 7340 16386
rect 7288 16322 7340 16328
rect 7102 16022 7158 16031
rect 6920 15972 6972 15978
rect 7102 15957 7158 15966
rect 6920 15914 6972 15920
rect 6656 15796 6868 15824
rect 6184 15428 6236 15434
rect 6184 15370 6236 15376
rect 6840 15298 6868 15796
rect 7300 15787 7328 16322
rect 7470 16022 7526 16031
rect 7470 15957 7526 15966
rect 8680 15960 8708 16748
rect 8864 16522 8892 17410
rect 9036 17264 9088 17270
rect 9036 17206 9088 17212
rect 8852 16516 8904 16522
rect 8852 16458 8904 16464
rect 9048 16386 9076 17206
rect 9240 17164 9860 17184
rect 9240 17108 9282 17164
rect 9338 17108 9362 17164
rect 9418 17108 9442 17164
rect 9498 17108 9522 17164
rect 9578 17108 9602 17164
rect 9658 17108 9682 17164
rect 9738 17108 9762 17164
rect 9818 17108 9860 17164
rect 9240 17088 9860 17108
rect 9968 16504 9996 17836
rect 10324 17808 10376 17814
rect 10324 17750 10376 17756
rect 10140 17468 10192 17474
rect 10140 17410 10192 17416
rect 10152 17066 10180 17410
rect 10336 17406 10364 17750
rect 10704 17474 10732 18430
rect 11336 18012 11388 18018
rect 11336 17954 11388 17960
rect 10968 17808 11020 17814
rect 10968 17750 11020 17756
rect 10692 17468 10744 17474
rect 10692 17410 10744 17416
rect 10324 17400 10376 17406
rect 10324 17342 10376 17348
rect 10324 17264 10376 17270
rect 10324 17206 10376 17212
rect 10140 17060 10192 17066
rect 10140 17002 10192 17008
rect 10336 16862 10364 17206
rect 10704 16912 10732 17410
rect 10876 16924 10928 16930
rect 10704 16884 10876 16912
rect 10324 16856 10376 16862
rect 10324 16798 10376 16804
rect 9876 16476 9996 16504
rect 9036 16380 9088 16386
rect 9036 16322 9088 16328
rect 9876 16318 9904 16476
rect 8852 16312 8904 16318
rect 8852 16254 8904 16260
rect 9864 16312 9916 16318
rect 9864 16254 9916 16260
rect 8864 15978 8892 16254
rect 9220 16244 9272 16250
rect 9140 16204 9220 16232
rect 9036 16176 9088 16182
rect 9036 16118 9088 16124
rect 8852 15972 8904 15978
rect 7286 15778 7342 15787
rect 7196 15768 7248 15774
rect 7196 15710 7248 15716
rect 7484 15774 7512 15957
rect 8680 15932 8800 15960
rect 8666 15778 8722 15787
rect 7286 15713 7342 15722
rect 7472 15768 7524 15774
rect 7208 15552 7236 15710
rect 7300 15552 7328 15713
rect 7472 15710 7524 15716
rect 7932 15768 7984 15774
rect 7932 15710 7984 15716
rect 8666 15713 8722 15722
rect 7208 15524 7328 15552
rect 6828 15292 6880 15298
rect 6828 15234 6880 15240
rect 7300 14872 7328 15524
rect 7944 15298 7972 15710
rect 8000 15532 8620 15552
rect 8000 15476 8042 15532
rect 8098 15476 8122 15532
rect 8178 15476 8202 15532
rect 8258 15476 8282 15532
rect 8338 15476 8362 15532
rect 8418 15476 8442 15532
rect 8498 15476 8522 15532
rect 8578 15476 8620 15532
rect 8000 15456 8620 15476
rect 8680 15298 8708 15713
rect 8772 15638 8800 15932
rect 8852 15914 8904 15920
rect 9048 15910 9076 16118
rect 9140 15960 9168 16204
rect 9220 16186 9272 16192
rect 9240 16076 9860 16096
rect 9240 16020 9282 16076
rect 9338 16020 9362 16076
rect 9418 16020 9442 16076
rect 9498 16020 9522 16076
rect 9578 16020 9602 16076
rect 9658 16020 9682 16076
rect 9738 16020 9762 16076
rect 9818 16020 9860 16076
rect 9240 16000 9860 16020
rect 9140 15932 9260 15960
rect 9036 15904 9088 15910
rect 9036 15846 9088 15852
rect 8944 15768 8996 15774
rect 8944 15710 8996 15716
rect 8760 15632 8812 15638
rect 8760 15574 8812 15580
rect 8956 15298 8984 15710
rect 9232 15434 9260 15932
rect 9968 15892 9996 16476
rect 10600 16380 10652 16386
rect 10704 16368 10732 16884
rect 10876 16866 10928 16872
rect 10980 16454 11008 17750
rect 11348 17066 11376 17954
rect 11336 17060 11388 17066
rect 11336 17002 11388 17008
rect 11624 16862 11652 18974
rect 12084 18884 12112 19110
rect 12268 18884 12296 19400
rect 12728 19360 12756 19518
rect 13176 19440 13228 19446
rect 13176 19382 13228 19388
rect 12728 19332 12848 19360
rect 12820 19224 12848 19332
rect 11992 18856 12112 18884
rect 12176 18856 12296 18884
rect 12636 19196 12848 19224
rect 11992 18272 12020 18856
rect 12176 18698 12204 18856
rect 12164 18692 12216 18698
rect 12164 18634 12216 18640
rect 11992 18244 12112 18272
rect 11980 18080 12032 18086
rect 11980 18022 12032 18028
rect 11992 17066 12020 18022
rect 12084 18018 12112 18244
rect 12072 18012 12124 18018
rect 12072 17954 12124 17960
rect 12176 17950 12204 18634
rect 12636 18272 12664 19196
rect 12992 19168 13044 19174
rect 12992 19110 13044 19116
rect 13004 18426 13032 19110
rect 13188 18698 13216 19382
rect 13372 19038 13400 19604
rect 13648 19088 13676 19604
rect 14188 19440 14240 19446
rect 14188 19382 14240 19388
rect 14200 19174 14228 19382
rect 14188 19168 14240 19174
rect 14188 19110 14240 19116
rect 13556 19060 13676 19088
rect 13360 19032 13412 19038
rect 13360 18974 13412 18980
rect 13556 18952 13584 19060
rect 13464 18924 13584 18952
rect 14200 18952 14228 19110
rect 14384 18952 14412 21014
rect 14476 20670 14504 21150
rect 14740 21072 14792 21078
rect 14740 21014 14792 21020
rect 14464 20664 14516 20670
rect 14464 20606 14516 20612
rect 14752 19990 14780 21014
rect 15120 20738 15148 21150
rect 15488 20874 15516 21564
rect 15948 21418 15976 21762
rect 16488 21752 16540 21758
rect 16488 21694 16540 21700
rect 15936 21412 15988 21418
rect 15936 21354 15988 21360
rect 16500 21282 16528 21694
rect 17408 21616 17460 21622
rect 17408 21558 17460 21564
rect 17132 21344 17184 21350
rect 17132 21286 17184 21292
rect 16488 21276 16540 21282
rect 16488 21218 16540 21224
rect 15936 21208 15988 21214
rect 15936 21150 15988 21156
rect 15476 20868 15528 20874
rect 15476 20810 15528 20816
rect 15108 20732 15160 20738
rect 15108 20674 15160 20680
rect 15948 20670 15976 21150
rect 16120 21140 16172 21146
rect 16120 21082 16172 21088
rect 15936 20664 15988 20670
rect 15936 20606 15988 20612
rect 15470 20476 15476 20528
rect 15528 20476 15534 20528
rect 14840 20428 15460 20448
rect 14840 20372 14882 20428
rect 14938 20372 14962 20428
rect 15018 20372 15042 20428
rect 15098 20372 15122 20428
rect 15178 20372 15202 20428
rect 15258 20372 15282 20428
rect 15338 20372 15362 20428
rect 15418 20372 15460 20428
rect 14840 20352 15460 20372
rect 15488 20058 15516 20476
rect 15948 20179 15976 20606
rect 15934 20170 15990 20179
rect 15934 20105 15936 20114
rect 15988 20105 15990 20114
rect 15936 20062 15988 20068
rect 15476 20052 15528 20058
rect 15476 19994 15528 20000
rect 14740 19984 14792 19990
rect 14740 19926 14792 19932
rect 16028 19984 16080 19990
rect 16028 19926 16080 19932
rect 16040 19632 16068 19926
rect 16132 19786 16160 21082
rect 16212 21072 16264 21078
rect 16212 21014 16264 21020
rect 16224 20806 16252 21014
rect 16212 20800 16264 20806
rect 16212 20742 16264 20748
rect 17144 20534 17172 21286
rect 17420 21282 17448 21558
rect 18248 21418 18276 21762
rect 18420 21684 18472 21690
rect 18420 21626 18472 21632
rect 18236 21412 18288 21418
rect 18236 21354 18288 21360
rect 17408 21276 17460 21282
rect 17408 21218 17460 21224
rect 18432 21146 18460 21626
rect 18708 21264 18736 21780
rect 20364 21758 20392 21813
rect 21272 21762 21324 21768
rect 19616 21752 19668 21758
rect 19616 21694 19668 21700
rect 20352 21752 20404 21758
rect 20352 21694 20404 21700
rect 21088 21752 21140 21758
rect 21088 21694 21140 21700
rect 19156 21616 19208 21622
rect 19156 21558 19208 21564
rect 19168 21350 19196 21558
rect 19156 21344 19208 21350
rect 19156 21286 19208 21292
rect 19628 21282 19656 21694
rect 19892 21616 19944 21622
rect 19892 21558 19944 21564
rect 19984 21616 20036 21622
rect 19984 21558 20036 21564
rect 18616 21236 18736 21264
rect 19616 21276 19668 21282
rect 18420 21140 18472 21146
rect 18420 21082 18472 21088
rect 17684 21072 17736 21078
rect 17684 21014 17736 21020
rect 17696 20534 17724 21014
rect 17132 20528 17184 20534
rect 17132 20470 17184 20476
rect 17684 20528 17736 20534
rect 17684 20470 17736 20476
rect 16304 20052 16356 20058
rect 16304 19994 16356 20000
rect 16316 19786 16344 19994
rect 16120 19780 16172 19786
rect 16120 19722 16172 19728
rect 16304 19780 16356 19786
rect 16304 19722 16356 19728
rect 16856 19644 16908 19650
rect 16040 19604 16160 19632
rect 14556 19440 14608 19446
rect 14556 19382 14608 19388
rect 14568 19106 14596 19382
rect 14840 19340 15460 19360
rect 14840 19284 14882 19340
rect 14938 19284 14962 19340
rect 15018 19284 15042 19340
rect 15098 19284 15122 19340
rect 15178 19284 15202 19340
rect 15258 19284 15282 19340
rect 15338 19284 15362 19340
rect 15418 19284 15460 19340
rect 14840 19264 15460 19284
rect 14832 19168 14884 19174
rect 14832 19110 14884 19116
rect 14556 19100 14608 19106
rect 14556 19042 14608 19048
rect 14200 18924 14320 18952
rect 14384 18924 14596 18952
rect 13176 18692 13228 18698
rect 13176 18634 13228 18640
rect 13464 18562 13492 18924
rect 13600 18796 14220 18816
rect 13600 18740 13642 18796
rect 13698 18740 13722 18796
rect 13778 18740 13802 18796
rect 13858 18740 13882 18796
rect 13938 18740 13962 18796
rect 14018 18740 14042 18796
rect 14098 18740 14122 18796
rect 14178 18740 14220 18796
rect 13600 18720 14220 18740
rect 13452 18556 13504 18562
rect 13452 18498 13504 18504
rect 12992 18420 13044 18426
rect 12992 18362 13044 18368
rect 12636 18244 12848 18272
rect 12256 18012 12308 18018
rect 12256 17954 12308 17960
rect 12164 17944 12216 17950
rect 12164 17886 12216 17892
rect 12268 17610 12296 17954
rect 12256 17604 12308 17610
rect 12256 17546 12308 17552
rect 12820 17456 12848 18244
rect 13268 18148 13320 18154
rect 13188 18108 13268 18136
rect 12992 17468 13044 17474
rect 12820 17428 12992 17456
rect 11980 17060 12032 17066
rect 11980 17002 12032 17008
rect 12072 16992 12124 16998
rect 12072 16934 12124 16940
rect 11612 16856 11664 16862
rect 11612 16798 11664 16804
rect 11796 16856 11848 16862
rect 11796 16798 11848 16804
rect 11888 16856 11940 16862
rect 11888 16798 11940 16804
rect 11624 16522 11652 16798
rect 11612 16516 11664 16522
rect 11612 16458 11664 16464
rect 10968 16448 11020 16454
rect 10968 16390 11020 16396
rect 10652 16340 10732 16368
rect 10600 16322 10652 16328
rect 10232 16244 10284 16250
rect 10232 16186 10284 16192
rect 10048 16176 10100 16182
rect 10048 16118 10100 16124
rect 9876 15864 9996 15892
rect 9494 15778 9550 15787
rect 9494 15716 9496 15722
rect 9548 15716 9550 15722
rect 9494 15713 9550 15716
rect 9496 15710 9548 15713
rect 9220 15428 9272 15434
rect 9220 15370 9272 15376
rect 7932 15292 7984 15298
rect 7932 15234 7984 15240
rect 8668 15292 8720 15298
rect 8668 15234 8720 15240
rect 8944 15292 8996 15298
rect 8944 15234 8996 15240
rect 9876 15144 9904 15864
rect 10060 15774 10088 16118
rect 10244 15824 10272 16186
rect 10152 15796 10272 15824
rect 10048 15768 10100 15774
rect 10048 15710 10100 15716
rect 9876 15116 9996 15144
rect 9240 14988 9860 15008
rect 9240 14932 9282 14988
rect 9338 14932 9362 14988
rect 9418 14932 9442 14988
rect 9498 14932 9522 14988
rect 9578 14932 9602 14988
rect 9658 14932 9682 14988
rect 9738 14932 9762 14988
rect 9818 14932 9860 14988
rect 9240 14912 9860 14932
rect 6932 14844 7328 14872
rect 18 14802 74 14811
rect 6932 14754 6960 14844
rect 18 14737 74 14746
rect 6920 14748 6972 14754
rect 6920 14690 6972 14696
rect 6736 14680 6788 14686
rect 6736 14622 6788 14628
rect 6552 14544 6604 14550
rect 6552 14486 6604 14492
rect 6564 14210 6592 14486
rect 6552 14204 6604 14210
rect 6552 14146 6604 14152
rect 5814 13826 5870 13835
rect 6748 13802 6776 14622
rect 7300 14210 7328 14844
rect 9036 14816 9088 14822
rect 9036 14758 9088 14764
rect 8000 14444 8620 14464
rect 8000 14388 8042 14444
rect 8098 14388 8122 14444
rect 8178 14388 8202 14444
rect 8258 14388 8282 14444
rect 8338 14388 8362 14444
rect 8418 14388 8442 14444
rect 8498 14388 8522 14444
rect 8578 14388 8620 14444
rect 8000 14368 8620 14388
rect 7288 14204 7340 14210
rect 7288 14146 7340 14152
rect 7932 14204 7984 14210
rect 7932 14146 7984 14152
rect 6920 14136 6972 14142
rect 6920 14078 6972 14084
rect 5814 13761 5870 13770
rect 6736 13796 6788 13802
rect 5828 13648 5856 13761
rect 6736 13738 6788 13744
rect 6368 13660 6420 13666
rect 5828 13620 5948 13648
rect 5920 7546 5948 13620
rect 6368 13602 6420 13608
rect 6184 13456 6236 13462
rect 6184 13398 6236 13404
rect 6196 11422 6224 13398
rect 6380 13122 6408 13602
rect 6932 13598 6960 14078
rect 6920 13592 6972 13598
rect 6920 13534 6972 13540
rect 6736 13524 6788 13530
rect 6736 13466 6788 13472
rect 6748 13122 6776 13466
rect 6932 13258 6960 13534
rect 6920 13252 6972 13258
rect 6920 13194 6972 13200
rect 6368 13116 6420 13122
rect 6368 13058 6420 13064
rect 6736 13116 6788 13122
rect 6736 13058 6788 13064
rect 6380 12374 6408 13058
rect 7300 13054 7328 14146
rect 7944 13802 7972 14146
rect 9048 13802 9076 14758
rect 9128 14000 9180 14006
rect 9128 13942 9180 13948
rect 7932 13796 7984 13802
rect 7932 13738 7984 13744
rect 9036 13796 9088 13802
rect 9036 13738 9088 13744
rect 9140 13666 9168 13942
rect 9240 13900 9860 13920
rect 9240 13844 9282 13900
rect 9338 13844 9362 13900
rect 9418 13844 9442 13900
rect 9498 13844 9522 13900
rect 9578 13844 9602 13900
rect 9658 13844 9682 13900
rect 9738 13844 9762 13900
rect 9818 13844 9860 13900
rect 9240 13824 9860 13844
rect 9128 13660 9180 13666
rect 9128 13602 9180 13608
rect 9496 13592 9548 13598
rect 9496 13534 9548 13540
rect 8000 13356 8620 13376
rect 8000 13300 8042 13356
rect 8098 13300 8122 13356
rect 8178 13300 8202 13356
rect 8258 13300 8282 13356
rect 8338 13300 8362 13356
rect 8418 13300 8442 13356
rect 8498 13300 8522 13356
rect 8578 13300 8620 13356
rect 8000 13280 8620 13300
rect 9508 13258 9536 13534
rect 9496 13252 9548 13258
rect 9968 13240 9996 15116
rect 10152 14890 10180 15796
rect 10704 15787 10732 16340
rect 11612 16380 11664 16386
rect 11612 16322 11664 16328
rect 10968 16176 11020 16182
rect 10968 16118 11020 16124
rect 10690 15778 10746 15787
rect 10690 15713 10746 15722
rect 10784 15768 10836 15774
rect 10784 15710 10836 15716
rect 10416 15700 10468 15706
rect 10416 15642 10468 15648
rect 10232 15632 10284 15638
rect 10232 15574 10284 15580
rect 10244 15298 10272 15574
rect 10232 15292 10284 15298
rect 10232 15234 10284 15240
rect 10428 15230 10456 15642
rect 10796 15298 10824 15710
rect 10784 15292 10836 15298
rect 10784 15234 10836 15240
rect 10416 15224 10468 15230
rect 10416 15166 10468 15172
rect 10692 15224 10744 15230
rect 10692 15166 10744 15172
rect 10428 14890 10456 15166
rect 10704 14890 10732 15166
rect 10140 14884 10192 14890
rect 10140 14826 10192 14832
rect 10416 14884 10468 14890
rect 10416 14826 10468 14832
rect 10692 14884 10744 14890
rect 10692 14826 10744 14832
rect 10598 14802 10654 14811
rect 10598 14737 10654 14746
rect 10612 14346 10640 14737
rect 10980 14686 11008 16118
rect 11152 15972 11204 15978
rect 11152 15914 11204 15920
rect 11164 15756 11192 15914
rect 11624 15774 11652 16322
rect 11808 15978 11836 16798
rect 11900 16250 11928 16798
rect 12084 16776 12112 16934
rect 12084 16748 12296 16776
rect 11980 16380 12032 16386
rect 11980 16322 12032 16328
rect 11888 16244 11940 16250
rect 11888 16186 11940 16192
rect 11796 15972 11848 15978
rect 11796 15914 11848 15920
rect 11992 15824 12020 16322
rect 12268 15960 12296 16748
rect 12820 16454 12848 17428
rect 12992 17410 13044 17416
rect 12900 16924 12952 16930
rect 12952 16884 13032 16912
rect 12900 16866 12952 16872
rect 12808 16448 12860 16454
rect 12808 16390 12860 16396
rect 12716 16176 12768 16182
rect 12716 16118 12768 16124
rect 11900 15796 12020 15824
rect 12084 15932 12296 15960
rect 11612 15768 11664 15774
rect 11164 15728 11284 15756
rect 11256 15280 11284 15728
rect 11612 15710 11664 15716
rect 11900 15298 11928 15796
rect 12084 15366 12112 15932
rect 12348 15768 12400 15774
rect 12348 15710 12400 15716
rect 12072 15360 12124 15366
rect 12072 15302 12124 15308
rect 11164 15252 11284 15280
rect 11888 15292 11940 15298
rect 10876 14680 10928 14686
rect 10876 14622 10928 14628
rect 10968 14680 11020 14686
rect 10968 14622 11020 14628
rect 10600 14340 10652 14346
rect 10600 14282 10652 14288
rect 10888 13920 10916 14622
rect 11164 14210 11192 15252
rect 11888 15234 11940 15240
rect 11796 15224 11848 15230
rect 11796 15166 11848 15172
rect 11336 15088 11388 15094
rect 11336 15030 11388 15036
rect 11348 14872 11376 15030
rect 11348 14844 11468 14872
rect 11152 14204 11204 14210
rect 11152 14146 11204 14152
rect 11440 14056 11468 14844
rect 11808 14346 11836 15166
rect 12360 14686 12388 15710
rect 12440 15700 12492 15706
rect 12728 15688 12756 16118
rect 13004 15978 13032 16884
rect 13084 16720 13136 16726
rect 13084 16662 13136 16668
rect 13096 16522 13124 16662
rect 13084 16516 13136 16522
rect 13084 16458 13136 16464
rect 12992 15972 13044 15978
rect 12992 15914 13044 15920
rect 12492 15660 12756 15688
rect 12440 15642 12492 15648
rect 12624 15292 12676 15298
rect 12544 15252 12624 15280
rect 12348 14680 12400 14686
rect 12348 14622 12400 14628
rect 11796 14340 11848 14346
rect 11796 14282 11848 14288
rect 12360 14142 12388 14622
rect 12348 14136 12400 14142
rect 12348 14078 12400 14084
rect 11348 14028 11468 14056
rect 10888 13892 11008 13920
rect 10232 13728 10284 13734
rect 10232 13670 10284 13676
rect 10784 13728 10836 13734
rect 10784 13670 10836 13676
rect 9968 13212 10088 13240
rect 9496 13194 9548 13200
rect 7288 13048 7340 13054
rect 7288 12990 7340 12996
rect 6552 12504 6604 12510
rect 6552 12446 6604 12452
rect 6368 12368 6420 12374
rect 6368 12310 6420 12316
rect 6564 12034 6592 12446
rect 6736 12436 6788 12442
rect 6736 12378 6788 12384
rect 6748 12170 6776 12378
rect 6736 12164 6788 12170
rect 6736 12106 6788 12112
rect 6552 12028 6604 12034
rect 6552 11970 6604 11976
rect 6564 11880 6592 11970
rect 7300 11960 7328 12990
rect 10060 12986 10088 13212
rect 10048 12980 10100 12986
rect 10048 12922 10100 12928
rect 9240 12812 9860 12832
rect 9240 12756 9282 12812
rect 9338 12756 9362 12812
rect 9418 12756 9442 12812
rect 9498 12756 9522 12812
rect 9578 12756 9602 12812
rect 9658 12756 9682 12812
rect 9738 12756 9762 12812
rect 9818 12756 9860 12812
rect 9240 12736 9860 12756
rect 10060 12628 10088 12922
rect 10244 12714 10272 13670
rect 10692 13456 10744 13462
rect 10692 13398 10744 13404
rect 10704 13054 10732 13398
rect 10796 13190 10824 13670
rect 10980 13598 11008 13892
rect 11348 13802 11376 14028
rect 11796 14000 11848 14006
rect 11796 13942 11848 13948
rect 11336 13796 11388 13802
rect 11336 13738 11388 13744
rect 10968 13592 11020 13598
rect 10968 13534 11020 13540
rect 11612 13456 11664 13462
rect 11612 13398 11664 13404
rect 11624 13240 11652 13398
rect 11532 13212 11652 13240
rect 10784 13184 10836 13190
rect 10784 13126 10836 13132
rect 10692 13048 10744 13054
rect 10692 12990 10744 12996
rect 10784 12980 10836 12986
rect 10784 12922 10836 12928
rect 10232 12708 10284 12714
rect 10232 12650 10284 12656
rect 9968 12600 10088 12628
rect 10416 12640 10468 12646
rect 7932 12572 7984 12578
rect 7932 12514 7984 12520
rect 7282 11908 7288 11960
rect 7340 11908 7346 11960
rect 6564 11852 6868 11880
rect 6368 11824 6420 11830
rect 6368 11766 6420 11772
rect 6380 11558 6408 11766
rect 6368 11552 6420 11558
rect 6368 11494 6420 11500
rect 6184 11416 6236 11422
rect 6184 11358 6236 11364
rect 6644 11416 6696 11422
rect 6644 11358 6696 11364
rect 6656 10946 6684 11358
rect 6840 11268 6868 11852
rect 7196 11416 7248 11422
rect 7300 11404 7328 11908
rect 7944 11626 7972 12514
rect 8852 12504 8904 12510
rect 8852 12446 8904 12452
rect 8000 12268 8620 12288
rect 8000 12212 8042 12268
rect 8098 12212 8122 12268
rect 8178 12212 8202 12268
rect 8258 12212 8282 12268
rect 8338 12212 8362 12268
rect 8418 12212 8442 12268
rect 8498 12212 8522 12268
rect 8578 12212 8620 12268
rect 8000 12192 8620 12212
rect 8864 12170 8892 12446
rect 8852 12164 8904 12170
rect 9968 12152 9996 12600
rect 10416 12582 10468 12588
rect 10232 12368 10284 12374
rect 10232 12310 10284 12316
rect 9968 12124 10088 12152
rect 8852 12106 8904 12112
rect 10060 11966 10088 12124
rect 10244 11966 10272 12310
rect 10048 11960 10100 11966
rect 10048 11902 10100 11908
rect 10232 11960 10284 11966
rect 10232 11902 10284 11908
rect 9240 11724 9860 11744
rect 9240 11668 9282 11724
rect 9338 11668 9362 11724
rect 9418 11668 9442 11724
rect 9498 11668 9522 11724
rect 9578 11668 9602 11724
rect 9658 11668 9682 11724
rect 9738 11668 9762 11724
rect 9818 11668 9860 11724
rect 9240 11648 9860 11668
rect 7932 11620 7984 11626
rect 7932 11562 7984 11568
rect 8852 11552 8904 11558
rect 8852 11494 8904 11500
rect 7248 11376 7328 11404
rect 7196 11358 7248 11364
rect 6840 11240 6960 11268
rect 6644 10940 6696 10946
rect 6644 10882 6696 10888
rect 6656 10724 6684 10882
rect 6564 10696 6684 10724
rect 6564 10248 6592 10696
rect 6932 10520 6960 11240
rect 7300 10878 7328 11376
rect 8668 11416 8720 11422
rect 8668 11358 8720 11364
rect 8000 11180 8620 11200
rect 8000 11124 8042 11180
rect 8098 11124 8122 11180
rect 8178 11124 8202 11180
rect 8258 11124 8282 11180
rect 8338 11124 8362 11180
rect 8418 11124 8442 11180
rect 8498 11124 8522 11180
rect 8578 11124 8620 11180
rect 8000 11104 8620 11124
rect 7288 10872 7340 10878
rect 7288 10814 7340 10820
rect 6840 10492 6960 10520
rect 6840 10334 6868 10492
rect 6828 10328 6880 10334
rect 6828 10270 6880 10276
rect 6564 10220 6684 10248
rect 6460 9988 6512 9994
rect 6460 9930 6512 9936
rect 6472 9772 6500 9930
rect 6380 9744 6500 9772
rect 6380 8956 6408 9744
rect 6656 9314 6684 10220
rect 6644 9308 6696 9314
rect 6644 9250 6696 9256
rect 6380 8928 6500 8956
rect 6472 8770 6500 8928
rect 6460 8764 6512 8770
rect 6460 8706 6512 8712
rect 6656 8158 6684 9250
rect 7196 9240 7248 9246
rect 7300 9228 7328 10814
rect 8680 10742 8708 11358
rect 8668 10736 8720 10742
rect 8668 10678 8720 10684
rect 8680 10470 8708 10678
rect 8668 10464 8720 10470
rect 8668 10406 8720 10412
rect 8000 10092 8620 10112
rect 8000 10036 8042 10092
rect 8098 10036 8122 10092
rect 8178 10036 8202 10092
rect 8258 10036 8282 10092
rect 8338 10036 8362 10092
rect 8418 10036 8442 10092
rect 8498 10036 8522 10092
rect 8578 10036 8620 10092
rect 8000 10016 8620 10036
rect 8864 9994 8892 11494
rect 9036 11280 9088 11286
rect 9036 11222 9088 11228
rect 9048 10878 9076 11222
rect 10060 10946 10088 11902
rect 10428 11626 10456 12582
rect 10796 12102 10824 12922
rect 10784 12096 10836 12102
rect 10784 12038 10836 12044
rect 10600 11892 10652 11898
rect 10600 11834 10652 11840
rect 10612 11676 10640 11834
rect 10612 11648 10732 11676
rect 10416 11620 10468 11626
rect 10416 11562 10468 11568
rect 10508 11416 10560 11422
rect 10508 11358 10560 11364
rect 10520 10946 10548 11358
rect 10704 11200 10732 11648
rect 11532 11608 11560 13212
rect 11532 11580 11652 11608
rect 11624 11422 11652 11580
rect 11612 11416 11664 11422
rect 11612 11358 11664 11364
rect 10612 11172 10732 11200
rect 10612 11014 10640 11172
rect 11336 11076 11388 11082
rect 11336 11018 11388 11024
rect 10600 11008 10652 11014
rect 10600 10950 10652 10956
rect 10048 10940 10100 10946
rect 10048 10882 10100 10888
rect 10508 10940 10560 10946
rect 10508 10882 10560 10888
rect 9036 10872 9088 10878
rect 9036 10814 9088 10820
rect 9036 10736 9088 10742
rect 9036 10678 9088 10684
rect 9048 10266 9076 10678
rect 9240 10636 9860 10656
rect 9240 10580 9282 10636
rect 9338 10580 9362 10636
rect 9418 10580 9442 10636
rect 9498 10580 9522 10636
rect 9578 10580 9602 10636
rect 9658 10580 9682 10636
rect 9738 10580 9762 10636
rect 9818 10580 9860 10636
rect 9240 10560 9860 10580
rect 9128 10328 9180 10334
rect 10060 10297 10088 10882
rect 10520 10538 10548 10882
rect 10876 10804 10928 10810
rect 10876 10746 10928 10752
rect 10508 10532 10560 10538
rect 10508 10474 10560 10480
rect 9128 10270 9180 10276
rect 10046 10288 10102 10297
rect 9036 10260 9088 10266
rect 9036 10202 9088 10208
rect 8852 9988 8904 9994
rect 8852 9930 8904 9936
rect 8300 9784 8352 9790
rect 8300 9726 8352 9732
rect 8208 9716 8260 9722
rect 8208 9658 8260 9664
rect 7248 9200 7328 9228
rect 7196 9182 7248 9188
rect 6644 8152 6696 8158
rect 6644 8094 6696 8100
rect 7196 8152 7248 8158
rect 7300 8140 7328 9200
rect 8220 9160 8248 9658
rect 8312 9450 8340 9726
rect 8300 9444 8352 9450
rect 8300 9386 8352 9392
rect 9140 9314 9168 10270
rect 10046 10223 10102 10232
rect 10060 9790 10088 10223
rect 10692 9852 10744 9858
rect 10692 9794 10744 9800
rect 10048 9784 10100 9790
rect 10048 9726 10100 9732
rect 9240 9548 9860 9568
rect 9240 9492 9282 9548
rect 9338 9492 9362 9548
rect 9418 9492 9442 9548
rect 9498 9492 9522 9548
rect 9578 9492 9602 9548
rect 9658 9492 9682 9548
rect 9738 9492 9762 9548
rect 9818 9492 9860 9548
rect 9240 9472 9860 9492
rect 9128 9308 9180 9314
rect 9128 9250 9180 9256
rect 8220 9132 8708 9160
rect 8000 9004 8620 9024
rect 8000 8948 8042 9004
rect 8098 8948 8122 9004
rect 8178 8948 8202 9004
rect 8258 8948 8282 9004
rect 8338 8948 8362 9004
rect 8418 8948 8442 9004
rect 8498 8948 8522 9004
rect 8578 8948 8620 9004
rect 8000 8928 8620 8948
rect 7840 8764 7892 8770
rect 7840 8706 7892 8712
rect 7248 8112 7328 8140
rect 7196 8094 7248 8100
rect 6656 7682 6684 8094
rect 7300 7682 7328 8112
rect 6644 7676 6696 7682
rect 6644 7618 6696 7624
rect 7288 7676 7340 7682
rect 7288 7618 7340 7624
rect 5908 7540 5960 7546
rect 5908 7482 5960 7488
rect 6368 7540 6420 7546
rect 6368 7482 6420 7488
rect 6092 7472 6144 7478
rect 6092 7414 6144 7420
rect 6104 7274 6132 7414
rect 6380 7274 6408 7482
rect 6092 7268 6144 7274
rect 6092 7210 6144 7216
rect 6368 7268 6420 7274
rect 6368 7210 6420 7216
rect 6104 6662 6132 7210
rect 6092 6656 6144 6662
rect 6092 6598 6144 6604
rect 6656 6440 6684 7618
rect 6920 7132 6972 7138
rect 7300 7120 7328 7618
rect 6972 7092 7328 7120
rect 6920 7074 6972 7080
rect 7012 6996 7064 7002
rect 7012 6938 7064 6944
rect 6828 6928 6880 6934
rect 6828 6870 6880 6876
rect 6840 6594 6868 6870
rect 6828 6588 6880 6594
rect 6828 6530 6880 6536
rect 6656 6412 6776 6440
rect 6552 6384 6604 6390
rect 6552 6326 6604 6332
rect 6564 6050 6592 6326
rect 6552 6044 6604 6050
rect 6552 5986 6604 5992
rect 6748 5982 6776 6412
rect 7024 6186 7052 6938
rect 7300 6637 7328 7092
rect 7472 6928 7524 6934
rect 7472 6870 7524 6876
rect 7286 6628 7342 6637
rect 7286 6563 7342 6572
rect 7484 6526 7512 6870
rect 7852 6662 7880 8706
rect 8680 8566 8708 9132
rect 8852 8900 8904 8906
rect 8852 8842 8904 8848
rect 8300 8560 8352 8566
rect 8300 8502 8352 8508
rect 8668 8560 8720 8566
rect 8668 8502 8720 8508
rect 8312 8362 8340 8502
rect 8300 8356 8352 8362
rect 8300 8298 8352 8304
rect 8000 7916 8620 7936
rect 8000 7860 8042 7916
rect 8098 7860 8122 7916
rect 8178 7860 8202 7916
rect 8258 7860 8282 7916
rect 8338 7860 8362 7916
rect 8418 7860 8442 7916
rect 8498 7860 8522 7916
rect 8578 7860 8620 7916
rect 8000 7840 8620 7860
rect 8864 7614 8892 8842
rect 9140 8158 9168 9250
rect 9240 8460 9860 8480
rect 9240 8404 9282 8460
rect 9338 8404 9362 8460
rect 9418 8404 9442 8460
rect 9498 8404 9522 8460
rect 9578 8404 9602 8460
rect 9658 8404 9682 8460
rect 9738 8404 9762 8460
rect 9818 8404 9860 8460
rect 9240 8384 9860 8404
rect 9128 8152 9180 8158
rect 9128 8094 9180 8100
rect 9140 7735 9168 8094
rect 9404 8084 9456 8090
rect 9404 8026 9456 8032
rect 9416 7818 9444 8026
rect 10060 7818 10088 9726
rect 10324 9648 10376 9654
rect 10324 9590 10376 9596
rect 10336 9382 10364 9590
rect 10704 9450 10732 9794
rect 10888 9722 10916 10746
rect 11348 10470 11376 11018
rect 11336 10464 11388 10470
rect 11336 10406 11388 10412
rect 11624 10402 11652 11358
rect 11808 11336 11836 13942
rect 12360 13054 12388 14078
rect 12544 13666 12572 15252
rect 12624 15234 12676 15240
rect 13188 15230 13216 18108
rect 13268 18090 13320 18096
rect 14292 17882 14320 18924
rect 14568 18494 14596 18924
rect 14844 18630 14872 19110
rect 16132 19106 16160 19604
rect 16856 19586 16908 19592
rect 16868 19203 16896 19586
rect 16854 19194 16910 19203
rect 16854 19129 16910 19138
rect 16120 19100 16172 19106
rect 16120 19042 16172 19048
rect 16132 18630 16160 19042
rect 17144 19038 17172 20470
rect 17696 19650 17724 20470
rect 17868 19984 17920 19990
rect 17868 19926 17920 19932
rect 17684 19644 17736 19650
rect 17684 19586 17736 19592
rect 17880 19582 17908 19926
rect 17868 19576 17920 19582
rect 17868 19518 17920 19524
rect 17592 19440 17644 19446
rect 17592 19382 17644 19388
rect 17604 19242 17632 19382
rect 17592 19236 17644 19242
rect 17592 19178 17644 19184
rect 17880 19038 17908 19518
rect 17132 19032 17184 19038
rect 17132 18974 17184 18980
rect 17316 19032 17368 19038
rect 17316 18974 17368 18980
rect 17868 19032 17920 19038
rect 17868 18974 17920 18980
rect 14832 18624 14884 18630
rect 14832 18566 14884 18572
rect 16120 18624 16172 18630
rect 16120 18566 16172 18572
rect 15568 18556 15620 18562
rect 15568 18498 15620 18504
rect 14556 18488 14608 18494
rect 14556 18430 14608 18436
rect 14568 18272 14596 18430
rect 14568 18244 14688 18272
rect 14280 17876 14332 17882
rect 14280 17818 14332 17824
rect 14464 17876 14516 17882
rect 14464 17818 14516 17824
rect 13360 17808 13412 17814
rect 13360 17750 13412 17756
rect 13372 17338 13400 17750
rect 13600 17708 14220 17728
rect 13600 17652 13642 17708
rect 13698 17652 13722 17708
rect 13778 17652 13802 17708
rect 13858 17652 13882 17708
rect 13938 17652 13962 17708
rect 14018 17652 14042 17708
rect 14098 17652 14122 17708
rect 14178 17652 14220 17708
rect 13600 17632 14220 17652
rect 14096 17536 14148 17542
rect 14096 17478 14148 17484
rect 14278 17486 14334 17495
rect 13360 17332 13412 17338
rect 13360 17274 13412 17280
rect 14108 16862 14136 17478
rect 14476 17474 14504 17818
rect 14278 17421 14334 17430
rect 14464 17468 14516 17474
rect 14292 16930 14320 17421
rect 14464 17410 14516 17416
rect 14280 16924 14332 16930
rect 14280 16866 14332 16872
rect 14476 16862 14504 17410
rect 14660 16862 14688 18244
rect 14840 18252 15460 18272
rect 14840 18196 14882 18252
rect 14938 18196 14962 18252
rect 15018 18196 15042 18252
rect 15098 18196 15122 18252
rect 15178 18196 15202 18252
rect 15258 18196 15282 18252
rect 15338 18196 15362 18252
rect 15418 18196 15460 18252
rect 14840 18176 15460 18196
rect 15580 17950 15608 18498
rect 17328 18494 17356 18974
rect 18616 18902 18644 21236
rect 19616 21218 19668 21224
rect 18880 21072 18932 21078
rect 18880 21014 18932 21020
rect 18892 20806 18920 21014
rect 19200 20972 19820 20992
rect 19200 20916 19242 20972
rect 19298 20916 19322 20972
rect 19378 20916 19402 20972
rect 19458 20916 19482 20972
rect 19538 20916 19562 20972
rect 19618 20916 19642 20972
rect 19698 20916 19722 20972
rect 19778 20916 19820 20972
rect 19200 20896 19820 20916
rect 19904 20806 19932 21558
rect 19996 21418 20024 21558
rect 19984 21412 20036 21418
rect 20364 21400 20392 21694
rect 20440 21516 21060 21536
rect 20440 21460 20482 21516
rect 20538 21460 20562 21516
rect 20618 21460 20642 21516
rect 20698 21460 20722 21516
rect 20778 21460 20802 21516
rect 20858 21460 20882 21516
rect 20938 21460 20962 21516
rect 21018 21460 21060 21516
rect 20440 21440 21060 21460
rect 20364 21372 20484 21400
rect 19984 21354 20036 21360
rect 20076 21208 20128 21214
rect 20076 21150 20128 21156
rect 18880 20800 18932 20806
rect 18880 20742 18932 20748
rect 19892 20800 19944 20806
rect 19892 20742 19944 20748
rect 20088 20670 20116 21150
rect 20456 20874 20484 21372
rect 20444 20868 20496 20874
rect 20444 20810 20496 20816
rect 19156 20664 19208 20670
rect 19156 20606 19208 20612
rect 20076 20664 20128 20670
rect 20076 20606 20128 20612
rect 19168 20179 19196 20606
rect 20088 20179 20116 20606
rect 20456 20584 20484 20810
rect 20364 20556 20484 20584
rect 19154 20170 19210 20179
rect 19154 20105 19210 20114
rect 20074 20170 20130 20179
rect 20074 20105 20076 20114
rect 20128 20105 20130 20114
rect 20364 20108 20392 20556
rect 20440 20428 21060 20448
rect 20440 20372 20482 20428
rect 20538 20372 20562 20428
rect 20618 20372 20642 20428
rect 20698 20372 20722 20428
rect 20778 20372 20802 20428
rect 20858 20372 20882 20428
rect 20938 20372 20962 20428
rect 21018 20372 21060 20428
rect 20440 20352 21060 20372
rect 20364 20080 20484 20108
rect 20076 20062 20128 20068
rect 18880 20052 18932 20058
rect 18880 19994 18932 20000
rect 18892 19786 18920 19994
rect 20168 19984 20220 19990
rect 20168 19926 20220 19932
rect 19200 19884 19820 19904
rect 19200 19828 19242 19884
rect 19298 19828 19322 19884
rect 19378 19828 19402 19884
rect 19458 19828 19482 19884
rect 19538 19828 19562 19884
rect 19618 19828 19642 19884
rect 19698 19828 19722 19884
rect 19778 19828 19820 19884
rect 19200 19808 19820 19828
rect 18880 19780 18932 19786
rect 20180 19768 20208 19926
rect 18880 19722 18932 19728
rect 20088 19740 20208 19768
rect 19062 19682 19118 19691
rect 19062 19617 19118 19626
rect 19076 19496 19104 19617
rect 18984 19468 19104 19496
rect 18984 19020 19012 19468
rect 19248 19440 19300 19446
rect 19248 19382 19300 19388
rect 19260 19174 19288 19382
rect 20088 19292 20116 19740
rect 20456 19496 20484 20080
rect 20364 19468 20484 19496
rect 20088 19264 20208 19292
rect 19248 19168 19300 19174
rect 19248 19110 19300 19116
rect 20180 19106 20208 19264
rect 20168 19100 20220 19106
rect 20168 19042 20220 19048
rect 18984 18992 19104 19020
rect 17776 18896 17828 18902
rect 17776 18838 17828 18844
rect 18604 18896 18656 18902
rect 18604 18838 18656 18844
rect 17788 18630 17816 18838
rect 17592 18624 17644 18630
rect 17592 18566 17644 18572
rect 17776 18624 17828 18630
rect 17776 18566 17828 18572
rect 17316 18488 17368 18494
rect 17316 18430 17368 18436
rect 17604 18408 17632 18566
rect 17868 18556 17920 18562
rect 17868 18498 17920 18504
rect 17684 18488 17736 18494
rect 17684 18430 17736 18436
rect 17512 18380 17632 18408
rect 15752 18352 15804 18358
rect 15752 18294 15804 18300
rect 15764 17950 15792 18294
rect 16488 18080 16540 18086
rect 16488 18022 16540 18028
rect 15568 17944 15620 17950
rect 15568 17886 15620 17892
rect 15752 17944 15804 17950
rect 15752 17886 15804 17892
rect 15844 17944 15896 17950
rect 15844 17886 15896 17892
rect 16028 17944 16080 17950
rect 16028 17886 16080 17892
rect 14832 17808 14884 17814
rect 14832 17750 14884 17756
rect 14844 17495 14872 17750
rect 14830 17486 14886 17495
rect 14830 17421 14886 17430
rect 15580 17456 15608 17886
rect 15660 17468 15712 17474
rect 15580 17428 15660 17456
rect 14740 17264 14792 17270
rect 14740 17206 14792 17212
rect 14752 17048 14780 17206
rect 14840 17164 15460 17184
rect 14840 17108 14882 17164
rect 14938 17108 14962 17164
rect 15018 17108 15042 17164
rect 15098 17108 15122 17164
rect 15178 17108 15202 17164
rect 15258 17108 15282 17164
rect 15338 17108 15362 17164
rect 15418 17108 15460 17164
rect 14840 17088 15460 17108
rect 14752 17020 14872 17048
rect 13268 16856 13320 16862
rect 13268 16798 13320 16804
rect 14096 16856 14148 16862
rect 14096 16798 14148 16804
rect 14464 16856 14516 16862
rect 14464 16798 14516 16804
rect 14648 16856 14700 16862
rect 14648 16798 14700 16804
rect 13280 16522 13308 16798
rect 13600 16620 14220 16640
rect 13600 16564 13642 16620
rect 13698 16564 13722 16620
rect 13778 16564 13802 16620
rect 13858 16564 13882 16620
rect 13938 16564 13962 16620
rect 14018 16564 14042 16620
rect 14098 16564 14122 16620
rect 14178 16564 14220 16620
rect 13600 16544 14220 16564
rect 13268 16516 13320 16522
rect 13268 16458 13320 16464
rect 13360 16380 13412 16386
rect 13360 16322 13412 16328
rect 13372 16164 13400 16322
rect 13372 16136 13492 16164
rect 13464 15688 13492 16136
rect 14476 15774 14504 16798
rect 14844 16454 14872 17020
rect 15286 17008 15292 17060
rect 15344 17008 15350 17060
rect 15304 16776 15332 17008
rect 15580 16862 15608 17428
rect 15660 17410 15712 17416
rect 15856 17270 15884 17886
rect 15844 17264 15896 17270
rect 15844 17206 15896 17212
rect 15568 16856 15620 16862
rect 15568 16798 15620 16804
rect 15304 16748 15424 16776
rect 15396 16454 15424 16748
rect 15580 16504 15608 16798
rect 15752 16516 15804 16522
rect 15580 16476 15752 16504
rect 14832 16448 14884 16454
rect 14832 16390 14884 16396
rect 15384 16448 15436 16454
rect 15384 16390 15436 16396
rect 14840 16076 15460 16096
rect 14840 16020 14882 16076
rect 14938 16020 14962 16076
rect 15018 16020 15042 16076
rect 15098 16020 15122 16076
rect 15178 16020 15202 16076
rect 15258 16020 15282 16076
rect 15338 16020 15362 16076
rect 15418 16020 15460 16076
rect 14840 16000 15460 16020
rect 15580 15892 15608 16476
rect 16040 16504 16068 17886
rect 16304 17876 16356 17882
rect 16500 17864 16528 18022
rect 17316 17944 17368 17950
rect 17316 17886 17368 17892
rect 16500 17836 16620 17864
rect 16304 17818 16356 17824
rect 16316 17066 16344 17818
rect 16304 17060 16356 17066
rect 16304 17002 16356 17008
rect 16592 16980 16620 17836
rect 17132 17400 17184 17406
rect 17132 17342 17184 17348
rect 16856 17264 16908 17270
rect 16856 17206 16908 17212
rect 15752 16458 15804 16464
rect 15856 16476 16068 16504
rect 16500 16952 16620 16980
rect 15856 15960 15884 16476
rect 15936 16380 15988 16386
rect 15988 16340 16252 16368
rect 15936 16322 15988 16328
rect 15856 15932 15976 15960
rect 15488 15864 15608 15892
rect 15750 15900 15806 15909
rect 14464 15768 14516 15774
rect 14464 15710 14516 15716
rect 13372 15660 13492 15688
rect 13176 15224 13228 15230
rect 13176 15166 13228 15172
rect 12808 15088 12860 15094
rect 12808 15030 12860 15036
rect 12820 14210 12848 15030
rect 13188 15008 13216 15166
rect 13096 14980 13216 15008
rect 12808 14204 12860 14210
rect 12808 14146 12860 14152
rect 12532 13660 12584 13666
rect 12532 13602 12584 13608
rect 12716 13660 12768 13666
rect 13096 13648 13124 14980
rect 13372 14686 13400 15660
rect 14280 15632 14332 15638
rect 14280 15574 14332 15580
rect 13600 15532 14220 15552
rect 13600 15476 13642 15532
rect 13698 15476 13722 15532
rect 13778 15476 13802 15532
rect 13858 15476 13882 15532
rect 13938 15476 13962 15532
rect 14018 15476 14042 15532
rect 14098 15476 14122 15532
rect 14178 15476 14220 15532
rect 13600 15456 14220 15476
rect 14292 15348 14320 15574
rect 14200 15320 14320 15348
rect 13360 14680 13412 14686
rect 13360 14622 13412 14628
rect 13096 13620 13216 13648
rect 12716 13602 12768 13608
rect 12544 13258 12572 13602
rect 12532 13252 12584 13258
rect 12532 13194 12584 13200
rect 12728 13190 12756 13602
rect 12992 13456 13044 13462
rect 12992 13398 13044 13404
rect 12716 13184 12768 13190
rect 12716 13126 12768 13132
rect 11980 13048 12032 13054
rect 11980 12990 12032 12996
rect 12348 13048 12400 13054
rect 12348 12990 12400 12996
rect 11992 12714 12020 12990
rect 11980 12708 12032 12714
rect 11980 12650 12032 12656
rect 12360 12615 12388 12990
rect 12346 12606 12402 12615
rect 12346 12541 12402 12550
rect 11980 11960 12032 11966
rect 11980 11902 12032 11908
rect 11992 11558 12020 11902
rect 11980 11552 12032 11558
rect 11980 11494 12032 11500
rect 12360 11422 12388 12541
rect 13004 12510 13032 13398
rect 13188 13104 13216 13620
rect 13372 13598 13400 14622
rect 14200 14600 14228 15320
rect 14476 15162 14504 15710
rect 15488 15416 15516 15864
rect 15750 15835 15806 15844
rect 15488 15388 15608 15416
rect 14740 15292 14792 15298
rect 14740 15234 14792 15240
rect 15580 15280 15608 15388
rect 15660 15292 15712 15298
rect 15580 15252 15660 15280
rect 14464 15156 14516 15162
rect 14464 15098 14516 15104
rect 14476 14686 14504 15098
rect 14464 14680 14516 14686
rect 14464 14622 14516 14628
rect 14200 14572 14320 14600
rect 13452 14544 13504 14550
rect 13452 14486 13504 14492
rect 13464 14278 13492 14486
rect 13600 14444 14220 14464
rect 13600 14388 13642 14444
rect 13698 14388 13722 14444
rect 13778 14388 13802 14444
rect 13858 14388 13882 14444
rect 13938 14388 13962 14444
rect 14018 14388 14042 14444
rect 14098 14388 14122 14444
rect 14178 14388 14220 14444
rect 13600 14368 14220 14388
rect 14292 14278 14320 14572
rect 14556 14544 14608 14550
rect 14556 14486 14608 14492
rect 14568 14346 14596 14486
rect 14556 14340 14608 14346
rect 14556 14282 14608 14288
rect 13452 14272 13504 14278
rect 13452 14214 13504 14220
rect 14280 14272 14332 14278
rect 14280 14214 14332 14220
rect 14372 14204 14424 14210
rect 14372 14146 14424 14152
rect 14556 14204 14608 14210
rect 14752 14201 14780 15234
rect 14840 14988 15460 15008
rect 14840 14932 14882 14988
rect 14938 14932 14962 14988
rect 15018 14932 15042 14988
rect 15098 14932 15122 14988
rect 15178 14932 15202 14988
rect 15258 14932 15282 14988
rect 15338 14932 15362 14988
rect 15418 14932 15460 14988
rect 14840 14912 15460 14932
rect 15200 14612 15252 14618
rect 15200 14554 15252 14560
rect 15212 14210 15240 14554
rect 15200 14204 15252 14210
rect 14556 14146 14608 14152
rect 14738 14192 14794 14201
rect 14384 13802 14412 14146
rect 14372 13796 14424 13802
rect 14372 13738 14424 13744
rect 14568 13713 14596 14146
rect 15200 14146 15252 14152
rect 15580 14142 15608 15252
rect 15660 15234 15712 15240
rect 15764 14210 15792 15835
rect 15948 15094 15976 15932
rect 16028 15224 16080 15230
rect 16028 15166 16080 15172
rect 15936 15088 15988 15094
rect 15936 15030 15988 15036
rect 15844 14544 15896 14550
rect 15844 14486 15896 14492
rect 15752 14204 15804 14210
rect 15750 14192 15752 14201
rect 15804 14192 15806 14201
rect 14738 14127 14794 14136
rect 15568 14136 15620 14142
rect 14554 13704 14610 13713
rect 14554 13639 14610 13648
rect 13360 13592 13412 13598
rect 13360 13534 13412 13540
rect 13452 13456 13504 13462
rect 13452 13398 13504 13404
rect 13464 13190 13492 13398
rect 13600 13356 14220 13376
rect 13600 13300 13642 13356
rect 13698 13300 13722 13356
rect 13778 13300 13802 13356
rect 13858 13300 13882 13356
rect 13938 13300 13962 13356
rect 14018 13300 14042 13356
rect 14098 13300 14122 13356
rect 14178 13300 14220 13356
rect 13600 13280 14220 13300
rect 13452 13184 13504 13190
rect 13452 13126 13504 13132
rect 14556 13184 14608 13190
rect 14556 13126 14608 13132
rect 13360 13116 13412 13122
rect 13188 13076 13360 13104
rect 13360 13058 13412 13064
rect 14568 12968 14596 13126
rect 14476 12940 14596 12968
rect 13266 12606 13322 12615
rect 13266 12541 13268 12550
rect 13320 12541 13322 12550
rect 13268 12514 13320 12520
rect 12992 12504 13044 12510
rect 12992 12446 13044 12452
rect 13452 12504 13504 12510
rect 13452 12446 13504 12452
rect 13268 12096 13320 12102
rect 13268 12038 13320 12044
rect 13280 11626 13308 12038
rect 13464 12034 13492 12446
rect 14476 12356 14504 12940
rect 14476 12328 14596 12356
rect 13600 12268 14220 12288
rect 13600 12212 13642 12268
rect 13698 12212 13722 12268
rect 13778 12212 13802 12268
rect 13858 12212 13882 12268
rect 13938 12212 13962 12268
rect 14018 12212 14042 12268
rect 14098 12212 14122 12268
rect 14178 12212 14220 12268
rect 13600 12192 14220 12212
rect 14568 12170 14596 12328
rect 14556 12164 14608 12170
rect 14556 12106 14608 12112
rect 13452 12028 13504 12034
rect 13452 11970 13504 11976
rect 14002 11996 14058 12005
rect 13268 11620 13320 11626
rect 13268 11562 13320 11568
rect 12348 11416 12400 11422
rect 12348 11358 12400 11364
rect 11808 11308 11928 11336
rect 11612 10396 11664 10402
rect 11612 10338 11664 10344
rect 11336 9784 11388 9790
rect 11336 9726 11388 9732
rect 10876 9716 10928 9722
rect 10876 9658 10928 9664
rect 11060 9716 11112 9722
rect 11060 9658 11112 9664
rect 10692 9444 10744 9450
rect 10692 9386 10744 9392
rect 10324 9376 10376 9382
rect 10324 9318 10376 9324
rect 11072 8906 11100 9658
rect 11348 9450 11376 9726
rect 11624 9450 11652 10338
rect 11336 9444 11388 9450
rect 11336 9386 11388 9392
rect 11612 9444 11664 9450
rect 11612 9386 11664 9392
rect 11900 9296 11928 11308
rect 12360 10334 12388 11358
rect 13464 10946 13492 11970
rect 14002 11931 14058 11940
rect 14016 11490 14044 11931
rect 14004 11484 14056 11490
rect 14004 11426 14056 11432
rect 14556 11416 14608 11422
rect 14556 11358 14608 11364
rect 13600 11180 14220 11200
rect 13600 11124 13642 11180
rect 13698 11124 13722 11180
rect 13778 11124 13802 11180
rect 13858 11124 13882 11180
rect 13938 11124 13962 11180
rect 14018 11124 14042 11180
rect 14098 11124 14122 11180
rect 14178 11124 14220 11180
rect 13600 11104 14220 11124
rect 13452 10940 13504 10946
rect 13452 10882 13504 10888
rect 13268 10872 13320 10878
rect 13268 10814 13320 10820
rect 13280 10538 13308 10814
rect 13268 10532 13320 10538
rect 13268 10474 13320 10480
rect 12348 10328 12400 10334
rect 12348 10270 12400 10276
rect 13268 10328 13320 10334
rect 13268 10270 13320 10276
rect 12360 9790 12388 10270
rect 12624 9852 12676 9858
rect 12624 9794 12676 9800
rect 12348 9784 12400 9790
rect 12348 9726 12400 9732
rect 11808 9268 11928 9296
rect 11060 8900 11112 8906
rect 11060 8842 11112 8848
rect 10692 8764 10744 8770
rect 10692 8706 10744 8712
rect 10416 8628 10468 8634
rect 10416 8570 10468 8576
rect 9404 7812 9456 7818
rect 9404 7754 9456 7760
rect 10048 7812 10100 7818
rect 10048 7754 10100 7760
rect 9126 7726 9182 7735
rect 9126 7661 9182 7670
rect 10060 7614 10088 7754
rect 8852 7608 8904 7614
rect 8852 7550 8904 7556
rect 10048 7608 10100 7614
rect 10048 7550 10100 7556
rect 9128 7472 9180 7478
rect 9128 7414 9180 7420
rect 8000 6828 8620 6848
rect 8000 6772 8042 6828
rect 8098 6772 8122 6828
rect 8178 6772 8202 6828
rect 8258 6772 8282 6828
rect 8338 6772 8362 6828
rect 8418 6772 8442 6828
rect 8498 6772 8522 6828
rect 8578 6772 8620 6828
rect 8000 6752 8620 6772
rect 7656 6656 7708 6662
rect 7656 6598 7708 6604
rect 7840 6656 7892 6662
rect 7840 6598 7892 6604
rect 7472 6520 7524 6526
rect 7472 6462 7524 6468
rect 7012 6180 7064 6186
rect 7012 6122 7064 6128
rect 7668 6050 7696 6598
rect 7852 6526 7880 6598
rect 8484 6588 8536 6594
rect 8484 6530 8536 6536
rect 7840 6520 7892 6526
rect 7840 6462 7892 6468
rect 8208 6520 8260 6526
rect 8208 6462 8260 6468
rect 8220 6393 8248 6462
rect 8496 6440 8524 6530
rect 8404 6412 8524 6440
rect 7748 6384 7800 6390
rect 7748 6326 7800 6332
rect 8206 6384 8262 6393
rect 7760 6186 7788 6326
rect 8206 6319 8262 6328
rect 8404 6186 8432 6412
rect 9140 6186 9168 7414
rect 9240 7372 9860 7392
rect 9240 7316 9282 7372
rect 9338 7316 9362 7372
rect 9418 7316 9442 7372
rect 9498 7316 9522 7372
rect 9578 7316 9602 7372
rect 9658 7316 9682 7372
rect 9738 7316 9762 7372
rect 9818 7316 9860 7372
rect 9240 7296 9860 7316
rect 9306 7012 9312 7064
rect 9364 7012 9370 7064
rect 9306 6994 9370 7012
rect 9306 6938 9310 6994
rect 9366 6938 9370 6994
rect 10232 6996 10284 7002
rect 10232 6938 10284 6944
rect 9306 6929 9370 6938
rect 10244 6637 10272 6938
rect 10428 6662 10456 8570
rect 10704 8362 10732 8706
rect 10692 8356 10744 8362
rect 10692 8298 10744 8304
rect 10692 8220 10744 8226
rect 10692 8162 10744 8168
rect 10704 7735 10732 8162
rect 11808 8158 11836 9268
rect 12360 9160 12388 9726
rect 12440 9172 12492 9178
rect 12360 9132 12440 9160
rect 11796 8152 11848 8158
rect 11796 8094 11848 8100
rect 11336 8084 11388 8090
rect 11336 8026 11388 8032
rect 11348 7818 11376 8026
rect 11980 8016 12032 8022
rect 11980 7958 12032 7964
rect 11336 7812 11388 7818
rect 11336 7754 11388 7760
rect 10690 7726 10746 7735
rect 10690 7661 10746 7670
rect 10876 7676 10928 7682
rect 10876 7618 10928 7624
rect 10416 6656 10468 6662
rect 10230 6628 10286 6637
rect 10416 6598 10468 6604
rect 10230 6563 10286 6572
rect 10324 6520 10376 6526
rect 10324 6462 10376 6468
rect 9956 6384 10008 6390
rect 9956 6326 10008 6332
rect 9240 6284 9860 6304
rect 9240 6228 9282 6284
rect 9338 6228 9362 6284
rect 9418 6228 9442 6284
rect 9498 6228 9522 6284
rect 9578 6228 9602 6284
rect 9658 6228 9682 6284
rect 9738 6228 9762 6284
rect 9818 6228 9860 6284
rect 9240 6208 9860 6228
rect 7748 6180 7800 6186
rect 7748 6122 7800 6128
rect 8392 6180 8444 6186
rect 8392 6122 8444 6128
rect 9128 6180 9180 6186
rect 9968 6168 9996 6326
rect 10336 6186 10364 6462
rect 9128 6122 9180 6128
rect 9600 6140 9996 6168
rect 10324 6180 10376 6186
rect 7656 6044 7708 6050
rect 7656 5986 7708 5992
rect 6736 5976 6788 5982
rect 6736 5918 6788 5924
rect 8000 5740 8620 5760
rect 8000 5684 8042 5740
rect 8098 5684 8122 5740
rect 8178 5684 8202 5740
rect 8258 5684 8282 5740
rect 8338 5684 8362 5740
rect 8418 5684 8442 5740
rect 8498 5684 8522 5740
rect 8578 5684 8620 5740
rect 8000 5664 8620 5684
rect 20 196 72 202
rect 20 138 72 144
rect 32 0 60 138
rect 9600 0 9628 6140
rect 10324 6122 10376 6128
rect 10888 4214 10916 7618
rect 11612 7540 11664 7546
rect 11612 7482 11664 7488
rect 11244 6996 11296 7002
rect 11244 6938 11296 6944
rect 11256 6458 11284 6938
rect 11624 6730 11652 7482
rect 11992 7324 12020 7958
rect 12360 7735 12388 9132
rect 12440 9114 12492 9120
rect 12636 8906 12664 9794
rect 12992 9648 13044 9654
rect 12992 9590 13044 9596
rect 13004 9382 13032 9590
rect 12992 9376 13044 9382
rect 12992 9318 13044 9324
rect 13084 9308 13136 9314
rect 13084 9250 13136 9256
rect 12624 8900 12676 8906
rect 12624 8842 12676 8848
rect 13096 8702 13124 9250
rect 13280 8906 13308 10270
rect 13464 9308 13492 10882
rect 14464 10736 14516 10742
rect 14464 10678 14516 10684
rect 14476 10334 14504 10678
rect 14568 10538 14596 11358
rect 14556 10532 14608 10538
rect 14556 10474 14608 10480
rect 14188 10328 14240 10334
rect 14464 10328 14516 10334
rect 14240 10288 14320 10316
rect 14188 10270 14240 10276
rect 13600 10092 14220 10112
rect 13600 10036 13642 10092
rect 13698 10036 13722 10092
rect 13778 10036 13802 10092
rect 13858 10036 13882 10092
rect 13938 10036 13962 10092
rect 14018 10036 14042 10092
rect 14098 10036 14122 10092
rect 14178 10036 14220 10092
rect 13600 10016 14220 10036
rect 14292 9790 14320 10288
rect 14464 10270 14516 10276
rect 14556 10192 14608 10198
rect 14556 10134 14608 10140
rect 14280 9784 14332 9790
rect 14280 9726 14332 9732
rect 14280 9648 14332 9654
rect 14280 9590 14332 9596
rect 13446 9256 13452 9308
rect 13504 9256 13510 9308
rect 13268 8900 13320 8906
rect 13268 8842 13320 8848
rect 13464 8833 13492 9256
rect 13600 9004 14220 9024
rect 13600 8948 13642 9004
rect 13698 8948 13722 9004
rect 13778 8948 13802 9004
rect 13858 8948 13882 9004
rect 13938 8948 13962 9004
rect 14018 8948 14042 9004
rect 14098 8948 14122 9004
rect 14178 8948 14220 9004
rect 13600 8928 14220 8948
rect 14292 8838 14320 9590
rect 14568 9450 14596 10134
rect 14556 9444 14608 9450
rect 14556 9386 14608 9392
rect 13450 8824 13506 8833
rect 13268 8764 13320 8770
rect 14280 8832 14332 8838
rect 14280 8774 14332 8780
rect 13450 8764 13506 8768
rect 13450 8759 13452 8764
rect 13268 8706 13320 8712
rect 13504 8759 13506 8764
rect 13452 8706 13504 8712
rect 13084 8696 13136 8702
rect 13084 8638 13136 8644
rect 13096 8480 13124 8638
rect 13004 8452 13124 8480
rect 13004 7868 13032 8452
rect 13280 8362 13308 8706
rect 13268 8356 13320 8362
rect 13268 8298 13320 8304
rect 13004 7840 13124 7868
rect 12346 7726 12402 7735
rect 12346 7661 12402 7670
rect 12900 7676 12952 7682
rect 12360 7614 12388 7661
rect 13096 7664 13124 7840
rect 13280 7750 13308 8298
rect 14280 8152 14332 8158
rect 14280 8094 14332 8100
rect 13452 8016 13504 8022
rect 13452 7958 13504 7964
rect 13268 7744 13320 7750
rect 13268 7686 13320 7692
rect 13096 7636 13216 7664
rect 12900 7618 12952 7624
rect 12348 7608 12400 7614
rect 12348 7550 12400 7556
rect 11900 7296 12020 7324
rect 11900 6780 11928 7296
rect 12164 7200 12216 7206
rect 12164 7142 12216 7148
rect 11900 6752 12020 6780
rect 11612 6724 11664 6730
rect 11612 6666 11664 6672
rect 11992 6594 12020 6752
rect 11980 6588 12032 6594
rect 12176 6576 12204 7142
rect 12360 6594 12388 7550
rect 12532 7472 12584 7478
rect 12912 7460 12940 7618
rect 12532 7414 12584 7420
rect 12820 7432 12940 7460
rect 13084 7472 13136 7478
rect 12544 7138 12572 7414
rect 12532 7132 12584 7138
rect 12532 7074 12584 7080
rect 12820 6916 12848 7432
rect 13084 7414 13136 7420
rect 13096 7070 13124 7414
rect 13188 7274 13216 7636
rect 13176 7268 13228 7274
rect 13176 7210 13228 7216
rect 13084 7064 13136 7070
rect 13084 7006 13136 7012
rect 13268 6928 13320 6934
rect 12820 6888 12940 6916
rect 12348 6588 12400 6594
rect 12176 6548 12296 6576
rect 11980 6530 12032 6536
rect 11244 6452 11296 6458
rect 11244 6394 11296 6400
rect 12268 6186 12296 6548
rect 12348 6530 12400 6536
rect 12256 6180 12308 6186
rect 12256 6122 12308 6128
rect 12268 6027 12296 6122
rect 12254 6018 12310 6027
rect 12912 5982 12940 6888
rect 13268 6870 13320 6876
rect 13280 6730 13308 6870
rect 13268 6724 13320 6730
rect 13268 6666 13320 6672
rect 13266 6018 13322 6027
rect 12254 5953 12310 5962
rect 12900 5976 12952 5982
rect 13266 5953 13268 5962
rect 12900 5918 12952 5924
rect 13320 5953 13322 5962
rect 13268 5918 13320 5924
rect 10876 4208 10928 4214
rect 10876 4150 10928 4156
rect 13464 202 13492 7958
rect 13600 7916 14220 7936
rect 13600 7860 13642 7916
rect 13698 7860 13722 7916
rect 13778 7860 13802 7916
rect 13858 7860 13882 7916
rect 13938 7860 13962 7916
rect 14018 7860 14042 7916
rect 14098 7860 14122 7916
rect 14178 7860 14220 7916
rect 13600 7840 14220 7860
rect 13634 7726 13690 7735
rect 13634 7661 13690 7670
rect 14004 7676 14056 7682
rect 13648 7070 13676 7661
rect 14004 7618 14056 7624
rect 13636 7064 13688 7070
rect 13636 7006 13688 7012
rect 14016 7002 14044 7618
rect 14004 6996 14056 7002
rect 14004 6938 14056 6944
rect 13600 6828 14220 6848
rect 13600 6772 13642 6828
rect 13698 6772 13722 6828
rect 13778 6772 13802 6828
rect 13858 6772 13882 6828
rect 13938 6772 13962 6828
rect 14018 6772 14042 6828
rect 14098 6772 14122 6828
rect 14178 6772 14220 6828
rect 13600 6752 14220 6772
rect 13820 6656 13872 6662
rect 13820 6598 13872 6604
rect 13832 6186 13860 6598
rect 13820 6180 13872 6186
rect 13820 6122 13872 6128
rect 14292 6050 14320 8094
rect 14752 8072 14780 14127
rect 15750 14127 15806 14136
rect 15568 14078 15620 14084
rect 15476 14068 15528 14074
rect 15476 14010 15528 14016
rect 14840 13900 15460 13920
rect 14840 13844 14882 13900
rect 14938 13844 14962 13900
rect 15018 13844 15042 13900
rect 15098 13844 15122 13900
rect 15178 13844 15202 13900
rect 15258 13844 15282 13900
rect 15338 13844 15362 13900
rect 15418 13844 15460 13900
rect 14840 13824 15460 13844
rect 15290 13704 15346 13713
rect 15290 13639 15346 13648
rect 15304 13122 15332 13639
rect 15488 13225 15516 14010
rect 15474 13216 15530 13225
rect 15474 13151 15530 13160
rect 15292 13116 15344 13122
rect 15292 13058 15344 13064
rect 15304 12981 15332 13058
rect 15290 12972 15346 12981
rect 15290 12907 15346 12916
rect 14840 12812 15460 12832
rect 14840 12756 14882 12812
rect 14938 12756 14962 12812
rect 15018 12756 15042 12812
rect 15098 12756 15122 12812
rect 15178 12756 15202 12812
rect 15258 12756 15282 12812
rect 15338 12756 15362 12812
rect 15418 12756 15460 12812
rect 14840 12736 15460 12756
rect 15488 12034 15516 13151
rect 15568 13116 15620 13122
rect 15568 13058 15620 13064
rect 15580 12510 15608 13058
rect 15660 12912 15712 12918
rect 15660 12854 15712 12860
rect 15568 12504 15620 12510
rect 15568 12446 15620 12452
rect 15580 12034 15608 12446
rect 15672 12102 15700 12854
rect 15856 12578 15884 14486
rect 16040 13252 16068 15166
rect 16224 14689 16252 16340
rect 16304 15088 16356 15094
rect 16304 15030 16356 15036
rect 16210 14680 16266 14689
rect 16210 14615 16266 14624
rect 16022 13200 16028 13252
rect 16080 13200 16086 13252
rect 16120 13184 16172 13190
rect 16120 13126 16172 13132
rect 15844 12572 15896 12578
rect 15844 12514 15896 12520
rect 15842 12362 15898 12371
rect 15842 12297 15898 12306
rect 15660 12096 15712 12102
rect 15660 12038 15712 12044
rect 15476 12028 15528 12034
rect 15474 11996 15476 12005
rect 15568 12028 15620 12034
rect 15528 11996 15530 12005
rect 15568 11970 15620 11976
rect 15474 11931 15530 11940
rect 15580 11880 15608 11970
rect 15488 11852 15608 11880
rect 14840 11724 15460 11744
rect 14840 11668 14882 11724
rect 14938 11668 14962 11724
rect 15018 11668 15042 11724
rect 15098 11668 15122 11724
rect 15178 11668 15202 11724
rect 15258 11668 15282 11724
rect 15338 11668 15362 11724
rect 15418 11668 15460 11724
rect 14840 11648 15460 11668
rect 15488 11422 15516 11852
rect 15856 11422 15884 12297
rect 15476 11416 15528 11422
rect 15476 11358 15528 11364
rect 15844 11416 15896 11422
rect 15844 11358 15896 11364
rect 14840 10636 15460 10656
rect 14840 10580 14882 10636
rect 14938 10580 14962 10636
rect 15018 10580 15042 10636
rect 15098 10580 15122 10636
rect 15178 10580 15202 10636
rect 15258 10580 15282 10636
rect 15338 10580 15362 10636
rect 15418 10580 15460 10636
rect 14840 10560 15460 10580
rect 15488 10520 15516 11358
rect 15752 11348 15804 11354
rect 15752 11290 15804 11296
rect 15764 11082 15792 11290
rect 15752 11076 15804 11082
rect 15752 11018 15804 11024
rect 15856 10928 15884 11358
rect 15304 10492 15516 10520
rect 15764 10900 15884 10928
rect 15936 10940 15988 10946
rect 15304 10334 15332 10492
rect 15764 10419 15792 10900
rect 15936 10882 15988 10888
rect 15750 10410 15806 10419
rect 15750 10345 15806 10354
rect 15292 10328 15344 10334
rect 15292 10270 15344 10276
rect 14924 10192 14976 10198
rect 14924 10134 14976 10140
rect 14936 9926 14964 10134
rect 14924 9920 14976 9926
rect 14924 9862 14976 9868
rect 15304 9858 15332 10270
rect 15292 9852 15344 9858
rect 15292 9794 15344 9800
rect 15568 9852 15620 9858
rect 15568 9794 15620 9800
rect 14840 9548 15460 9568
rect 14840 9492 14882 9548
rect 14938 9492 14962 9548
rect 15018 9492 15042 9548
rect 15098 9492 15122 9548
rect 15178 9492 15202 9548
rect 15258 9492 15282 9548
rect 15338 9492 15362 9548
rect 15418 9492 15460 9548
rect 14840 9472 15460 9492
rect 15580 9432 15608 9794
rect 15764 9790 15792 10345
rect 15752 9784 15804 9790
rect 15752 9726 15804 9732
rect 15764 9568 15792 9726
rect 15948 9722 15976 10882
rect 16132 10538 16160 13126
rect 16120 10532 16172 10538
rect 16120 10474 16172 10480
rect 16120 10260 16172 10266
rect 16120 10202 16172 10208
rect 16028 9852 16080 9858
rect 16028 9794 16080 9800
rect 15936 9716 15988 9722
rect 15936 9658 15988 9664
rect 15764 9540 15884 9568
rect 15396 9404 15608 9432
rect 15658 9434 15714 9443
rect 15396 8906 15424 9404
rect 15658 9369 15714 9378
rect 15384 8900 15436 8906
rect 15384 8842 15436 8848
rect 15474 8824 15530 8833
rect 15474 8764 15530 8768
rect 15474 8759 15476 8764
rect 15528 8759 15530 8764
rect 15476 8706 15528 8712
rect 14840 8460 15460 8480
rect 14840 8404 14882 8460
rect 14938 8404 14962 8460
rect 15018 8404 15042 8460
rect 15098 8404 15122 8460
rect 15178 8404 15202 8460
rect 15258 8404 15282 8460
rect 15338 8404 15362 8460
rect 15418 8404 15460 8460
rect 14840 8384 15460 8404
rect 15016 8152 15068 8158
rect 15016 8094 15068 8100
rect 14832 8084 14884 8090
rect 14752 8044 14832 8072
rect 14464 8016 14516 8022
rect 14464 7958 14516 7964
rect 14476 7682 14504 7958
rect 14646 7726 14702 7735
rect 14464 7676 14516 7682
rect 14752 7682 14780 8044
rect 14832 8026 14884 8032
rect 14646 7661 14702 7670
rect 14740 7676 14792 7682
rect 14464 7618 14516 7624
rect 14660 6594 14688 7661
rect 14740 7618 14792 7624
rect 15028 7528 15056 8094
rect 15200 8084 15252 8090
rect 15200 8026 15252 8032
rect 15212 7818 15240 8026
rect 15200 7812 15252 7818
rect 15200 7754 15252 7760
rect 14752 7500 15056 7528
rect 14752 7274 14780 7500
rect 14840 7372 15460 7392
rect 14840 7316 14882 7372
rect 14938 7316 14962 7372
rect 15018 7316 15042 7372
rect 15098 7316 15122 7372
rect 15178 7316 15202 7372
rect 15258 7316 15282 7372
rect 15338 7316 15362 7372
rect 15418 7316 15460 7372
rect 14840 7296 15460 7316
rect 14740 7268 14792 7274
rect 14740 7210 14792 7216
rect 15672 7206 15700 9369
rect 15856 9246 15884 9540
rect 15844 9240 15896 9246
rect 15844 9182 15896 9188
rect 16040 8833 16068 9794
rect 16132 9450 16160 10202
rect 16316 9687 16344 15030
rect 16500 14686 16528 16952
rect 16672 16788 16724 16794
rect 16672 16730 16724 16736
rect 16684 16522 16712 16730
rect 16672 16516 16724 16522
rect 16672 16458 16724 16464
rect 16670 16388 16726 16397
rect 16670 16328 16672 16332
rect 16724 16328 16726 16332
rect 16670 16323 16726 16328
rect 16672 16322 16724 16323
rect 16684 16300 16712 16322
rect 16868 16318 16896 17206
rect 16856 16312 16908 16318
rect 16856 16254 16908 16260
rect 16868 15910 16896 16254
rect 16856 15904 16908 15910
rect 16856 15846 16908 15852
rect 16672 15836 16724 15842
rect 16672 15778 16724 15784
rect 16488 14680 16540 14686
rect 16488 14622 16540 14628
rect 16684 14464 16712 15778
rect 16868 15298 16896 15846
rect 16948 15768 17000 15774
rect 16948 15710 17000 15716
rect 16960 15434 16988 15710
rect 16948 15428 17000 15434
rect 16948 15370 17000 15376
rect 16856 15292 16908 15298
rect 16856 15234 16908 15240
rect 16592 14436 16712 14464
rect 16592 14142 16620 14436
rect 16960 14210 16988 15370
rect 17144 14346 17172 17342
rect 17328 15909 17356 17886
rect 17314 15900 17370 15909
rect 17314 15835 17370 15844
rect 17328 15700 17356 15835
rect 17512 15824 17540 18380
rect 17696 18086 17724 18430
rect 17880 18340 17908 18498
rect 18420 18352 18472 18358
rect 17880 18312 18000 18340
rect 17684 18080 17736 18086
rect 17684 18022 17736 18028
rect 17696 17861 17724 18022
rect 17682 17852 17738 17861
rect 17682 17787 17738 17796
rect 17696 17474 17724 17787
rect 17972 17660 18000 18312
rect 18420 18294 18472 18300
rect 18880 18352 18932 18358
rect 18880 18294 18932 18300
rect 17880 17632 18000 17660
rect 17880 17495 17908 17632
rect 17866 17486 17922 17495
rect 17684 17468 17736 17474
rect 17866 17421 17922 17430
rect 17684 17410 17736 17416
rect 17880 17270 17908 17421
rect 17868 17264 17920 17270
rect 17868 17206 17920 17212
rect 18144 16924 18196 16930
rect 17972 16884 18144 16912
rect 17776 16788 17828 16794
rect 17776 16730 17828 16736
rect 17788 16522 17816 16730
rect 17776 16516 17828 16522
rect 17776 16458 17828 16464
rect 17972 16318 18000 16884
rect 18144 16866 18196 16872
rect 18432 16862 18460 18294
rect 18892 18136 18920 18294
rect 18800 18108 18920 18136
rect 18800 17456 18828 18108
rect 18800 17428 18920 17456
rect 18604 17264 18656 17270
rect 18604 17206 18656 17212
rect 18420 16856 18472 16862
rect 18420 16798 18472 16804
rect 18616 16454 18644 17206
rect 18604 16448 18656 16454
rect 18604 16390 18656 16396
rect 17960 16312 18012 16318
rect 17960 16254 18012 16260
rect 17420 15796 17540 15824
rect 17310 15648 17316 15700
rect 17368 15648 17374 15700
rect 17316 15088 17368 15094
rect 17316 15030 17368 15036
rect 17328 14668 17356 15030
rect 17420 14890 17448 15796
rect 17776 15632 17828 15638
rect 17776 15574 17828 15580
rect 17408 14884 17460 14890
rect 17408 14826 17460 14832
rect 17328 14640 17448 14668
rect 17132 14340 17184 14346
rect 17132 14282 17184 14288
rect 16948 14204 17000 14210
rect 17420 14192 17448 14640
rect 16948 14146 17000 14152
rect 17328 14164 17448 14192
rect 16580 14136 16632 14142
rect 16580 14078 16632 14084
rect 16396 9920 16448 9926
rect 16396 9862 16448 9868
rect 16302 9678 16358 9687
rect 16302 9613 16358 9622
rect 16120 9444 16172 9450
rect 16120 9386 16172 9392
rect 16408 9296 16436 9862
rect 16362 9268 16436 9296
rect 16592 9296 16620 14078
rect 16960 13648 16988 14146
rect 16868 13620 16988 13648
rect 16868 13172 16896 13620
rect 17132 13524 17184 13530
rect 17132 13466 17184 13472
rect 16868 13144 16942 13172
rect 16762 12972 16818 12981
rect 16762 12907 16818 12916
rect 16776 12714 16804 12907
rect 16764 12708 16816 12714
rect 16764 12650 16816 12656
rect 16762 12606 16818 12615
rect 16762 12541 16818 12550
rect 16776 12510 16804 12541
rect 16764 12504 16816 12510
rect 16764 12446 16816 12452
rect 16764 12368 16816 12374
rect 16764 12310 16816 12316
rect 16776 12170 16804 12310
rect 16764 12164 16816 12170
rect 16764 12106 16816 12112
rect 16914 11608 16942 13144
rect 17040 12912 17092 12918
rect 17040 12854 17092 12860
rect 17052 11812 17080 12854
rect 17144 12714 17172 13466
rect 17328 13258 17356 14164
rect 17788 13598 17816 15574
rect 17972 15230 18000 16254
rect 18604 15768 18656 15774
rect 18604 15710 18656 15716
rect 18616 15298 18644 15710
rect 18892 15416 18920 17428
rect 19076 17338 19104 18992
rect 19200 18796 19820 18816
rect 19200 18740 19242 18796
rect 19298 18740 19322 18796
rect 19378 18740 19402 18796
rect 19458 18740 19482 18796
rect 19538 18740 19562 18796
rect 19618 18740 19642 18796
rect 19698 18740 19722 18796
rect 19778 18740 19820 18796
rect 19200 18720 19820 18740
rect 20076 18692 20128 18698
rect 20076 18634 20128 18640
rect 19892 18488 19944 18494
rect 19892 18430 19944 18436
rect 19794 17892 19800 17944
rect 19852 17892 19858 17944
rect 19812 17861 19840 17892
rect 19798 17852 19854 17861
rect 19904 17838 19932 18430
rect 19854 17810 19932 17838
rect 19798 17787 19854 17796
rect 19200 17708 19820 17728
rect 19200 17652 19242 17708
rect 19298 17652 19322 17708
rect 19378 17652 19402 17708
rect 19458 17652 19482 17708
rect 19538 17652 19562 17708
rect 19618 17652 19642 17708
rect 19698 17652 19722 17708
rect 19778 17652 19820 17708
rect 19200 17632 19820 17652
rect 19708 17536 19760 17542
rect 19522 17486 19578 17495
rect 19708 17478 19760 17484
rect 19522 17421 19524 17430
rect 19576 17421 19578 17430
rect 19524 17410 19576 17416
rect 19064 17332 19116 17338
rect 19064 17274 19116 17280
rect 19076 16436 19104 17274
rect 19536 16885 19564 17410
rect 19720 17066 19748 17478
rect 19708 17060 19760 17066
rect 19708 17002 19760 17008
rect 19522 16876 19578 16885
rect 19522 16811 19578 16820
rect 19200 16620 19820 16640
rect 19200 16564 19242 16620
rect 19298 16564 19322 16620
rect 19378 16564 19402 16620
rect 19458 16564 19482 16620
rect 19538 16564 19562 16620
rect 19618 16564 19642 16620
rect 19698 16564 19722 16620
rect 19778 16564 19820 16620
rect 19200 16544 19820 16564
rect 19076 16408 19196 16436
rect 19168 15960 19196 16408
rect 19904 16386 19932 17810
rect 20088 16930 20116 18634
rect 20180 18630 20208 19042
rect 20364 19038 20392 19468
rect 20440 19340 21060 19360
rect 20440 19284 20482 19340
rect 20538 19284 20562 19340
rect 20618 19284 20642 19340
rect 20698 19284 20722 19340
rect 20778 19284 20802 19340
rect 20858 19284 20882 19340
rect 20938 19284 20962 19340
rect 21018 19284 21060 19340
rect 20440 19264 21060 19284
rect 20352 19032 20404 19038
rect 20352 18974 20404 18980
rect 20904 18896 20956 18902
rect 20904 18838 20956 18844
rect 20916 18698 20944 18838
rect 20904 18692 20956 18698
rect 20904 18634 20956 18640
rect 20168 18624 20220 18630
rect 20168 18566 20220 18572
rect 20352 18352 20404 18358
rect 20352 18294 20404 18300
rect 20168 17264 20220 17270
rect 20168 17206 20220 17212
rect 20076 16924 20128 16930
rect 20076 16866 20128 16872
rect 20180 16726 20208 17206
rect 20076 16720 20128 16726
rect 20076 16662 20128 16668
rect 20168 16720 20220 16726
rect 20168 16662 20220 16668
rect 20088 16397 20116 16662
rect 20364 16454 20392 18294
rect 20440 18252 21060 18272
rect 20440 18196 20482 18252
rect 20538 18196 20562 18252
rect 20618 18196 20642 18252
rect 20698 18196 20722 18252
rect 20778 18196 20802 18252
rect 20858 18196 20882 18252
rect 20938 18196 20962 18252
rect 21018 18196 21060 18252
rect 20440 18176 21060 18196
rect 21100 18068 21128 21694
rect 21284 21214 21312 21762
rect 21640 21616 21692 21622
rect 21640 21558 21692 21564
rect 21456 21276 21508 21282
rect 21456 21218 21508 21224
rect 21272 21208 21324 21214
rect 21272 21150 21324 21156
rect 21468 20992 21496 21218
rect 21376 20964 21496 20992
rect 21376 19088 21404 20964
rect 21376 19060 21496 19088
rect 21272 18896 21324 18902
rect 21272 18838 21324 18844
rect 21008 18040 21128 18068
rect 21008 17524 21036 18040
rect 21008 17496 21128 17524
rect 21100 17338 21128 17496
rect 21088 17332 21140 17338
rect 21088 17274 21140 17280
rect 20440 17164 21060 17184
rect 20440 17108 20482 17164
rect 20538 17108 20562 17164
rect 20618 17108 20642 17164
rect 20698 17108 20722 17164
rect 20778 17108 20802 17164
rect 20858 17108 20882 17164
rect 20938 17108 20962 17164
rect 21018 17108 21060 17164
rect 20440 17088 21060 17108
rect 20902 16876 20958 16885
rect 20902 16811 20904 16820
rect 20956 16811 20958 16820
rect 20904 16798 20956 16804
rect 20720 16788 20772 16794
rect 20916 16788 20944 16798
rect 20720 16730 20772 16736
rect 20732 16522 20760 16730
rect 20996 16720 21048 16726
rect 20996 16662 21048 16668
rect 20720 16516 20772 16522
rect 20720 16458 20772 16464
rect 20352 16448 20404 16454
rect 20074 16388 20130 16397
rect 20352 16390 20404 16396
rect 19892 16380 19944 16386
rect 19892 16322 19944 16328
rect 20074 16323 20130 16332
rect 19076 15932 19196 15960
rect 19076 15774 19104 15932
rect 20088 15842 20116 16323
rect 20076 15836 20128 15842
rect 20076 15778 20128 15784
rect 19064 15768 19116 15774
rect 19064 15710 19116 15716
rect 19064 15632 19116 15638
rect 19064 15574 19116 15580
rect 18972 15428 19024 15434
rect 18892 15388 18972 15416
rect 18972 15370 19024 15376
rect 18604 15292 18656 15298
rect 18604 15234 18656 15240
rect 17960 15224 18012 15230
rect 17960 15166 18012 15172
rect 18510 15168 18566 15177
rect 17972 14872 18000 15166
rect 18510 15103 18566 15112
rect 18524 14872 18552 15103
rect 17972 14844 18552 14872
rect 17972 14689 18000 14844
rect 18236 14748 18288 14754
rect 18236 14690 18288 14696
rect 17958 14680 18014 14689
rect 17958 14615 18014 14624
rect 17972 13666 18000 14615
rect 18248 13920 18276 14690
rect 18524 14686 18552 14844
rect 19076 14811 19104 15574
rect 19200 15532 19820 15552
rect 19200 15476 19242 15532
rect 19298 15476 19322 15532
rect 19378 15476 19402 15532
rect 19458 15476 19482 15532
rect 19538 15476 19562 15532
rect 19618 15476 19642 15532
rect 19698 15476 19722 15532
rect 19778 15476 19820 15532
rect 19200 15456 19820 15476
rect 19800 15156 19852 15162
rect 19800 15098 19852 15104
rect 19062 14802 19118 14811
rect 18782 14696 18788 14748
rect 18840 14696 18846 14748
rect 19062 14737 19118 14746
rect 18512 14680 18564 14686
rect 18512 14622 18564 14628
rect 18604 14612 18656 14618
rect 18604 14554 18656 14560
rect 18616 14210 18644 14554
rect 18800 14210 18828 14696
rect 18972 14612 19024 14618
rect 18972 14554 19024 14560
rect 18984 14346 19012 14554
rect 18972 14340 19024 14346
rect 18972 14282 19024 14288
rect 19076 14210 19104 14737
rect 19812 14600 19840 15098
rect 19984 15088 20036 15094
rect 19984 15030 20036 15036
rect 19996 14618 20024 15030
rect 20088 14680 20116 15778
rect 20364 14822 20392 16390
rect 21008 16232 21036 16662
rect 21284 16397 21312 18838
rect 21468 17950 21496 19060
rect 21652 18630 21680 21558
rect 21640 18624 21692 18630
rect 21640 18566 21692 18572
rect 21836 18358 21864 25229
rect 26422 22732 26478 22741
rect 26422 22667 26478 22676
rect 22742 21878 22798 21887
rect 22742 21820 22798 21822
rect 22742 21813 22744 21820
rect 22796 21813 22798 21820
rect 22744 21762 22796 21768
rect 22008 21752 22060 21758
rect 22008 21694 22060 21700
rect 22020 21418 22048 21694
rect 22376 21616 22428 21622
rect 22376 21558 22428 21564
rect 22008 21412 22060 21418
rect 22388 21400 22416 21558
rect 22388 21372 22508 21400
rect 22008 21354 22060 21360
rect 22192 21344 22244 21350
rect 22192 21286 22244 21292
rect 22008 20664 22060 20670
rect 22008 20606 22060 20612
rect 22020 19904 22048 20606
rect 22204 19972 22232 21286
rect 22480 20924 22508 21372
rect 22388 20896 22508 20924
rect 22204 19944 22278 19972
rect 22020 19876 22140 19904
rect 22008 19780 22060 19786
rect 22008 19722 22060 19728
rect 22020 19564 22048 19722
rect 21974 19536 22048 19564
rect 21974 19020 22002 19536
rect 22112 19203 22140 19876
rect 22250 19428 22278 19944
rect 22204 19400 22278 19428
rect 22204 19242 22232 19400
rect 22192 19236 22244 19242
rect 22098 19194 22154 19203
rect 22192 19178 22244 19184
rect 22098 19129 22154 19138
rect 22112 19088 22140 19129
rect 22112 19060 22232 19088
rect 21974 18992 22048 19020
rect 21824 18352 21876 18358
rect 22020 18340 22048 18992
rect 22204 18562 22232 19060
rect 22192 18556 22244 18562
rect 22192 18498 22244 18504
rect 22020 18312 22140 18340
rect 21824 18294 21876 18300
rect 21456 17944 21508 17950
rect 21456 17886 21508 17892
rect 21456 17808 21508 17814
rect 21456 17750 21508 17756
rect 21468 16794 21496 17750
rect 21638 17730 21694 17739
rect 21638 17665 21694 17674
rect 21652 17388 21680 17665
rect 21836 17610 21864 18294
rect 22112 17660 22140 18312
rect 22020 17632 22140 17660
rect 21824 17604 21876 17610
rect 21824 17546 21876 17552
rect 21652 17360 21772 17388
rect 21456 16788 21508 16794
rect 21456 16730 21508 16736
rect 21744 16708 21772 17360
rect 21652 16680 21772 16708
rect 21652 16522 21680 16680
rect 21640 16516 21692 16522
rect 21640 16458 21692 16464
rect 21270 16388 21326 16397
rect 21270 16323 21326 16332
rect 21008 16204 21128 16232
rect 20440 16076 21060 16096
rect 20440 16020 20482 16076
rect 20538 16020 20562 16076
rect 20618 16020 20642 16076
rect 20698 16020 20722 16076
rect 20778 16020 20802 16076
rect 20858 16020 20882 16076
rect 20938 16020 20962 16076
rect 21018 16020 21060 16076
rect 20440 16000 21060 16020
rect 21100 15960 21128 16204
rect 21272 16176 21324 16182
rect 21272 16118 21324 16124
rect 21008 15932 21128 15960
rect 21008 15774 21036 15932
rect 20996 15768 21048 15774
rect 20996 15710 21048 15716
rect 21088 15360 21140 15366
rect 21088 15302 21140 15308
rect 20440 14988 21060 15008
rect 20440 14932 20482 14988
rect 20538 14932 20562 14988
rect 20618 14932 20642 14988
rect 20698 14932 20722 14988
rect 20778 14932 20802 14988
rect 20858 14932 20882 14988
rect 20938 14932 20962 14988
rect 21018 14932 21060 14988
rect 20440 14912 21060 14932
rect 20990 14832 20996 14884
rect 21048 14872 21054 14884
rect 21100 14872 21128 15302
rect 21048 14844 21128 14872
rect 21048 14832 21054 14844
rect 20352 14816 20404 14822
rect 20352 14758 20404 14764
rect 20626 14802 20682 14811
rect 20444 14748 20496 14754
rect 20626 14737 20682 14746
rect 20444 14690 20496 14696
rect 20070 14628 20076 14680
rect 20128 14628 20134 14680
rect 20346 14628 20352 14680
rect 20404 14628 20410 14680
rect 19984 14612 20036 14618
rect 19812 14572 19932 14600
rect 19200 14444 19820 14464
rect 19200 14388 19242 14444
rect 19298 14388 19322 14444
rect 19378 14388 19402 14444
rect 19458 14388 19482 14444
rect 19538 14388 19562 14444
rect 19618 14388 19642 14444
rect 19698 14388 19722 14444
rect 19778 14388 19820 14444
rect 19200 14368 19820 14388
rect 18604 14204 18656 14210
rect 18604 14146 18656 14152
rect 18788 14204 18840 14210
rect 18788 14146 18840 14152
rect 19064 14204 19116 14210
rect 19064 14146 19116 14152
rect 18248 13892 18368 13920
rect 18340 13802 18368 13892
rect 18328 13796 18380 13802
rect 18328 13738 18380 13744
rect 17960 13660 18012 13666
rect 18800 13660 18828 14146
rect 19076 13713 19104 14146
rect 19904 14142 19932 14572
rect 19984 14554 20036 14560
rect 20168 14544 20220 14550
rect 20168 14486 20220 14492
rect 19892 14136 19944 14142
rect 19892 14078 19944 14084
rect 19062 13704 19118 13713
rect 18782 13608 18788 13660
rect 18840 13608 18846 13660
rect 19062 13639 19118 13648
rect 19892 13660 19944 13666
rect 17960 13602 18012 13608
rect 17776 13592 17828 13598
rect 17776 13534 17828 13540
rect 17316 13252 17368 13258
rect 18800 13225 18828 13608
rect 19892 13602 19944 13608
rect 19200 13356 19820 13376
rect 19200 13300 19242 13356
rect 19298 13300 19322 13356
rect 19378 13300 19402 13356
rect 19458 13300 19482 13356
rect 19538 13300 19562 13356
rect 19618 13300 19642 13356
rect 19698 13300 19722 13356
rect 19778 13300 19820 13356
rect 19200 13280 19820 13300
rect 17316 13194 17368 13200
rect 17498 13216 17554 13225
rect 17498 13151 17554 13160
rect 18786 13216 18842 13225
rect 18786 13151 18842 13160
rect 17512 13122 17540 13151
rect 18800 13122 18828 13151
rect 17224 13116 17276 13122
rect 17500 13116 17552 13122
rect 17276 13076 17356 13104
rect 17224 13058 17276 13064
rect 17132 12708 17184 12714
rect 17132 12650 17184 12656
rect 17132 12504 17184 12510
rect 17132 12446 17184 12452
rect 17144 12034 17172 12446
rect 17132 12028 17184 12034
rect 17132 11970 17184 11976
rect 17328 11898 17356 13076
rect 17500 13058 17552 13064
rect 18788 13116 18840 13122
rect 18788 13058 18840 13064
rect 17500 12912 17552 12918
rect 17500 12854 17552 12860
rect 17512 12615 17540 12854
rect 17498 12606 17554 12615
rect 17498 12541 17554 12550
rect 18602 12606 18658 12615
rect 18800 12578 18828 13058
rect 18602 12541 18658 12550
rect 18788 12572 18840 12578
rect 17960 12368 18012 12374
rect 17960 12310 18012 12316
rect 17972 12102 18000 12310
rect 17500 12096 17552 12102
rect 17500 12038 17552 12044
rect 17960 12096 18012 12102
rect 17960 12038 18012 12044
rect 17316 11892 17368 11898
rect 17512 11880 17540 12038
rect 18512 11960 18564 11966
rect 18512 11902 18564 11908
rect 17316 11834 17368 11840
rect 17466 11852 17540 11880
rect 18236 11892 18288 11898
rect 17052 11784 17172 11812
rect 16914 11580 16988 11608
rect 16856 11416 16908 11422
rect 16856 11358 16908 11364
rect 16868 10878 16896 11358
rect 16856 10872 16908 10878
rect 16856 10814 16908 10820
rect 16868 10663 16896 10814
rect 16854 10654 16910 10663
rect 16854 10589 16910 10598
rect 16868 10334 16896 10589
rect 16856 10328 16908 10334
rect 16856 10270 16908 10276
rect 16960 10112 16988 11580
rect 17144 10384 17172 11784
rect 17316 11280 17368 11286
rect 17466 11268 17494 11852
rect 18236 11834 18288 11840
rect 17592 11824 17644 11830
rect 17592 11766 17644 11772
rect 17604 11422 17632 11766
rect 17592 11416 17644 11422
rect 17592 11358 17644 11364
rect 17868 11280 17920 11286
rect 17466 11240 17540 11268
rect 17316 11222 17368 11228
rect 16914 10084 16988 10112
rect 17098 10356 17172 10384
rect 16764 9852 16816 9858
rect 16764 9794 16816 9800
rect 16592 9268 16666 9296
rect 16026 8824 16082 8833
rect 16026 8759 16082 8768
rect 16212 8764 16264 8770
rect 16040 7818 16068 8759
rect 16362 8752 16390 9268
rect 16488 9172 16540 9178
rect 16488 9114 16540 9120
rect 16500 8906 16528 9114
rect 16488 8900 16540 8906
rect 16488 8842 16540 8848
rect 16638 8820 16666 9268
rect 16776 9246 16804 9794
rect 16914 9500 16942 10084
rect 17098 9840 17126 10356
rect 17328 10266 17356 11222
rect 17316 10260 17368 10266
rect 17316 10202 17368 10208
rect 17224 10192 17276 10198
rect 17224 10134 17276 10140
rect 17052 9812 17126 9840
rect 17052 9654 17080 9812
rect 17040 9648 17092 9654
rect 17040 9590 17092 9596
rect 16914 9472 16988 9500
rect 16764 9240 16816 9246
rect 16764 9182 16816 9188
rect 16592 8792 16666 8820
rect 16362 8724 16436 8752
rect 16212 8706 16264 8712
rect 16224 8589 16252 8706
rect 16210 8580 16266 8589
rect 16210 8515 16266 8524
rect 16028 7812 16080 7818
rect 16028 7754 16080 7760
rect 16210 7726 16266 7735
rect 16210 7661 16266 7670
rect 15660 7200 15712 7206
rect 15660 7142 15712 7148
rect 16224 7138 16252 7661
rect 16212 7132 16264 7138
rect 16212 7074 16264 7080
rect 14648 6588 14700 6594
rect 14648 6530 14700 6536
rect 16212 6384 16264 6390
rect 16212 6326 16264 6332
rect 14840 6284 15460 6304
rect 14840 6228 14882 6284
rect 14938 6228 14962 6284
rect 15018 6228 15042 6284
rect 15098 6228 15122 6284
rect 15178 6228 15202 6284
rect 15258 6228 15282 6284
rect 15338 6228 15362 6284
rect 15418 6228 15460 6284
rect 14840 6208 15460 6228
rect 16224 6118 16252 6326
rect 16408 6168 16436 8724
rect 16592 8616 16620 8792
rect 16672 8628 16724 8634
rect 16592 8588 16672 8616
rect 16592 7546 16620 8588
rect 16672 8570 16724 8576
rect 16776 8294 16804 9182
rect 16960 8838 16988 9472
rect 16948 8832 17000 8838
rect 16948 8774 17000 8780
rect 17038 8580 17094 8589
rect 17038 8515 17094 8524
rect 16764 8288 16816 8294
rect 16764 8230 16816 8236
rect 17052 8072 17080 8515
rect 17236 8362 17264 10134
rect 17512 9994 17540 11240
rect 17868 11222 17920 11228
rect 18052 11280 18104 11286
rect 18052 11222 18104 11228
rect 17684 10464 17736 10470
rect 17684 10406 17736 10412
rect 17500 9988 17552 9994
rect 17500 9930 17552 9936
rect 17408 9648 17460 9654
rect 17408 9590 17460 9596
rect 17224 8356 17276 8362
rect 17224 8298 17276 8304
rect 16868 8044 17080 8072
rect 16580 7540 16632 7546
rect 16580 7482 16632 7488
rect 16868 7460 16896 8044
rect 17130 7970 17186 7979
rect 17130 7905 17186 7914
rect 17144 7614 17172 7905
rect 17420 7614 17448 9590
rect 17696 9246 17724 10406
rect 17684 9240 17736 9246
rect 17684 9182 17736 9188
rect 17592 8560 17644 8566
rect 17592 8502 17644 8508
rect 17604 8294 17632 8502
rect 17592 8288 17644 8294
rect 17592 8230 17644 8236
rect 17880 8072 17908 11222
rect 17958 10410 18014 10419
rect 17958 10345 17960 10354
rect 18012 10345 18014 10354
rect 17960 10338 18012 10344
rect 17972 10322 18000 10338
rect 18064 10334 18092 11222
rect 18248 10538 18276 11834
rect 18420 10940 18472 10946
rect 18524 10928 18552 11902
rect 18472 10900 18552 10928
rect 18420 10882 18472 10888
rect 18524 10663 18552 10900
rect 18510 10654 18566 10663
rect 18510 10589 18566 10598
rect 18236 10532 18288 10538
rect 18236 10474 18288 10480
rect 18052 10328 18104 10334
rect 18052 10270 18104 10276
rect 18144 10192 18196 10198
rect 18142 10166 18144 10175
rect 18196 10166 18198 10175
rect 18142 10101 18198 10110
rect 18248 9994 18276 10474
rect 18052 9988 18104 9994
rect 18052 9931 18104 9936
rect 18236 9988 18288 9994
rect 18050 9922 18106 9931
rect 18236 9930 18288 9936
rect 18050 9857 18106 9866
rect 18064 8344 18092 9857
rect 18328 9852 18380 9858
rect 18328 9794 18380 9800
rect 18340 8770 18368 9794
rect 18524 9172 18552 10589
rect 18506 9120 18512 9172
rect 18564 9120 18570 9172
rect 18328 8764 18380 8770
rect 18328 8706 18380 8712
rect 18236 8356 18288 8362
rect 18064 8316 18236 8344
rect 18236 8298 18288 8304
rect 18052 8152 18104 8158
rect 18052 8094 18104 8100
rect 17788 8044 17908 8072
rect 17132 7608 17184 7614
rect 17132 7550 17184 7556
rect 17408 7608 17460 7614
rect 17408 7550 17460 7556
rect 17788 7460 17816 8044
rect 18064 7614 18092 8094
rect 18340 7682 18368 8706
rect 18524 8634 18552 9120
rect 18512 8628 18564 8634
rect 18512 8570 18564 8576
rect 18524 8158 18552 8570
rect 18512 8152 18564 8158
rect 18512 8094 18564 8100
rect 18616 7682 18644 12541
rect 18788 12514 18840 12520
rect 18972 12436 19024 12442
rect 18972 12378 19024 12384
rect 18788 11416 18840 11422
rect 18788 11358 18840 11364
rect 18800 10396 18828 11358
rect 18782 10344 18788 10396
rect 18840 10344 18846 10396
rect 18696 9240 18748 9246
rect 18696 9182 18748 9188
rect 18708 8833 18736 9182
rect 18694 8824 18750 8833
rect 18694 8759 18750 8768
rect 18800 7735 18828 10344
rect 18984 8362 19012 12378
rect 19200 12268 19820 12288
rect 19200 12212 19242 12268
rect 19298 12212 19322 12268
rect 19378 12212 19402 12268
rect 19458 12212 19482 12268
rect 19538 12212 19562 12268
rect 19618 12212 19642 12268
rect 19698 12212 19722 12268
rect 19778 12212 19820 12268
rect 19200 12192 19820 12212
rect 19904 12084 19932 13602
rect 20180 13462 20208 14486
rect 20364 14210 20392 14628
rect 20456 14567 20484 14690
rect 20442 14558 20498 14567
rect 20640 14550 20668 14737
rect 21284 14567 21312 16118
rect 21456 15768 21508 15774
rect 21456 15710 21508 15716
rect 21468 15230 21496 15710
rect 21916 15700 21968 15706
rect 22020 15688 22048 17632
rect 22192 17468 22244 17474
rect 22192 17410 22244 17416
rect 22204 16522 22232 17410
rect 22388 16522 22416 20896
rect 22560 20732 22612 20738
rect 22560 20674 22612 20680
rect 22572 18136 22600 20674
rect 22928 20188 22980 20194
rect 22742 20170 22798 20179
rect 22742 20105 22798 20114
rect 22848 20148 22928 20176
rect 22756 20040 22784 20105
rect 22848 20040 22876 20148
rect 22928 20130 22980 20136
rect 22756 20012 22876 20040
rect 22928 20052 22980 20058
rect 22756 19582 22784 20012
rect 22928 19994 22980 20000
rect 22940 19836 22968 19994
rect 22940 19808 23060 19836
rect 22744 19576 22796 19582
rect 22744 19518 22796 19524
rect 22756 19038 22784 19518
rect 22744 19032 22796 19038
rect 22744 18974 22796 18980
rect 22480 18108 22600 18136
rect 22480 17950 22508 18108
rect 22756 18012 22784 18974
rect 23032 18884 23060 19808
rect 22940 18856 23060 18884
rect 22940 18698 22968 18856
rect 22928 18692 22980 18698
rect 22928 18634 22980 18640
rect 22928 18556 22980 18562
rect 22928 18498 22980 18504
rect 22940 18340 22968 18498
rect 22940 18312 23060 18340
rect 22738 17960 22744 18012
rect 22796 17960 22802 18012
rect 22468 17944 22520 17950
rect 22468 17886 22520 17892
rect 22756 17474 22784 17960
rect 22744 17468 22796 17474
rect 22744 17410 22796 17416
rect 22192 16516 22244 16522
rect 22192 16458 22244 16464
rect 22376 16516 22428 16522
rect 22376 16458 22428 16464
rect 22284 16312 22336 16318
rect 22284 16254 22336 16260
rect 22020 15660 22140 15688
rect 21916 15642 21968 15648
rect 21732 15632 21784 15638
rect 21732 15574 21784 15580
rect 21456 15224 21508 15230
rect 21454 15172 21456 15177
rect 21508 15172 21510 15177
rect 21454 15168 21510 15172
rect 21454 15103 21510 15112
rect 21270 14558 21326 14567
rect 20442 14493 20498 14502
rect 20628 14544 20680 14550
rect 21270 14493 21326 14502
rect 20628 14486 20680 14492
rect 21270 14314 21326 14323
rect 21270 14249 21326 14258
rect 21284 14210 21312 14249
rect 20352 14204 20404 14210
rect 20352 14146 20404 14152
rect 21272 14204 21324 14210
rect 21272 14146 21324 14152
rect 21456 14204 21508 14210
rect 21456 14146 21508 14152
rect 20364 13784 20392 14146
rect 20440 13900 21060 13920
rect 20440 13844 20482 13900
rect 20538 13844 20562 13900
rect 20618 13844 20642 13900
rect 20698 13844 20722 13900
rect 20778 13844 20802 13900
rect 20858 13844 20882 13900
rect 20938 13844 20962 13900
rect 21018 13844 21060 13900
rect 20440 13824 21060 13844
rect 20364 13756 20760 13784
rect 20442 13704 20498 13713
rect 20442 13639 20498 13648
rect 20456 13598 20484 13639
rect 20732 13598 20760 13756
rect 20444 13592 20496 13598
rect 20444 13534 20496 13540
rect 20720 13592 20772 13598
rect 20720 13534 20772 13540
rect 20168 13456 20220 13462
rect 20168 13398 20220 13404
rect 20456 13122 20484 13534
rect 20536 13524 20588 13530
rect 20536 13466 20588 13472
rect 20548 13258 20576 13466
rect 20732 13376 20760 13534
rect 20732 13348 20852 13376
rect 20536 13252 20588 13258
rect 20824 13225 20852 13348
rect 20536 13194 20588 13200
rect 20810 13216 20866 13225
rect 20444 13116 20496 13122
rect 20364 13076 20444 13104
rect 20168 12912 20220 12918
rect 20168 12854 20220 12860
rect 20180 12696 20208 12854
rect 20088 12668 20208 12696
rect 20088 12102 20116 12668
rect 20166 12606 20222 12615
rect 20166 12541 20222 12550
rect 20180 12510 20208 12541
rect 20168 12504 20220 12510
rect 20168 12446 20220 12452
rect 19812 12056 19932 12084
rect 20076 12096 20128 12102
rect 19812 11948 19840 12056
rect 20076 12038 20128 12044
rect 19720 11920 19840 11948
rect 19720 11472 19748 11920
rect 19984 11824 20036 11830
rect 19984 11766 20036 11772
rect 19996 11608 20024 11766
rect 19996 11580 20116 11608
rect 19720 11444 19840 11472
rect 19156 11348 19208 11354
rect 19076 11308 19156 11336
rect 19076 11064 19104 11308
rect 19812 11336 19840 11444
rect 19812 11308 19932 11336
rect 19156 11290 19208 11296
rect 19200 11180 19820 11200
rect 19200 11124 19242 11180
rect 19298 11124 19322 11180
rect 19378 11124 19402 11180
rect 19458 11124 19482 11180
rect 19538 11124 19562 11180
rect 19618 11124 19642 11180
rect 19698 11124 19722 11180
rect 19778 11124 19820 11180
rect 19200 11104 19820 11124
rect 19904 11064 19932 11308
rect 20088 11132 20116 11580
rect 19076 11036 19196 11064
rect 19168 10928 19196 11036
rect 19812 11036 19932 11064
rect 19996 11104 20116 11132
rect 20364 11336 20392 13076
rect 20444 13058 20496 13064
rect 20548 12981 20576 13194
rect 20810 13151 20866 13160
rect 21270 13216 21326 13225
rect 21270 13151 21326 13160
rect 20534 12972 20590 12981
rect 20534 12907 20590 12916
rect 20440 12812 21060 12832
rect 20440 12756 20482 12812
rect 20538 12756 20562 12812
rect 20618 12756 20642 12812
rect 20698 12756 20722 12812
rect 20778 12756 20802 12812
rect 20858 12756 20882 12812
rect 20938 12756 20962 12812
rect 21018 12756 21060 12812
rect 20440 12736 21060 12756
rect 21088 12504 21140 12510
rect 21086 12484 21088 12493
rect 21140 12484 21142 12493
rect 21086 12419 21142 12428
rect 21180 12028 21232 12034
rect 21178 11996 21180 12005
rect 21232 11996 21234 12005
rect 21178 11931 21234 11940
rect 21284 11880 21312 13151
rect 21468 13054 21496 14146
rect 21744 13920 21772 15574
rect 21928 14346 21956 15642
rect 21916 14340 21968 14346
rect 22112 14323 22140 15660
rect 22296 15230 22324 16254
rect 22756 15842 22784 17410
rect 23032 16504 23060 18312
rect 26436 18154 26464 22667
rect 26424 18148 26476 18154
rect 26424 18090 26476 18096
rect 23480 16924 23532 16930
rect 23480 16866 23532 16872
rect 22940 16476 23060 16504
rect 22940 16318 22968 16476
rect 22928 16312 22980 16318
rect 22928 16254 22980 16260
rect 22744 15836 22796 15842
rect 22744 15778 22796 15784
rect 22284 15224 22336 15230
rect 22284 15166 22336 15172
rect 21916 14282 21968 14288
rect 22098 14314 22154 14323
rect 22098 14249 22154 14258
rect 21744 13892 21956 13920
rect 21732 13796 21784 13802
rect 21732 13738 21784 13744
rect 21744 13258 21772 13738
rect 21732 13252 21784 13258
rect 21732 13194 21784 13200
rect 21640 13184 21692 13190
rect 21640 13126 21692 13132
rect 21456 13048 21508 13054
rect 21456 12990 21508 12996
rect 21468 11966 21496 12990
rect 21652 12714 21680 13126
rect 21824 13116 21876 13122
rect 21824 13058 21876 13064
rect 21640 12708 21692 12714
rect 21836 12696 21864 13058
rect 21640 12650 21692 12656
rect 21790 12668 21864 12696
rect 21640 12436 21692 12442
rect 21640 12378 21692 12384
rect 21652 12170 21680 12378
rect 21640 12164 21692 12170
rect 21640 12106 21692 12112
rect 21790 12016 21818 12668
rect 21744 11988 21818 12016
rect 21456 11960 21508 11966
rect 21456 11902 21508 11908
rect 21192 11852 21312 11880
rect 20440 11724 21060 11744
rect 20440 11668 20482 11724
rect 20538 11668 20562 11724
rect 20618 11668 20642 11724
rect 20698 11668 20722 11724
rect 20778 11668 20802 11724
rect 20858 11668 20882 11724
rect 20938 11668 20962 11724
rect 21018 11668 21060 11724
rect 20440 11648 21060 11668
rect 21192 11422 21220 11852
rect 21180 11416 21232 11422
rect 21180 11358 21232 11364
rect 20444 11348 20496 11354
rect 20364 11308 20444 11336
rect 19812 10928 19840 11036
rect 19168 10900 19288 10928
rect 19260 10384 19288 10900
rect 19168 10356 19288 10384
rect 19720 10900 19840 10928
rect 19720 10384 19748 10900
rect 19720 10356 19840 10384
rect 19168 10248 19196 10356
rect 19076 10220 19196 10248
rect 19812 10248 19840 10356
rect 19812 10220 19932 10248
rect 19076 8820 19104 10220
rect 19200 10092 19820 10112
rect 19200 10036 19242 10092
rect 19298 10036 19322 10092
rect 19378 10036 19402 10092
rect 19458 10036 19482 10092
rect 19538 10036 19562 10092
rect 19618 10036 19642 10092
rect 19698 10036 19722 10092
rect 19778 10036 19820 10092
rect 19200 10016 19820 10036
rect 19904 9976 19932 10220
rect 19812 9948 19932 9976
rect 19340 9852 19392 9858
rect 19812 9840 19840 9948
rect 19340 9794 19392 9800
rect 19720 9812 19840 9840
rect 19156 9716 19208 9722
rect 19154 9678 19156 9687
rect 19208 9678 19210 9687
rect 19154 9613 19210 9622
rect 19352 9104 19380 9794
rect 19720 9364 19748 9812
rect 19996 9382 20024 11104
rect 20168 10940 20220 10946
rect 20168 10882 20220 10888
rect 20180 10520 20208 10882
rect 20260 10532 20312 10538
rect 20180 10492 20260 10520
rect 20260 10474 20312 10480
rect 20364 10334 20392 11308
rect 20444 11290 20496 11296
rect 20536 11348 20588 11354
rect 20536 11290 20588 11296
rect 20812 11348 20864 11354
rect 20812 11290 20864 11296
rect 20548 10736 20576 11290
rect 20824 11082 20852 11290
rect 20812 11076 20864 11082
rect 21192 11064 21220 11358
rect 21364 11280 21416 11286
rect 21364 11222 21416 11228
rect 21192 11036 21312 11064
rect 20812 11018 20864 11024
rect 21088 11008 21140 11014
rect 21088 10950 21140 10956
rect 20530 10684 20536 10736
rect 20588 10684 20594 10736
rect 20440 10636 21060 10656
rect 20440 10580 20482 10636
rect 20538 10580 20562 10636
rect 20618 10580 20642 10636
rect 20698 10580 20722 10636
rect 20778 10580 20802 10636
rect 20858 10580 20882 10636
rect 20938 10580 20962 10636
rect 21018 10580 21060 10636
rect 20440 10560 21060 10580
rect 20352 10328 20404 10334
rect 20350 10288 20352 10297
rect 20628 10328 20680 10334
rect 20404 10288 20406 10297
rect 20628 10270 20680 10276
rect 20350 10223 20406 10232
rect 20168 9852 20220 9858
rect 20168 9794 20220 9800
rect 20180 9450 20208 9794
rect 20168 9444 20220 9450
rect 20168 9386 20220 9392
rect 19984 9376 20036 9382
rect 19720 9336 19840 9364
rect 19812 9178 19840 9336
rect 19984 9318 20036 9324
rect 20166 9312 20222 9321
rect 20166 9247 20222 9256
rect 19800 9172 19852 9178
rect 19800 9114 19852 9120
rect 19984 9172 20036 9178
rect 19984 9114 20036 9120
rect 19334 9052 19340 9104
rect 19392 9052 19398 9104
rect 19200 9004 19820 9024
rect 19200 8948 19242 9004
rect 19298 8948 19322 9004
rect 19378 8948 19402 9004
rect 19458 8948 19482 9004
rect 19538 8948 19562 9004
rect 19618 8948 19642 9004
rect 19698 8948 19722 9004
rect 19778 8948 19820 9004
rect 19200 8928 19820 8948
rect 19996 8820 20024 9114
rect 20180 8906 20208 9247
rect 20364 9246 20392 10223
rect 20640 9994 20668 10270
rect 20812 10192 20864 10198
rect 20812 10134 20864 10140
rect 20628 9988 20680 9994
rect 20628 9930 20680 9936
rect 20824 9858 20852 10134
rect 20812 9852 20864 9858
rect 20812 9794 20864 9800
rect 20440 9548 21060 9568
rect 20440 9492 20482 9548
rect 20538 9492 20562 9548
rect 20618 9492 20642 9548
rect 20698 9492 20722 9548
rect 20778 9492 20802 9548
rect 20858 9492 20882 9548
rect 20938 9492 20962 9548
rect 21018 9492 21060 9548
rect 20440 9472 21060 9492
rect 21100 9364 21128 10950
rect 21284 10402 21312 11036
rect 21376 11014 21404 11222
rect 21364 11008 21416 11014
rect 21364 10950 21416 10956
rect 21468 10878 21496 11902
rect 21744 11830 21772 11988
rect 21732 11824 21784 11830
rect 21732 11766 21784 11772
rect 21744 11608 21772 11766
rect 21744 11580 21818 11608
rect 21640 11552 21692 11558
rect 21640 11494 21692 11500
rect 21456 10872 21508 10878
rect 21456 10814 21508 10820
rect 21272 10396 21324 10402
rect 21272 10338 21324 10344
rect 21008 9336 21128 9364
rect 20352 9240 20404 9246
rect 21008 9228 21036 9336
rect 21284 9296 21312 10338
rect 21468 10334 21496 10814
rect 21456 10328 21508 10334
rect 21456 10270 21508 10276
rect 21468 9931 21496 10270
rect 21652 10248 21680 11494
rect 21790 10384 21818 11580
rect 21928 10878 21956 13892
rect 22006 13216 22062 13225
rect 22006 13151 22062 13160
rect 22020 13122 22048 13151
rect 22008 13116 22060 13122
rect 22008 13058 22060 13064
rect 22112 12220 22140 14249
rect 22296 14210 22324 15166
rect 22468 15088 22520 15094
rect 22468 15030 22520 15036
rect 22480 14686 22508 15030
rect 22756 14748 22784 15778
rect 22926 15290 22982 15299
rect 22926 15225 22982 15234
rect 22940 15076 22968 15225
rect 22940 15048 23060 15076
rect 22738 14696 22744 14748
rect 22796 14696 22802 14748
rect 22468 14680 22520 14686
rect 22468 14622 22520 14628
rect 22284 14204 22336 14210
rect 22284 14146 22336 14152
rect 22066 12192 22140 12220
rect 22066 11676 22094 12192
rect 22296 12152 22324 14146
rect 22756 13660 22784 14696
rect 23032 14192 23060 15048
rect 22940 14164 23060 14192
rect 22940 14006 22968 14164
rect 22928 14000 22980 14006
rect 22928 13942 22980 13948
rect 22738 13608 22744 13660
rect 22796 13608 22802 13660
rect 22468 13592 22520 13598
rect 22468 13534 22520 13540
rect 22204 12124 22324 12152
rect 22204 11966 22232 12124
rect 22192 11960 22244 11966
rect 22192 11902 22244 11908
rect 22204 11744 22232 11902
rect 22204 11716 22324 11744
rect 22066 11648 22140 11676
rect 21916 10872 21968 10878
rect 21916 10814 21968 10820
rect 21790 10356 21864 10384
rect 21836 10297 21864 10356
rect 21822 10288 21878 10297
rect 21652 10220 21772 10248
rect 21928 10266 21956 10814
rect 21822 10223 21878 10232
rect 21916 10260 21968 10266
rect 21454 9922 21510 9931
rect 21454 9857 21510 9866
rect 20352 9182 20404 9188
rect 20916 9200 21036 9228
rect 21192 9268 21312 9296
rect 20168 8900 20220 8906
rect 20168 8842 20220 8848
rect 19076 8792 19196 8820
rect 18972 8356 19024 8362
rect 19168 8344 19196 8792
rect 18972 8298 19024 8304
rect 19076 8316 19196 8344
rect 19904 8792 20024 8820
rect 19076 8158 19104 8316
rect 19904 8208 19932 8792
rect 20260 8696 20312 8702
rect 20260 8638 20312 8644
rect 20168 8628 20220 8634
rect 20272 8589 20300 8638
rect 20168 8570 20220 8576
rect 20258 8580 20314 8589
rect 19904 8180 20116 8208
rect 19064 8152 19116 8158
rect 19064 8094 19116 8100
rect 19984 8084 20036 8090
rect 19984 8026 20036 8032
rect 19200 7916 19820 7936
rect 19200 7860 19242 7916
rect 19298 7860 19322 7916
rect 19378 7860 19402 7916
rect 19458 7860 19482 7916
rect 19538 7860 19562 7916
rect 19618 7860 19642 7916
rect 19698 7860 19722 7916
rect 19778 7860 19820 7916
rect 19200 7840 19820 7860
rect 18972 7812 19024 7818
rect 18972 7754 19024 7760
rect 18786 7726 18842 7735
rect 18328 7676 18380 7682
rect 18328 7618 18380 7624
rect 18604 7676 18656 7682
rect 18786 7661 18842 7670
rect 18604 7618 18656 7624
rect 18052 7608 18104 7614
rect 18052 7550 18104 7556
rect 18144 7472 18196 7478
rect 16868 7432 16988 7460
rect 17788 7432 17908 7460
rect 16960 7274 16988 7432
rect 17880 7274 17908 7432
rect 18144 7414 18196 7420
rect 16948 7268 17000 7274
rect 16948 7210 17000 7216
rect 17868 7268 17920 7274
rect 17868 7210 17920 7216
rect 17776 7064 17828 7070
rect 18156 7052 18184 7414
rect 17776 7006 17828 7012
rect 18064 7024 18184 7052
rect 16408 6140 16896 6168
rect 16212 6112 16264 6118
rect 16212 6054 16264 6060
rect 14280 6044 14332 6050
rect 16868 6027 16896 6140
rect 14280 5986 14332 5992
rect 16854 6018 16910 6027
rect 17788 5982 17816 7006
rect 18064 6440 18092 7024
rect 18340 6594 18368 7618
rect 18616 7003 18644 7618
rect 18984 7268 19012 7754
rect 19246 7726 19302 7735
rect 19246 7661 19302 7670
rect 19798 7726 19854 7735
rect 19996 7682 20024 8026
rect 19798 7661 19854 7670
rect 19984 7676 20036 7682
rect 18966 7216 18972 7268
rect 19024 7216 19030 7268
rect 19260 7138 19288 7661
rect 19812 7546 19840 7661
rect 19984 7618 20036 7624
rect 19800 7540 19852 7546
rect 19800 7482 19852 7488
rect 19248 7132 19300 7138
rect 19248 7074 19300 7080
rect 18602 6994 18658 7003
rect 18602 6929 18658 6938
rect 18328 6588 18380 6594
rect 18328 6530 18380 6536
rect 18616 6526 18644 6929
rect 18972 6928 19024 6934
rect 18972 6870 19024 6876
rect 18604 6520 18656 6526
rect 18604 6462 18656 6468
rect 18786 6506 18842 6515
rect 18786 6441 18842 6450
rect 18064 6412 18184 6440
rect 18156 6050 18184 6412
rect 18800 6186 18828 6441
rect 18984 6186 19012 6870
rect 19200 6828 19820 6848
rect 19200 6772 19242 6828
rect 19298 6772 19322 6828
rect 19378 6772 19402 6828
rect 19458 6772 19482 6828
rect 19538 6772 19562 6828
rect 19618 6772 19642 6828
rect 19698 6772 19722 6828
rect 19778 6772 19820 6828
rect 19200 6752 19820 6772
rect 19800 6520 19852 6526
rect 19800 6462 19852 6468
rect 19812 6186 19840 6462
rect 18788 6180 18840 6186
rect 18788 6122 18840 6128
rect 18972 6180 19024 6186
rect 18972 6122 19024 6128
rect 19800 6180 19852 6186
rect 19800 6122 19852 6128
rect 20088 6050 20116 8180
rect 20180 7750 20208 8570
rect 20258 8515 20314 8524
rect 20364 8158 20392 9182
rect 20916 8752 20944 9200
rect 21192 9110 21220 9268
rect 21180 9104 21232 9110
rect 21180 9046 21232 9052
rect 20916 8724 21036 8752
rect 21008 8616 21036 8724
rect 21008 8588 21128 8616
rect 20440 8460 21060 8480
rect 20440 8404 20482 8460
rect 20538 8404 20562 8460
rect 20618 8404 20642 8460
rect 20698 8404 20722 8460
rect 20778 8404 20802 8460
rect 20858 8404 20882 8460
rect 20938 8404 20962 8460
rect 21018 8404 21060 8460
rect 20440 8384 21060 8404
rect 21100 8276 21128 8588
rect 21192 8362 21220 9046
rect 21180 8356 21232 8362
rect 21180 8298 21232 8304
rect 21270 8336 21326 8345
rect 21008 8248 21128 8276
rect 21270 8271 21326 8280
rect 20352 8152 20404 8158
rect 20536 8152 20588 8158
rect 20352 8094 20404 8100
rect 20534 8100 20536 8101
rect 20588 8100 20590 8101
rect 20534 8092 20590 8100
rect 20534 8027 20590 8036
rect 20720 8084 20772 8090
rect 20720 8026 20772 8032
rect 20168 7744 20220 7750
rect 20168 7686 20220 7692
rect 20260 7608 20312 7614
rect 20260 7550 20312 7556
rect 20272 7274 20300 7550
rect 20732 7528 20760 8026
rect 20364 7500 20760 7528
rect 21008 7528 21036 8248
rect 21008 7500 21128 7528
rect 20260 7268 20312 7274
rect 20260 7210 20312 7216
rect 18144 6044 18196 6050
rect 18144 5986 18196 5992
rect 20076 6044 20128 6050
rect 20076 5986 20128 5992
rect 20364 5982 20392 7500
rect 20440 7372 21060 7392
rect 20440 7316 20482 7372
rect 20538 7316 20562 7372
rect 20618 7316 20642 7372
rect 20698 7316 20722 7372
rect 20778 7316 20802 7372
rect 20858 7316 20882 7372
rect 20938 7316 20962 7372
rect 21018 7316 21060 7372
rect 20440 7296 21060 7316
rect 21100 7256 21128 7500
rect 21008 7228 21128 7256
rect 20720 7132 20772 7138
rect 20720 7074 20772 7080
rect 20732 6730 20760 7074
rect 20720 6724 20772 6730
rect 20720 6666 20772 6672
rect 21008 6594 21036 7228
rect 20996 6588 21048 6594
rect 20996 6530 21048 6536
rect 20440 6284 21060 6304
rect 20440 6228 20482 6284
rect 20538 6228 20562 6284
rect 20618 6228 20642 6284
rect 20698 6228 20722 6284
rect 20778 6228 20802 6284
rect 20858 6228 20882 6284
rect 20938 6228 20962 6284
rect 21018 6228 21060 6284
rect 20440 6208 21060 6228
rect 21284 6050 21312 8271
rect 21468 8158 21496 9857
rect 21744 9840 21772 10220
rect 21916 10202 21968 10208
rect 22112 10044 22140 11648
rect 22296 10044 22324 11716
rect 22480 11268 22508 13534
rect 22756 12493 22784 13608
rect 22928 12708 22980 12714
rect 22928 12650 22980 12656
rect 22742 12484 22798 12493
rect 22940 12492 22968 12650
rect 22940 12464 23060 12492
rect 22742 12419 22798 12428
rect 22756 11490 22784 12419
rect 22744 11484 22796 11490
rect 22744 11426 22796 11432
rect 23032 11336 23060 12464
rect 22940 11308 23060 11336
rect 22480 11240 22600 11268
rect 22572 10384 22600 11240
rect 22020 10016 22140 10044
rect 22204 10016 22324 10044
rect 22480 10356 22600 10384
rect 21744 9812 21864 9840
rect 21640 9716 21692 9722
rect 21640 9658 21692 9664
rect 21652 9450 21680 9658
rect 21640 9444 21692 9450
rect 21640 9386 21692 9392
rect 21836 9296 21864 9812
rect 22020 9500 22048 10016
rect 22204 9858 22232 10016
rect 22480 9994 22508 10356
rect 22744 10192 22796 10198
rect 22744 10134 22796 10140
rect 22468 9988 22520 9994
rect 22468 9930 22520 9936
rect 22192 9852 22244 9858
rect 22244 9812 22324 9840
rect 22192 9794 22244 9800
rect 22192 9716 22244 9722
rect 22192 9658 22244 9664
rect 22020 9472 22140 9500
rect 22112 9314 22140 9472
rect 21652 9268 21864 9296
rect 22100 9308 22152 9314
rect 21456 8152 21508 8158
rect 21456 8094 21508 8100
rect 21652 8090 21680 9268
rect 22100 9250 22152 9256
rect 22008 9172 22060 9178
rect 22008 9114 22060 9120
rect 21824 9104 21876 9110
rect 21824 9046 21876 9052
rect 21640 8084 21692 8090
rect 21640 8026 21692 8032
rect 21362 7726 21418 7735
rect 21362 7661 21418 7670
rect 21376 7138 21404 7661
rect 21548 7608 21600 7614
rect 21548 7550 21600 7556
rect 21560 7274 21588 7550
rect 21548 7268 21600 7274
rect 21548 7210 21600 7216
rect 21364 7132 21416 7138
rect 21364 7074 21416 7080
rect 21640 6996 21692 7002
rect 21640 6938 21692 6944
rect 21652 6515 21680 6938
rect 21836 6594 21864 9046
rect 22020 7735 22048 9114
rect 22006 7726 22062 7735
rect 22006 7661 22062 7670
rect 22008 7540 22060 7546
rect 22008 7482 22060 7488
rect 21824 6588 21876 6594
rect 21824 6530 21876 6536
rect 21638 6506 21694 6515
rect 21638 6441 21694 6450
rect 21824 6384 21876 6390
rect 21824 6326 21876 6332
rect 21836 6050 21864 6326
rect 22020 6186 22048 7482
rect 22008 6180 22060 6186
rect 22008 6122 22060 6128
rect 22204 6118 22232 9658
rect 22296 9432 22324 9812
rect 22296 9404 22508 9432
rect 22480 7868 22508 9404
rect 22756 8101 22784 10134
rect 22742 8092 22798 8101
rect 22742 8027 22798 8036
rect 22388 7840 22508 7868
rect 22388 7682 22416 7840
rect 22376 7676 22428 7682
rect 22376 7618 22428 7624
rect 22468 6928 22520 6934
rect 22468 6870 22520 6876
rect 22480 6271 22508 6870
rect 22940 6662 22968 11308
rect 23204 10328 23256 10334
rect 23204 10270 23256 10276
rect 23216 8362 23244 10270
rect 23388 9444 23440 9450
rect 23492 9432 23520 16866
rect 28736 12374 28764 27744
rect 28724 12368 28776 12374
rect 28724 12310 28776 12316
rect 26240 10736 26292 10742
rect 26240 10678 26292 10684
rect 23440 9404 23520 9432
rect 23388 9386 23440 9392
rect 23204 8356 23256 8362
rect 23204 8298 23256 8304
rect 22928 6656 22980 6662
rect 22928 6598 22980 6604
rect 22466 6262 22522 6271
rect 22466 6197 22522 6206
rect 22192 6112 22244 6118
rect 22192 6054 22244 6060
rect 21272 6044 21324 6050
rect 21272 5986 21324 5992
rect 21824 6044 21876 6050
rect 21824 5986 21876 5992
rect 16854 5953 16856 5962
rect 16908 5953 16910 5962
rect 17776 5976 17828 5982
rect 16856 5918 16908 5924
rect 17776 5918 17828 5924
rect 20352 5976 20404 5982
rect 20352 5918 20404 5924
rect 14096 5908 14148 5914
rect 14148 5868 14320 5896
rect 14096 5850 14148 5856
rect 13600 5740 14220 5760
rect 13600 5684 13642 5740
rect 13698 5684 13722 5740
rect 13778 5684 13802 5740
rect 13858 5684 13882 5740
rect 13938 5684 13962 5740
rect 14018 5684 14042 5740
rect 14098 5684 14122 5740
rect 14178 5684 14220 5740
rect 13600 5664 14220 5684
rect 13452 196 13504 202
rect 14292 171 14320 5868
rect 19200 5740 19820 5760
rect 19200 5684 19242 5740
rect 19298 5684 19322 5740
rect 19378 5684 19402 5740
rect 19458 5684 19482 5740
rect 19538 5684 19562 5740
rect 19618 5684 19642 5740
rect 19698 5684 19722 5740
rect 19778 5684 19820 5740
rect 19200 5664 19820 5684
rect 23216 5295 23244 8298
rect 23202 5286 23258 5295
rect 23202 5221 23258 5230
rect 19156 4140 19208 4146
rect 19156 4082 19208 4088
rect 13452 138 13504 144
rect 14278 162 14334 171
rect 14278 97 14334 106
rect 19168 0 19196 4082
rect 26252 2733 26280 10678
rect 28538 8092 28594 8101
rect 28538 8027 28594 8036
rect 26238 2724 26294 2733
rect 26238 2659 26294 2668
rect 28552 171 28580 8027
rect 28722 406 28778 415
rect 28722 341 28778 350
rect 28538 162 28594 171
rect 28538 97 28594 106
rect 28736 0 28764 341
<< via2 >>
rect 18602 27678 18658 27734
rect 8042 22004 8098 22060
rect 8122 22004 8178 22060
rect 8202 22004 8258 22060
rect 8282 22004 8338 22060
rect 8362 22004 8418 22060
rect 8442 22004 8498 22060
rect 8522 22004 8578 22060
rect 13642 22004 13698 22060
rect 13722 22004 13778 22060
rect 13802 22004 13858 22060
rect 13882 22004 13938 22060
rect 13962 22004 14018 22060
rect 14042 22004 14098 22060
rect 14122 22004 14178 22060
rect 21822 25238 21878 25294
rect 19242 22004 19298 22060
rect 19322 22004 19378 22060
rect 19402 22004 19458 22060
rect 19482 22004 19538 22060
rect 19562 22004 19618 22060
rect 19642 22004 19698 22060
rect 19722 22004 19778 22060
rect 20350 21822 20406 21878
rect 9282 21460 9338 21516
rect 9362 21460 9418 21516
rect 9442 21460 9498 21516
rect 9522 21460 9578 21516
rect 9602 21460 9658 21516
rect 9682 21460 9738 21516
rect 9762 21460 9818 21516
rect 8042 20916 8098 20972
rect 8122 20916 8178 20972
rect 8202 20916 8258 20972
rect 8282 20916 8338 20972
rect 8362 20916 8418 20972
rect 8442 20916 8498 20972
rect 8522 20916 8578 20972
rect 8042 19828 8098 19884
rect 8122 19828 8178 19884
rect 8202 19828 8258 19884
rect 8282 19828 8338 19884
rect 8362 19828 8418 19884
rect 8442 19828 8498 19884
rect 8522 19828 8578 19884
rect 9282 20372 9338 20428
rect 9362 20372 9418 20428
rect 9442 20372 9498 20428
rect 9522 20372 9578 20428
rect 9602 20372 9658 20428
rect 9682 20372 9738 20428
rect 9762 20372 9818 20428
rect 8042 18740 8098 18796
rect 8122 18740 8178 18796
rect 8202 18740 8258 18796
rect 8282 18740 8338 18796
rect 8362 18740 8418 18796
rect 8442 18740 8498 18796
rect 8522 18740 8578 18796
rect 9282 19284 9338 19340
rect 9362 19284 9418 19340
rect 9442 19284 9498 19340
rect 9522 19284 9578 19340
rect 9602 19284 9658 19340
rect 9682 19284 9738 19340
rect 9762 19284 9818 19340
rect 8042 17652 8098 17708
rect 8122 17652 8178 17708
rect 8202 17652 8258 17708
rect 8282 17652 8338 17708
rect 8362 17652 8418 17708
rect 8442 17652 8498 17708
rect 8522 17652 8578 17708
rect 9282 18196 9338 18252
rect 9362 18196 9418 18252
rect 9442 18196 9498 18252
rect 9522 18196 9578 18252
rect 9602 18196 9658 18252
rect 9682 18196 9738 18252
rect 9762 18196 9818 18252
rect 14882 21460 14938 21516
rect 14962 21460 15018 21516
rect 15042 21460 15098 21516
rect 15122 21460 15178 21516
rect 15202 21460 15258 21516
rect 15282 21460 15338 21516
rect 15362 21460 15418 21516
rect 13642 20916 13698 20972
rect 13722 20916 13778 20972
rect 13802 20916 13858 20972
rect 13882 20916 13938 20972
rect 13962 20916 14018 20972
rect 14042 20916 14098 20972
rect 14122 20916 14178 20972
rect 13642 19828 13698 19884
rect 13722 19828 13778 19884
rect 13802 19828 13858 19884
rect 13882 19828 13938 19884
rect 13962 19828 14018 19884
rect 14042 19828 14098 19884
rect 14122 19828 14178 19884
rect 8042 16564 8098 16620
rect 8122 16564 8178 16620
rect 8202 16564 8258 16620
rect 8282 16564 8338 16620
rect 8362 16564 8418 16620
rect 8442 16564 8498 16620
rect 8522 16564 8578 16620
rect 7102 15966 7158 16022
rect 7470 15966 7526 16022
rect 9282 17108 9338 17164
rect 9362 17108 9418 17164
rect 9442 17108 9498 17164
rect 9522 17108 9578 17164
rect 9602 17108 9658 17164
rect 9682 17108 9738 17164
rect 9762 17108 9818 17164
rect 7286 15722 7342 15778
rect 8666 15722 8722 15778
rect 8042 15476 8098 15532
rect 8122 15476 8178 15532
rect 8202 15476 8258 15532
rect 8282 15476 8338 15532
rect 8362 15476 8418 15532
rect 8442 15476 8498 15532
rect 8522 15476 8578 15532
rect 9282 16020 9338 16076
rect 9362 16020 9418 16076
rect 9442 16020 9498 16076
rect 9522 16020 9578 16076
rect 9602 16020 9658 16076
rect 9682 16020 9738 16076
rect 9762 16020 9818 16076
rect 14882 20372 14938 20428
rect 14962 20372 15018 20428
rect 15042 20372 15098 20428
rect 15122 20372 15178 20428
rect 15202 20372 15258 20428
rect 15282 20372 15338 20428
rect 15362 20372 15418 20428
rect 15934 20120 15990 20170
rect 15934 20114 15936 20120
rect 15936 20114 15988 20120
rect 15988 20114 15990 20120
rect 14882 19284 14938 19340
rect 14962 19284 15018 19340
rect 15042 19284 15098 19340
rect 15122 19284 15178 19340
rect 15202 19284 15258 19340
rect 15282 19284 15338 19340
rect 15362 19284 15418 19340
rect 13642 18740 13698 18796
rect 13722 18740 13778 18796
rect 13802 18740 13858 18796
rect 13882 18740 13938 18796
rect 13962 18740 14018 18796
rect 14042 18740 14098 18796
rect 14122 18740 14178 18796
rect 9494 15768 9550 15778
rect 9494 15722 9496 15768
rect 9496 15722 9548 15768
rect 9548 15722 9550 15768
rect 9282 14932 9338 14988
rect 9362 14932 9418 14988
rect 9442 14932 9498 14988
rect 9522 14932 9578 14988
rect 9602 14932 9658 14988
rect 9682 14932 9738 14988
rect 9762 14932 9818 14988
rect 18 14746 74 14802
rect 5814 13770 5870 13826
rect 8042 14388 8098 14444
rect 8122 14388 8178 14444
rect 8202 14388 8258 14444
rect 8282 14388 8338 14444
rect 8362 14388 8418 14444
rect 8442 14388 8498 14444
rect 8522 14388 8578 14444
rect 9282 13844 9338 13900
rect 9362 13844 9418 13900
rect 9442 13844 9498 13900
rect 9522 13844 9578 13900
rect 9602 13844 9658 13900
rect 9682 13844 9738 13900
rect 9762 13844 9818 13900
rect 8042 13300 8098 13356
rect 8122 13300 8178 13356
rect 8202 13300 8258 13356
rect 8282 13300 8338 13356
rect 8362 13300 8418 13356
rect 8442 13300 8498 13356
rect 8522 13300 8578 13356
rect 10690 15722 10746 15778
rect 10598 14746 10654 14802
rect 9282 12756 9338 12812
rect 9362 12756 9418 12812
rect 9442 12756 9498 12812
rect 9522 12756 9578 12812
rect 9602 12756 9658 12812
rect 9682 12756 9738 12812
rect 9762 12756 9818 12812
rect 8042 12212 8098 12268
rect 8122 12212 8178 12268
rect 8202 12212 8258 12268
rect 8282 12212 8338 12268
rect 8362 12212 8418 12268
rect 8442 12212 8498 12268
rect 8522 12212 8578 12268
rect 9282 11668 9338 11724
rect 9362 11668 9418 11724
rect 9442 11668 9498 11724
rect 9522 11668 9578 11724
rect 9602 11668 9658 11724
rect 9682 11668 9738 11724
rect 9762 11668 9818 11724
rect 8042 11124 8098 11180
rect 8122 11124 8178 11180
rect 8202 11124 8258 11180
rect 8282 11124 8338 11180
rect 8362 11124 8418 11180
rect 8442 11124 8498 11180
rect 8522 11124 8578 11180
rect 8042 10036 8098 10092
rect 8122 10036 8178 10092
rect 8202 10036 8258 10092
rect 8282 10036 8338 10092
rect 8362 10036 8418 10092
rect 8442 10036 8498 10092
rect 8522 10036 8578 10092
rect 9282 10580 9338 10636
rect 9362 10580 9418 10636
rect 9442 10580 9498 10636
rect 9522 10580 9578 10636
rect 9602 10580 9658 10636
rect 9682 10580 9738 10636
rect 9762 10580 9818 10636
rect 10046 10232 10102 10288
rect 9282 9492 9338 9548
rect 9362 9492 9418 9548
rect 9442 9492 9498 9548
rect 9522 9492 9578 9548
rect 9602 9492 9658 9548
rect 9682 9492 9738 9548
rect 9762 9492 9818 9548
rect 8042 8948 8098 9004
rect 8122 8948 8178 9004
rect 8202 8948 8258 9004
rect 8282 8948 8338 9004
rect 8362 8948 8418 9004
rect 8442 8948 8498 9004
rect 8522 8948 8578 9004
rect 7286 6572 7342 6628
rect 8042 7860 8098 7916
rect 8122 7860 8178 7916
rect 8202 7860 8258 7916
rect 8282 7860 8338 7916
rect 8362 7860 8418 7916
rect 8442 7860 8498 7916
rect 8522 7860 8578 7916
rect 9282 8404 9338 8460
rect 9362 8404 9418 8460
rect 9442 8404 9498 8460
rect 9522 8404 9578 8460
rect 9602 8404 9658 8460
rect 9682 8404 9738 8460
rect 9762 8404 9818 8460
rect 16854 19138 16910 19194
rect 13642 17652 13698 17708
rect 13722 17652 13778 17708
rect 13802 17652 13858 17708
rect 13882 17652 13938 17708
rect 13962 17652 14018 17708
rect 14042 17652 14098 17708
rect 14122 17652 14178 17708
rect 14278 17430 14334 17486
rect 14882 18196 14938 18252
rect 14962 18196 15018 18252
rect 15042 18196 15098 18252
rect 15122 18196 15178 18252
rect 15202 18196 15258 18252
rect 15282 18196 15338 18252
rect 15362 18196 15418 18252
rect 19242 20916 19298 20972
rect 19322 20916 19378 20972
rect 19402 20916 19458 20972
rect 19482 20916 19538 20972
rect 19562 20916 19618 20972
rect 19642 20916 19698 20972
rect 19722 20916 19778 20972
rect 20482 21460 20538 21516
rect 20562 21460 20618 21516
rect 20642 21460 20698 21516
rect 20722 21460 20778 21516
rect 20802 21460 20858 21516
rect 20882 21460 20938 21516
rect 20962 21460 21018 21516
rect 19154 20114 19210 20170
rect 20074 20120 20130 20170
rect 20074 20114 20076 20120
rect 20076 20114 20128 20120
rect 20128 20114 20130 20120
rect 20482 20372 20538 20428
rect 20562 20372 20618 20428
rect 20642 20372 20698 20428
rect 20722 20372 20778 20428
rect 20802 20372 20858 20428
rect 20882 20372 20938 20428
rect 20962 20372 21018 20428
rect 19242 19828 19298 19884
rect 19322 19828 19378 19884
rect 19402 19828 19458 19884
rect 19482 19828 19538 19884
rect 19562 19828 19618 19884
rect 19642 19828 19698 19884
rect 19722 19828 19778 19884
rect 19062 19626 19118 19682
rect 14830 17430 14886 17486
rect 14882 17108 14938 17164
rect 14962 17108 15018 17164
rect 15042 17108 15098 17164
rect 15122 17108 15178 17164
rect 15202 17108 15258 17164
rect 15282 17108 15338 17164
rect 15362 17108 15418 17164
rect 13642 16564 13698 16620
rect 13722 16564 13778 16620
rect 13802 16564 13858 16620
rect 13882 16564 13938 16620
rect 13962 16564 14018 16620
rect 14042 16564 14098 16620
rect 14122 16564 14178 16620
rect 14882 16020 14938 16076
rect 14962 16020 15018 16076
rect 15042 16020 15098 16076
rect 15122 16020 15178 16076
rect 15202 16020 15258 16076
rect 15282 16020 15338 16076
rect 15362 16020 15418 16076
rect 13642 15476 13698 15532
rect 13722 15476 13778 15532
rect 13802 15476 13858 15532
rect 13882 15476 13938 15532
rect 13962 15476 14018 15532
rect 14042 15476 14098 15532
rect 14122 15476 14178 15532
rect 12346 12550 12402 12606
rect 15750 15844 15806 15900
rect 13642 14388 13698 14444
rect 13722 14388 13778 14444
rect 13802 14388 13858 14444
rect 13882 14388 13938 14444
rect 13962 14388 14018 14444
rect 14042 14388 14098 14444
rect 14122 14388 14178 14444
rect 14882 14932 14938 14988
rect 14962 14932 15018 14988
rect 15042 14932 15098 14988
rect 15122 14932 15178 14988
rect 15202 14932 15258 14988
rect 15282 14932 15338 14988
rect 15362 14932 15418 14988
rect 14738 14136 14794 14192
rect 15750 14152 15752 14192
rect 15752 14152 15804 14192
rect 15804 14152 15806 14192
rect 14554 13648 14610 13704
rect 13642 13300 13698 13356
rect 13722 13300 13778 13356
rect 13802 13300 13858 13356
rect 13882 13300 13938 13356
rect 13962 13300 14018 13356
rect 14042 13300 14098 13356
rect 14122 13300 14178 13356
rect 13266 12572 13322 12606
rect 13266 12550 13268 12572
rect 13268 12550 13320 12572
rect 13320 12550 13322 12572
rect 13642 12212 13698 12268
rect 13722 12212 13778 12268
rect 13802 12212 13858 12268
rect 13882 12212 13938 12268
rect 13962 12212 14018 12268
rect 14042 12212 14098 12268
rect 14122 12212 14178 12268
rect 14002 11940 14058 11996
rect 13642 11124 13698 11180
rect 13722 11124 13778 11180
rect 13802 11124 13858 11180
rect 13882 11124 13938 11180
rect 13962 11124 14018 11180
rect 14042 11124 14098 11180
rect 14122 11124 14178 11180
rect 9126 7670 9182 7726
rect 8042 6772 8098 6828
rect 8122 6772 8178 6828
rect 8202 6772 8258 6828
rect 8282 6772 8338 6828
rect 8362 6772 8418 6828
rect 8442 6772 8498 6828
rect 8522 6772 8578 6828
rect 8206 6328 8262 6384
rect 9282 7316 9338 7372
rect 9362 7316 9418 7372
rect 9442 7316 9498 7372
rect 9522 7316 9578 7372
rect 9602 7316 9658 7372
rect 9682 7316 9738 7372
rect 9762 7316 9818 7372
rect 9310 6938 9366 6994
rect 10690 7670 10746 7726
rect 10230 6572 10286 6628
rect 9282 6228 9338 6284
rect 9362 6228 9418 6284
rect 9442 6228 9498 6284
rect 9522 6228 9578 6284
rect 9602 6228 9658 6284
rect 9682 6228 9738 6284
rect 9762 6228 9818 6284
rect 8042 5684 8098 5740
rect 8122 5684 8178 5740
rect 8202 5684 8258 5740
rect 8282 5684 8338 5740
rect 8362 5684 8418 5740
rect 8442 5684 8498 5740
rect 8522 5684 8578 5740
rect 13642 10036 13698 10092
rect 13722 10036 13778 10092
rect 13802 10036 13858 10092
rect 13882 10036 13938 10092
rect 13962 10036 14018 10092
rect 14042 10036 14098 10092
rect 14122 10036 14178 10092
rect 13642 8948 13698 9004
rect 13722 8948 13778 9004
rect 13802 8948 13858 9004
rect 13882 8948 13938 9004
rect 13962 8948 14018 9004
rect 14042 8948 14098 9004
rect 14122 8948 14178 9004
rect 13450 8768 13506 8824
rect 12346 7670 12402 7726
rect 12254 5962 12310 6018
rect 13266 5976 13322 6018
rect 13266 5962 13268 5976
rect 13268 5962 13320 5976
rect 13320 5962 13322 5976
rect 13642 7860 13698 7916
rect 13722 7860 13778 7916
rect 13802 7860 13858 7916
rect 13882 7860 13938 7916
rect 13962 7860 14018 7916
rect 14042 7860 14098 7916
rect 14122 7860 14178 7916
rect 13634 7670 13690 7726
rect 13642 6772 13698 6828
rect 13722 6772 13778 6828
rect 13802 6772 13858 6828
rect 13882 6772 13938 6828
rect 13962 6772 14018 6828
rect 14042 6772 14098 6828
rect 14122 6772 14178 6828
rect 15750 14136 15806 14152
rect 14882 13844 14938 13900
rect 14962 13844 15018 13900
rect 15042 13844 15098 13900
rect 15122 13844 15178 13900
rect 15202 13844 15258 13900
rect 15282 13844 15338 13900
rect 15362 13844 15418 13900
rect 15290 13648 15346 13704
rect 15474 13160 15530 13216
rect 15290 12916 15346 12972
rect 14882 12756 14938 12812
rect 14962 12756 15018 12812
rect 15042 12756 15098 12812
rect 15122 12756 15178 12812
rect 15202 12756 15258 12812
rect 15282 12756 15338 12812
rect 15362 12756 15418 12812
rect 16210 14628 16212 14680
rect 16212 14628 16264 14680
rect 16264 14628 16266 14680
rect 16210 14624 16266 14628
rect 15842 12306 15898 12362
rect 15474 11976 15476 11996
rect 15476 11976 15528 11996
rect 15528 11976 15530 11996
rect 15474 11940 15530 11976
rect 14882 11668 14938 11724
rect 14962 11668 15018 11724
rect 15042 11668 15098 11724
rect 15122 11668 15178 11724
rect 15202 11668 15258 11724
rect 15282 11668 15338 11724
rect 15362 11668 15418 11724
rect 14882 10580 14938 10636
rect 14962 10580 15018 10636
rect 15042 10580 15098 10636
rect 15122 10580 15178 10636
rect 15202 10580 15258 10636
rect 15282 10580 15338 10636
rect 15362 10580 15418 10636
rect 15750 10354 15806 10410
rect 14882 9492 14938 9548
rect 14962 9492 15018 9548
rect 15042 9492 15098 9548
rect 15122 9492 15178 9548
rect 15202 9492 15258 9548
rect 15282 9492 15338 9548
rect 15362 9492 15418 9548
rect 15658 9378 15714 9434
rect 15474 8768 15530 8824
rect 14882 8404 14938 8460
rect 14962 8404 15018 8460
rect 15042 8404 15098 8460
rect 15122 8404 15178 8460
rect 15202 8404 15258 8460
rect 15282 8404 15338 8460
rect 15362 8404 15418 8460
rect 14646 7670 14702 7726
rect 14882 7316 14938 7372
rect 14962 7316 15018 7372
rect 15042 7316 15098 7372
rect 15122 7316 15178 7372
rect 15202 7316 15258 7372
rect 15282 7316 15338 7372
rect 15362 7316 15418 7372
rect 16670 16380 16726 16388
rect 16670 16332 16672 16380
rect 16672 16332 16724 16380
rect 16724 16332 16726 16380
rect 17314 15844 17370 15900
rect 17682 17796 17738 17852
rect 17866 17430 17922 17486
rect 16302 9622 16358 9678
rect 16762 12916 16818 12972
rect 16762 12550 16818 12606
rect 19242 18740 19298 18796
rect 19322 18740 19378 18796
rect 19402 18740 19458 18796
rect 19482 18740 19538 18796
rect 19562 18740 19618 18796
rect 19642 18740 19698 18796
rect 19722 18740 19778 18796
rect 19798 17796 19854 17852
rect 19242 17652 19298 17708
rect 19322 17652 19378 17708
rect 19402 17652 19458 17708
rect 19482 17652 19538 17708
rect 19562 17652 19618 17708
rect 19642 17652 19698 17708
rect 19722 17652 19778 17708
rect 19522 17468 19578 17486
rect 19522 17430 19524 17468
rect 19524 17430 19576 17468
rect 19576 17430 19578 17468
rect 19522 16820 19578 16876
rect 19242 16564 19298 16620
rect 19322 16564 19378 16620
rect 19402 16564 19458 16620
rect 19482 16564 19538 16620
rect 19562 16564 19618 16620
rect 19642 16564 19698 16620
rect 19722 16564 19778 16620
rect 20482 19284 20538 19340
rect 20562 19284 20618 19340
rect 20642 19284 20698 19340
rect 20722 19284 20778 19340
rect 20802 19284 20858 19340
rect 20882 19284 20938 19340
rect 20962 19284 21018 19340
rect 20482 18196 20538 18252
rect 20562 18196 20618 18252
rect 20642 18196 20698 18252
rect 20722 18196 20778 18252
rect 20802 18196 20858 18252
rect 20882 18196 20938 18252
rect 20962 18196 21018 18252
rect 20482 17108 20538 17164
rect 20562 17108 20618 17164
rect 20642 17108 20698 17164
rect 20722 17108 20778 17164
rect 20802 17108 20858 17164
rect 20882 17108 20938 17164
rect 20962 17108 21018 17164
rect 20902 16856 20958 16876
rect 20902 16820 20904 16856
rect 20904 16820 20956 16856
rect 20956 16820 20958 16856
rect 20074 16332 20130 16388
rect 18510 15112 18566 15168
rect 17958 14624 18014 14680
rect 19242 15476 19298 15532
rect 19322 15476 19378 15532
rect 19402 15476 19458 15532
rect 19482 15476 19538 15532
rect 19562 15476 19618 15532
rect 19642 15476 19698 15532
rect 19722 15476 19778 15532
rect 19062 14746 19118 14802
rect 26422 22676 26478 22732
rect 22742 21822 22798 21878
rect 22098 19138 22154 19194
rect 21638 17674 21694 17730
rect 21270 16332 21326 16388
rect 20482 16020 20538 16076
rect 20562 16020 20618 16076
rect 20642 16020 20698 16076
rect 20722 16020 20778 16076
rect 20802 16020 20858 16076
rect 20882 16020 20938 16076
rect 20962 16020 21018 16076
rect 20482 14932 20538 14988
rect 20562 14932 20618 14988
rect 20642 14932 20698 14988
rect 20722 14932 20778 14988
rect 20802 14932 20858 14988
rect 20882 14932 20938 14988
rect 20962 14932 21018 14988
rect 20626 14746 20682 14802
rect 19242 14388 19298 14444
rect 19322 14388 19378 14444
rect 19402 14388 19458 14444
rect 19482 14388 19538 14444
rect 19562 14388 19618 14444
rect 19642 14388 19698 14444
rect 19722 14388 19778 14444
rect 19062 13648 19118 13704
rect 19242 13300 19298 13356
rect 19322 13300 19378 13356
rect 19402 13300 19458 13356
rect 19482 13300 19538 13356
rect 19562 13300 19618 13356
rect 19642 13300 19698 13356
rect 19722 13300 19778 13356
rect 17498 13160 17554 13216
rect 18786 13160 18842 13216
rect 17498 12550 17554 12606
rect 18602 12550 18658 12606
rect 16854 10598 16910 10654
rect 16026 8768 16082 8824
rect 16210 8524 16266 8580
rect 16210 7670 16266 7726
rect 14882 6228 14938 6284
rect 14962 6228 15018 6284
rect 15042 6228 15098 6284
rect 15122 6228 15178 6284
rect 15202 6228 15258 6284
rect 15282 6228 15338 6284
rect 15362 6228 15418 6284
rect 17038 8524 17094 8580
rect 17130 7914 17186 7970
rect 17958 10396 18014 10410
rect 17958 10354 17960 10396
rect 17960 10354 18012 10396
rect 18012 10354 18014 10396
rect 18510 10598 18566 10654
rect 18142 10140 18144 10166
rect 18144 10140 18196 10166
rect 18196 10140 18198 10166
rect 18142 10110 18198 10140
rect 18050 9866 18106 9922
rect 18694 8768 18750 8824
rect 19242 12212 19298 12268
rect 19322 12212 19378 12268
rect 19402 12212 19458 12268
rect 19482 12212 19538 12268
rect 19562 12212 19618 12268
rect 19642 12212 19698 12268
rect 19722 12212 19778 12268
rect 20442 14502 20498 14558
rect 22742 20114 22798 20170
rect 21454 15112 21510 15168
rect 21270 14502 21326 14558
rect 21270 14258 21326 14314
rect 20482 13844 20538 13900
rect 20562 13844 20618 13900
rect 20642 13844 20698 13900
rect 20722 13844 20778 13900
rect 20802 13844 20858 13900
rect 20882 13844 20938 13900
rect 20962 13844 21018 13900
rect 20442 13648 20498 13704
rect 20166 12550 20222 12606
rect 19242 11124 19298 11180
rect 19322 11124 19378 11180
rect 19402 11124 19458 11180
rect 19482 11124 19538 11180
rect 19562 11124 19618 11180
rect 19642 11124 19698 11180
rect 19722 11124 19778 11180
rect 20810 13160 20866 13216
rect 21270 13160 21326 13216
rect 20534 12916 20590 12972
rect 20482 12756 20538 12812
rect 20562 12756 20618 12812
rect 20642 12756 20698 12812
rect 20722 12756 20778 12812
rect 20802 12756 20858 12812
rect 20882 12756 20938 12812
rect 20962 12756 21018 12812
rect 21086 12452 21088 12484
rect 21088 12452 21140 12484
rect 21140 12452 21142 12484
rect 21086 12428 21142 12452
rect 21178 11976 21180 11996
rect 21180 11976 21232 11996
rect 21232 11976 21234 11996
rect 21178 11940 21234 11976
rect 22098 14258 22154 14314
rect 20482 11668 20538 11724
rect 20562 11668 20618 11724
rect 20642 11668 20698 11724
rect 20722 11668 20778 11724
rect 20802 11668 20858 11724
rect 20882 11668 20938 11724
rect 20962 11668 21018 11724
rect 19242 10036 19298 10092
rect 19322 10036 19378 10092
rect 19402 10036 19458 10092
rect 19482 10036 19538 10092
rect 19562 10036 19618 10092
rect 19642 10036 19698 10092
rect 19722 10036 19778 10092
rect 19154 9664 19156 9678
rect 19156 9664 19208 9678
rect 19208 9664 19210 9678
rect 19154 9622 19210 9664
rect 20482 10580 20538 10636
rect 20562 10580 20618 10636
rect 20642 10580 20698 10636
rect 20722 10580 20778 10636
rect 20802 10580 20858 10636
rect 20882 10580 20938 10636
rect 20962 10580 21018 10636
rect 20350 10276 20352 10288
rect 20352 10276 20404 10288
rect 20404 10276 20406 10288
rect 20350 10232 20406 10276
rect 20166 9256 20222 9312
rect 19242 8948 19298 9004
rect 19322 8948 19378 9004
rect 19402 8948 19458 9004
rect 19482 8948 19538 9004
rect 19562 8948 19618 9004
rect 19642 8948 19698 9004
rect 19722 8948 19778 9004
rect 20482 9492 20538 9548
rect 20562 9492 20618 9548
rect 20642 9492 20698 9548
rect 20722 9492 20778 9548
rect 20802 9492 20858 9548
rect 20882 9492 20938 9548
rect 20962 9492 21018 9548
rect 22006 13160 22062 13216
rect 22926 15234 22982 15290
rect 21822 10232 21878 10288
rect 21454 9866 21510 9922
rect 19242 7860 19298 7916
rect 19322 7860 19378 7916
rect 19402 7860 19458 7916
rect 19482 7860 19538 7916
rect 19562 7860 19618 7916
rect 19642 7860 19698 7916
rect 19722 7860 19778 7916
rect 18786 7670 18842 7726
rect 16854 5976 16910 6018
rect 19246 7670 19302 7726
rect 19798 7670 19854 7726
rect 18602 6938 18658 6994
rect 18786 6450 18842 6506
rect 19242 6772 19298 6828
rect 19322 6772 19378 6828
rect 19402 6772 19458 6828
rect 19482 6772 19538 6828
rect 19562 6772 19618 6828
rect 19642 6772 19698 6828
rect 19722 6772 19778 6828
rect 20258 8524 20314 8580
rect 20482 8404 20538 8460
rect 20562 8404 20618 8460
rect 20642 8404 20698 8460
rect 20722 8404 20778 8460
rect 20802 8404 20858 8460
rect 20882 8404 20938 8460
rect 20962 8404 21018 8460
rect 21270 8280 21326 8336
rect 20534 8036 20590 8092
rect 20482 7316 20538 7372
rect 20562 7316 20618 7372
rect 20642 7316 20698 7372
rect 20722 7316 20778 7372
rect 20802 7316 20858 7372
rect 20882 7316 20938 7372
rect 20962 7316 21018 7372
rect 20482 6228 20538 6284
rect 20562 6228 20618 6284
rect 20642 6228 20698 6284
rect 20722 6228 20778 6284
rect 20802 6228 20858 6284
rect 20882 6228 20938 6284
rect 20962 6228 21018 6284
rect 22742 12428 22798 12484
rect 21362 7670 21418 7726
rect 22006 7670 22062 7726
rect 21638 6450 21694 6506
rect 22742 8036 22798 8092
rect 22466 6206 22522 6262
rect 16854 5962 16856 5976
rect 16856 5962 16908 5976
rect 16908 5962 16910 5976
rect 13642 5684 13698 5740
rect 13722 5684 13778 5740
rect 13802 5684 13858 5740
rect 13882 5684 13938 5740
rect 13962 5684 14018 5740
rect 14042 5684 14098 5740
rect 14122 5684 14178 5740
rect 19242 5684 19298 5740
rect 19322 5684 19378 5740
rect 19402 5684 19458 5740
rect 19482 5684 19538 5740
rect 19562 5684 19618 5740
rect 19642 5684 19698 5740
rect 19722 5684 19778 5740
rect 23202 5230 23258 5286
rect 14278 106 14334 162
rect 28538 8036 28594 8092
rect 26238 2668 26294 2724
rect 28722 350 28778 406
rect 28538 106 28594 162
<< metal3 >>
rect 18597 27736 18663 27739
rect 18597 27734 28796 27736
rect 18597 27678 18602 27734
rect 18658 27678 28796 27734
rect 18597 27676 28796 27678
rect 18597 27673 18663 27676
rect 21817 25296 21883 25299
rect 21817 25294 28796 25296
rect 21817 25238 21822 25294
rect 21878 25238 28796 25294
rect 21817 25236 28796 25238
rect 21817 25233 21883 25236
rect 26417 22734 26483 22737
rect 26417 22732 28796 22734
rect 26417 22676 26422 22732
rect 26478 22676 28796 22732
rect 26417 22674 28796 22676
rect 26417 22671 26483 22674
rect 8000 22064 8620 22080
rect 8000 22000 8038 22064
rect 8102 22000 8118 22064
rect 8182 22000 8198 22064
rect 8262 22000 8278 22064
rect 8342 22000 8358 22064
rect 8422 22000 8438 22064
rect 8502 22000 8518 22064
rect 8582 22000 8620 22064
rect 8000 21984 8620 22000
rect 13600 22064 14220 22080
rect 13600 22000 13638 22064
rect 13702 22000 13718 22064
rect 13782 22000 13798 22064
rect 13862 22000 13878 22064
rect 13942 22000 13958 22064
rect 14022 22000 14038 22064
rect 14102 22000 14118 22064
rect 14182 22000 14220 22064
rect 13600 21984 14220 22000
rect 19200 22064 19820 22080
rect 19200 22000 19238 22064
rect 19302 22000 19318 22064
rect 19382 22000 19398 22064
rect 19462 22000 19478 22064
rect 19542 22000 19558 22064
rect 19622 22000 19638 22064
rect 19702 22000 19718 22064
rect 19782 22000 19820 22064
rect 19200 21984 19820 22000
rect 20345 21880 20411 21883
rect 22737 21880 22803 21883
rect 20345 21878 22803 21880
rect 20345 21822 20350 21878
rect 20406 21822 22742 21878
rect 22798 21822 22803 21878
rect 20345 21820 22803 21822
rect 20345 21817 20411 21820
rect 22737 21817 22803 21820
rect 9240 21520 9860 21536
rect 9240 21456 9278 21520
rect 9342 21456 9358 21520
rect 9422 21456 9438 21520
rect 9502 21456 9518 21520
rect 9582 21456 9598 21520
rect 9662 21456 9678 21520
rect 9742 21456 9758 21520
rect 9822 21456 9860 21520
rect 9240 21440 9860 21456
rect 14840 21520 15460 21536
rect 14840 21456 14878 21520
rect 14942 21456 14958 21520
rect 15022 21456 15038 21520
rect 15102 21456 15118 21520
rect 15182 21456 15198 21520
rect 15262 21456 15278 21520
rect 15342 21456 15358 21520
rect 15422 21456 15460 21520
rect 14840 21440 15460 21456
rect 20440 21520 21060 21536
rect 20440 21456 20478 21520
rect 20542 21456 20558 21520
rect 20622 21456 20638 21520
rect 20702 21456 20718 21520
rect 20782 21456 20798 21520
rect 20862 21456 20878 21520
rect 20942 21456 20958 21520
rect 21022 21456 21060 21520
rect 20440 21440 21060 21456
rect 8000 20976 8620 20992
rect 8000 20912 8038 20976
rect 8102 20912 8118 20976
rect 8182 20912 8198 20976
rect 8262 20912 8278 20976
rect 8342 20912 8358 20976
rect 8422 20912 8438 20976
rect 8502 20912 8518 20976
rect 8582 20912 8620 20976
rect 8000 20896 8620 20912
rect 13600 20976 14220 20992
rect 13600 20912 13638 20976
rect 13702 20912 13718 20976
rect 13782 20912 13798 20976
rect 13862 20912 13878 20976
rect 13942 20912 13958 20976
rect 14022 20912 14038 20976
rect 14102 20912 14118 20976
rect 14182 20912 14220 20976
rect 13600 20896 14220 20912
rect 19200 20976 19820 20992
rect 19200 20912 19238 20976
rect 19302 20912 19318 20976
rect 19382 20912 19398 20976
rect 19462 20912 19478 20976
rect 19542 20912 19558 20976
rect 19622 20912 19638 20976
rect 19702 20912 19718 20976
rect 19782 20912 19820 20976
rect 19200 20896 19820 20912
rect 9240 20432 9860 20448
rect 9240 20368 9278 20432
rect 9342 20368 9358 20432
rect 9422 20368 9438 20432
rect 9502 20368 9518 20432
rect 9582 20368 9598 20432
rect 9662 20368 9678 20432
rect 9742 20368 9758 20432
rect 9822 20368 9860 20432
rect 9240 20352 9860 20368
rect 14840 20432 15460 20448
rect 14840 20368 14878 20432
rect 14942 20368 14958 20432
rect 15022 20368 15038 20432
rect 15102 20368 15118 20432
rect 15182 20368 15198 20432
rect 15262 20368 15278 20432
rect 15342 20368 15358 20432
rect 15422 20368 15460 20432
rect 14840 20352 15460 20368
rect 20440 20432 21060 20448
rect 20440 20368 20478 20432
rect 20542 20368 20558 20432
rect 20622 20368 20638 20432
rect 20702 20368 20718 20432
rect 20782 20368 20798 20432
rect 20862 20368 20878 20432
rect 20942 20368 20958 20432
rect 21022 20368 21060 20432
rect 20440 20352 21060 20368
rect 23016 20234 28796 20294
rect 15929 20172 15995 20175
rect 19149 20172 19215 20175
rect 20069 20172 20135 20175
rect 22737 20172 22803 20175
rect 15929 20170 22803 20172
rect 15929 20114 15934 20170
rect 15990 20114 19154 20170
rect 19210 20114 20074 20170
rect 20130 20114 22742 20170
rect 22798 20114 22803 20170
rect 15929 20112 22803 20114
rect 15929 20109 15995 20112
rect 19149 20109 19215 20112
rect 20069 20109 20135 20112
rect 22737 20109 22803 20112
rect 8000 19888 8620 19904
rect 8000 19824 8038 19888
rect 8102 19824 8118 19888
rect 8182 19824 8198 19888
rect 8262 19824 8278 19888
rect 8342 19824 8358 19888
rect 8422 19824 8438 19888
rect 8502 19824 8518 19888
rect 8582 19824 8620 19888
rect 8000 19808 8620 19824
rect 13600 19888 14220 19904
rect 13600 19824 13638 19888
rect 13702 19824 13718 19888
rect 13782 19824 13798 19888
rect 13862 19824 13878 19888
rect 13942 19824 13958 19888
rect 14022 19824 14038 19888
rect 14102 19824 14118 19888
rect 14182 19824 14220 19888
rect 13600 19808 14220 19824
rect 19200 19888 19820 19904
rect 19200 19824 19238 19888
rect 19302 19824 19318 19888
rect 19382 19824 19398 19888
rect 19462 19824 19478 19888
rect 19542 19824 19558 19888
rect 19622 19824 19638 19888
rect 19702 19824 19718 19888
rect 19782 19824 19820 19888
rect 19200 19808 19820 19824
rect 19057 19684 19123 19687
rect 23016 19684 23076 20234
rect 19057 19682 23076 19684
rect 19057 19626 19062 19682
rect 19118 19626 23076 19682
rect 19057 19624 23076 19626
rect 19057 19621 19123 19624
rect 9240 19344 9860 19360
rect 9240 19280 9278 19344
rect 9342 19280 9358 19344
rect 9422 19280 9438 19344
rect 9502 19280 9518 19344
rect 9582 19280 9598 19344
rect 9662 19280 9678 19344
rect 9742 19280 9758 19344
rect 9822 19280 9860 19344
rect 9240 19264 9860 19280
rect 14840 19344 15460 19360
rect 14840 19280 14878 19344
rect 14942 19280 14958 19344
rect 15022 19280 15038 19344
rect 15102 19280 15118 19344
rect 15182 19280 15198 19344
rect 15262 19280 15278 19344
rect 15342 19280 15358 19344
rect 15422 19280 15460 19344
rect 14840 19264 15460 19280
rect 20440 19344 21060 19360
rect 20440 19280 20478 19344
rect 20542 19280 20558 19344
rect 20622 19280 20638 19344
rect 20702 19280 20718 19344
rect 20782 19280 20798 19344
rect 20862 19280 20878 19344
rect 20942 19280 20958 19344
rect 21022 19280 21060 19344
rect 20440 19264 21060 19280
rect 16849 19196 16915 19199
rect 22093 19196 22159 19199
rect 16849 19194 22159 19196
rect 16849 19138 16854 19194
rect 16910 19138 22098 19194
rect 22154 19138 22159 19194
rect 16849 19136 22159 19138
rect 16849 19133 16915 19136
rect 22093 19133 22159 19136
rect 8000 18800 8620 18816
rect 8000 18736 8038 18800
rect 8102 18736 8118 18800
rect 8182 18736 8198 18800
rect 8262 18736 8278 18800
rect 8342 18736 8358 18800
rect 8422 18736 8438 18800
rect 8502 18736 8518 18800
rect 8582 18736 8620 18800
rect 8000 18720 8620 18736
rect 13600 18800 14220 18816
rect 13600 18736 13638 18800
rect 13702 18736 13718 18800
rect 13782 18736 13798 18800
rect 13862 18736 13878 18800
rect 13942 18736 13958 18800
rect 14022 18736 14038 18800
rect 14102 18736 14118 18800
rect 14182 18736 14220 18800
rect 13600 18720 14220 18736
rect 19200 18800 19820 18816
rect 19200 18736 19238 18800
rect 19302 18736 19318 18800
rect 19382 18736 19398 18800
rect 19462 18736 19478 18800
rect 19542 18736 19558 18800
rect 19622 18736 19638 18800
rect 19702 18736 19718 18800
rect 19782 18736 19820 18800
rect 19200 18720 19820 18736
rect 9240 18256 9860 18272
rect 9240 18192 9278 18256
rect 9342 18192 9358 18256
rect 9422 18192 9438 18256
rect 9502 18192 9518 18256
rect 9582 18192 9598 18256
rect 9662 18192 9678 18256
rect 9742 18192 9758 18256
rect 9822 18192 9860 18256
rect 9240 18176 9860 18192
rect 14840 18256 15460 18272
rect 14840 18192 14878 18256
rect 14942 18192 14958 18256
rect 15022 18192 15038 18256
rect 15102 18192 15118 18256
rect 15182 18192 15198 18256
rect 15262 18192 15278 18256
rect 15342 18192 15358 18256
rect 15422 18192 15460 18256
rect 14840 18176 15460 18192
rect 20440 18256 21060 18272
rect 20440 18192 20478 18256
rect 20542 18192 20558 18256
rect 20622 18192 20638 18256
rect 20702 18192 20718 18256
rect 20782 18192 20798 18256
rect 20862 18192 20878 18256
rect 20942 18192 20958 18256
rect 21022 18192 21060 18256
rect 20440 18176 21060 18192
rect 17677 17854 17743 17857
rect 19793 17854 19859 17857
rect 17677 17852 19859 17854
rect 17677 17796 17682 17852
rect 17738 17796 19798 17852
rect 19854 17796 19859 17852
rect 17677 17794 19859 17796
rect 17677 17791 17743 17794
rect 19793 17791 19859 17794
rect 21633 17732 21699 17735
rect 21633 17730 28796 17732
rect 8000 17712 8620 17728
rect 8000 17648 8038 17712
rect 8102 17648 8118 17712
rect 8182 17648 8198 17712
rect 8262 17648 8278 17712
rect 8342 17648 8358 17712
rect 8422 17648 8438 17712
rect 8502 17648 8518 17712
rect 8582 17648 8620 17712
rect 8000 17632 8620 17648
rect 13600 17712 14220 17728
rect 13600 17648 13638 17712
rect 13702 17648 13718 17712
rect 13782 17648 13798 17712
rect 13862 17648 13878 17712
rect 13942 17648 13958 17712
rect 14022 17648 14038 17712
rect 14102 17648 14118 17712
rect 14182 17648 14220 17712
rect 13600 17632 14220 17648
rect 19200 17712 19820 17728
rect 19200 17648 19238 17712
rect 19302 17648 19318 17712
rect 19382 17648 19398 17712
rect 19462 17648 19478 17712
rect 19542 17648 19558 17712
rect 19622 17648 19638 17712
rect 19702 17648 19718 17712
rect 19782 17648 19820 17712
rect 21633 17674 21638 17730
rect 21694 17674 28796 17730
rect 21633 17672 28796 17674
rect 21633 17669 21699 17672
rect 19200 17632 19820 17648
rect 14273 17488 14339 17491
rect 14825 17488 14891 17491
rect 14273 17486 14891 17488
rect 14273 17430 14278 17486
rect 14334 17430 14830 17486
rect 14886 17430 14891 17486
rect 14273 17428 14891 17430
rect 14273 17425 14339 17428
rect 14825 17425 14891 17428
rect 17861 17488 17927 17491
rect 19517 17488 19583 17491
rect 17861 17486 19583 17488
rect 17861 17430 17866 17486
rect 17922 17430 19522 17486
rect 19578 17430 19583 17486
rect 17861 17428 19583 17430
rect 17861 17425 17927 17428
rect 19517 17425 19583 17428
rect 9240 17168 9860 17184
rect 9240 17104 9278 17168
rect 9342 17104 9358 17168
rect 9422 17104 9438 17168
rect 9502 17104 9518 17168
rect 9582 17104 9598 17168
rect 9662 17104 9678 17168
rect 9742 17104 9758 17168
rect 9822 17104 9860 17168
rect 9240 17088 9860 17104
rect 14840 17168 15460 17184
rect 14840 17104 14878 17168
rect 14942 17104 14958 17168
rect 15022 17104 15038 17168
rect 15102 17104 15118 17168
rect 15182 17104 15198 17168
rect 15262 17104 15278 17168
rect 15342 17104 15358 17168
rect 15422 17104 15460 17168
rect 14840 17088 15460 17104
rect 20440 17168 21060 17184
rect 20440 17104 20478 17168
rect 20542 17104 20558 17168
rect 20622 17104 20638 17168
rect 20702 17104 20718 17168
rect 20782 17104 20798 17168
rect 20862 17104 20878 17168
rect 20942 17104 20958 17168
rect 21022 17104 21060 17168
rect 20440 17088 21060 17104
rect 19517 16878 19583 16881
rect 20897 16878 20963 16881
rect 19517 16876 20963 16878
rect 19517 16820 19522 16876
rect 19578 16820 20902 16876
rect 20958 16820 20963 16876
rect 19517 16818 20963 16820
rect 19517 16815 19583 16818
rect 20897 16815 20963 16818
rect 8000 16624 8620 16640
rect 8000 16560 8038 16624
rect 8102 16560 8118 16624
rect 8182 16560 8198 16624
rect 8262 16560 8278 16624
rect 8342 16560 8358 16624
rect 8422 16560 8438 16624
rect 8502 16560 8518 16624
rect 8582 16560 8620 16624
rect 8000 16544 8620 16560
rect 13600 16624 14220 16640
rect 13600 16560 13638 16624
rect 13702 16560 13718 16624
rect 13782 16560 13798 16624
rect 13862 16560 13878 16624
rect 13942 16560 13958 16624
rect 14022 16560 14038 16624
rect 14102 16560 14118 16624
rect 14182 16560 14220 16624
rect 13600 16544 14220 16560
rect 19200 16624 19820 16640
rect 19200 16560 19238 16624
rect 19302 16560 19318 16624
rect 19382 16560 19398 16624
rect 19462 16560 19478 16624
rect 19542 16560 19558 16624
rect 19622 16560 19638 16624
rect 19702 16560 19718 16624
rect 19782 16560 19820 16624
rect 19200 16544 19820 16560
rect 16665 16390 16731 16393
rect 20069 16390 20135 16393
rect 21265 16392 21331 16393
rect 21260 16390 21266 16392
rect 16665 16388 20135 16390
rect 16665 16332 16670 16388
rect 16726 16332 20074 16388
rect 20130 16332 20135 16388
rect 16665 16330 20135 16332
rect 21176 16330 21266 16390
rect 16665 16327 16731 16330
rect 20069 16327 20135 16330
rect 21260 16328 21266 16330
rect 21330 16328 21336 16392
rect 21265 16327 21331 16328
rect 9240 16080 9860 16096
rect 7097 16024 7163 16027
rect 7465 16024 7531 16027
rect 7097 16022 7531 16024
rect 7097 15966 7102 16022
rect 7158 15966 7470 16022
rect 7526 15966 7531 16022
rect 9240 16016 9278 16080
rect 9342 16016 9358 16080
rect 9422 16016 9438 16080
rect 9502 16016 9518 16080
rect 9582 16016 9598 16080
rect 9662 16016 9678 16080
rect 9742 16016 9758 16080
rect 9822 16016 9860 16080
rect 9240 16000 9860 16016
rect 14840 16080 15460 16096
rect 14840 16016 14878 16080
rect 14942 16016 14958 16080
rect 15022 16016 15038 16080
rect 15102 16016 15118 16080
rect 15182 16016 15198 16080
rect 15262 16016 15278 16080
rect 15342 16016 15358 16080
rect 15422 16016 15460 16080
rect 14840 16000 15460 16016
rect 20440 16080 21060 16096
rect 20440 16016 20478 16080
rect 20542 16016 20558 16080
rect 20622 16016 20638 16080
rect 20702 16016 20718 16080
rect 20782 16016 20798 16080
rect 20862 16016 20878 16080
rect 20942 16016 20958 16080
rect 21022 16016 21060 16080
rect 20440 16000 21060 16016
rect 7097 15964 7531 15966
rect 7097 15961 7163 15964
rect 7465 15961 7531 15964
rect 15745 15902 15811 15905
rect 17309 15902 17375 15905
rect 15745 15900 17375 15902
rect 15745 15844 15750 15900
rect 15806 15844 17314 15900
rect 17370 15844 17375 15900
rect 15745 15842 17375 15844
rect 15745 15839 15811 15842
rect 17309 15839 17375 15842
rect 7281 15780 7347 15783
rect 8661 15780 8727 15783
rect 9489 15780 9555 15783
rect 10685 15780 10751 15783
rect 7281 15778 10751 15780
rect 7281 15722 7286 15778
rect 7342 15722 8666 15778
rect 8722 15722 9494 15778
rect 9550 15722 10690 15778
rect 10746 15722 10751 15778
rect 7281 15720 10751 15722
rect 7281 15717 7347 15720
rect 8661 15717 8727 15720
rect 9489 15717 9555 15720
rect 10685 15717 10751 15720
rect 8000 15536 8620 15552
rect 8000 15472 8038 15536
rect 8102 15472 8118 15536
rect 8182 15472 8198 15536
rect 8262 15472 8278 15536
rect 8342 15472 8358 15536
rect 8422 15472 8438 15536
rect 8502 15472 8518 15536
rect 8582 15472 8620 15536
rect 8000 15456 8620 15472
rect 13600 15536 14220 15552
rect 13600 15472 13638 15536
rect 13702 15472 13718 15536
rect 13782 15472 13798 15536
rect 13862 15472 13878 15536
rect 13942 15472 13958 15536
rect 14022 15472 14038 15536
rect 14102 15472 14118 15536
rect 14182 15472 14220 15536
rect 13600 15456 14220 15472
rect 19200 15536 19820 15552
rect 19200 15472 19238 15536
rect 19302 15472 19318 15536
rect 19382 15472 19398 15536
rect 19462 15472 19478 15536
rect 19542 15472 19558 15536
rect 19622 15472 19638 15536
rect 19702 15472 19718 15536
rect 19782 15472 19820 15536
rect 19200 15456 19820 15472
rect 22921 15292 22987 15295
rect 22921 15290 28796 15292
rect 22921 15234 22926 15290
rect 22982 15234 28796 15290
rect 22921 15232 28796 15234
rect 22921 15229 22987 15232
rect 18505 15170 18571 15173
rect 21449 15170 21515 15173
rect 18505 15168 21515 15170
rect 18505 15112 18510 15168
rect 18566 15112 21454 15168
rect 21510 15112 21515 15168
rect 18505 15110 21515 15112
rect 18505 15107 18571 15110
rect 21449 15107 21515 15110
rect 9240 14992 9860 15008
rect 9240 14928 9278 14992
rect 9342 14928 9358 14992
rect 9422 14928 9438 14992
rect 9502 14928 9518 14992
rect 9582 14928 9598 14992
rect 9662 14928 9678 14992
rect 9742 14928 9758 14992
rect 9822 14928 9860 14992
rect 9240 14912 9860 14928
rect 14840 14992 15460 15008
rect 14840 14928 14878 14992
rect 14942 14928 14958 14992
rect 15022 14928 15038 14992
rect 15102 14928 15118 14992
rect 15182 14928 15198 14992
rect 15262 14928 15278 14992
rect 15342 14928 15358 14992
rect 15422 14928 15460 14992
rect 14840 14912 15460 14928
rect 20440 14992 21060 15008
rect 20440 14928 20478 14992
rect 20542 14928 20558 14992
rect 20622 14928 20638 14992
rect 20702 14928 20718 14992
rect 20782 14928 20798 14992
rect 20862 14928 20878 14992
rect 20942 14928 20958 14992
rect 21022 14928 21060 14992
rect 20440 14912 21060 14928
rect 13 14804 79 14807
rect 10593 14804 10659 14807
rect 13 14802 10659 14804
rect 13 14746 18 14802
rect 74 14746 10598 14802
rect 10654 14746 10659 14802
rect 13 14744 10659 14746
rect 13 14741 79 14744
rect 10593 14741 10659 14744
rect 19057 14804 19123 14807
rect 20621 14804 20687 14807
rect 19057 14802 20687 14804
rect 19057 14746 19062 14802
rect 19118 14746 20626 14802
rect 20682 14746 20687 14802
rect 19057 14744 20687 14746
rect 19057 14741 19123 14744
rect 20621 14741 20687 14744
rect 16205 14682 16271 14685
rect 17953 14682 18019 14685
rect 16205 14680 18019 14682
rect 16205 14624 16210 14680
rect 16266 14624 17958 14680
rect 18014 14624 18019 14680
rect 16205 14622 18019 14624
rect 16205 14619 16271 14622
rect 17953 14619 18019 14622
rect 20437 14560 20503 14563
rect 21265 14560 21331 14563
rect 20437 14558 21331 14560
rect 20437 14502 20442 14558
rect 20498 14502 21270 14558
rect 21326 14502 21331 14558
rect 20437 14500 21331 14502
rect 20437 14497 20503 14500
rect 21265 14497 21331 14500
rect 8000 14448 8620 14464
rect 8000 14384 8038 14448
rect 8102 14384 8118 14448
rect 8182 14384 8198 14448
rect 8262 14384 8278 14448
rect 8342 14384 8358 14448
rect 8422 14384 8438 14448
rect 8502 14384 8518 14448
rect 8582 14384 8620 14448
rect 8000 14368 8620 14384
rect 13600 14448 14220 14464
rect 13600 14384 13638 14448
rect 13702 14384 13718 14448
rect 13782 14384 13798 14448
rect 13862 14384 13878 14448
rect 13942 14384 13958 14448
rect 14022 14384 14038 14448
rect 14102 14384 14118 14448
rect 14182 14384 14220 14448
rect 13600 14368 14220 14384
rect 19200 14448 19820 14464
rect 19200 14384 19238 14448
rect 19302 14384 19318 14448
rect 19382 14384 19398 14448
rect 19462 14384 19478 14448
rect 19542 14384 19558 14448
rect 19622 14384 19638 14448
rect 19702 14384 19718 14448
rect 19782 14384 19820 14448
rect 19200 14368 19820 14384
rect 21265 14316 21331 14319
rect 22093 14316 22159 14319
rect 21265 14314 22159 14316
rect 21265 14258 21270 14314
rect 21326 14258 22098 14314
rect 22154 14258 22159 14314
rect 21265 14256 22159 14258
rect 21265 14253 21331 14256
rect 22093 14253 22159 14256
rect 14733 14194 14799 14197
rect 15745 14194 15811 14197
rect 14733 14192 15811 14194
rect 14733 14136 14738 14192
rect 14794 14136 15750 14192
rect 15806 14136 15811 14192
rect 14733 14134 15811 14136
rect 14733 14131 14799 14134
rect 15745 14131 15811 14134
rect 9240 13904 9860 13920
rect 9240 13840 9278 13904
rect 9342 13840 9358 13904
rect 9422 13840 9438 13904
rect 9502 13840 9518 13904
rect 9582 13840 9598 13904
rect 9662 13840 9678 13904
rect 9742 13840 9758 13904
rect 9822 13840 9860 13904
rect 5809 13828 5875 13831
rect 0 13826 5875 13828
rect 0 13770 5814 13826
rect 5870 13770 5875 13826
rect 9240 13824 9860 13840
rect 14840 13904 15460 13920
rect 14840 13840 14878 13904
rect 14942 13840 14958 13904
rect 15022 13840 15038 13904
rect 15102 13840 15118 13904
rect 15182 13840 15198 13904
rect 15262 13840 15278 13904
rect 15342 13840 15358 13904
rect 15422 13840 15460 13904
rect 14840 13824 15460 13840
rect 20440 13904 21060 13920
rect 20440 13840 20478 13904
rect 20542 13840 20558 13904
rect 20622 13840 20638 13904
rect 20702 13840 20718 13904
rect 20782 13840 20798 13904
rect 20862 13840 20878 13904
rect 20942 13840 20958 13904
rect 21022 13840 21060 13904
rect 20440 13824 21060 13840
rect 0 13768 5875 13770
rect 5809 13765 5875 13768
rect 14549 13706 14615 13709
rect 15285 13706 15351 13709
rect 14549 13704 15351 13706
rect 14549 13648 14554 13704
rect 14610 13648 15290 13704
rect 15346 13648 15351 13704
rect 14549 13646 15351 13648
rect 14549 13643 14615 13646
rect 15285 13643 15351 13646
rect 19057 13706 19123 13709
rect 20437 13706 20503 13709
rect 19057 13704 20503 13706
rect 19057 13648 19062 13704
rect 19118 13648 20442 13704
rect 20498 13648 20503 13704
rect 19057 13646 20503 13648
rect 19057 13643 19123 13646
rect 20437 13643 20503 13646
rect 8000 13360 8620 13376
rect 8000 13296 8038 13360
rect 8102 13296 8118 13360
rect 8182 13296 8198 13360
rect 8262 13296 8278 13360
rect 8342 13296 8358 13360
rect 8422 13296 8438 13360
rect 8502 13296 8518 13360
rect 8582 13296 8620 13360
rect 8000 13280 8620 13296
rect 13600 13360 14220 13376
rect 13600 13296 13638 13360
rect 13702 13296 13718 13360
rect 13782 13296 13798 13360
rect 13862 13296 13878 13360
rect 13942 13296 13958 13360
rect 14022 13296 14038 13360
rect 14102 13296 14118 13360
rect 14182 13296 14220 13360
rect 13600 13280 14220 13296
rect 19200 13360 19820 13376
rect 19200 13296 19238 13360
rect 19302 13296 19318 13360
rect 19382 13296 19398 13360
rect 19462 13296 19478 13360
rect 19542 13296 19558 13360
rect 19622 13296 19638 13360
rect 19702 13296 19718 13360
rect 19782 13296 19820 13360
rect 19200 13280 19820 13296
rect 15469 13218 15535 13221
rect 17493 13218 17559 13221
rect 18781 13218 18847 13221
rect 15469 13216 18847 13218
rect 15469 13160 15474 13216
rect 15530 13160 17498 13216
rect 17554 13160 18786 13216
rect 18842 13160 18847 13216
rect 15469 13158 18847 13160
rect 15469 13155 15535 13158
rect 17493 13155 17559 13158
rect 18781 13155 18847 13158
rect 20805 13218 20871 13221
rect 21265 13218 21331 13221
rect 22001 13218 22067 13221
rect 20805 13216 22067 13218
rect 20805 13160 20810 13216
rect 20866 13160 21270 13216
rect 21326 13160 22006 13216
rect 22062 13160 22067 13216
rect 20805 13158 22067 13160
rect 20805 13155 20871 13158
rect 21265 13155 21331 13158
rect 22001 13155 22067 13158
rect 15285 12974 15351 12977
rect 16757 12974 16823 12977
rect 15285 12972 16823 12974
rect 15285 12916 15290 12972
rect 15346 12916 16762 12972
rect 16818 12916 16823 12972
rect 15285 12914 16823 12916
rect 15285 12911 15351 12914
rect 9240 12816 9860 12832
rect 9240 12752 9278 12816
rect 9342 12752 9358 12816
rect 9422 12752 9438 12816
rect 9502 12752 9518 12816
rect 9582 12752 9598 12816
rect 9662 12752 9678 12816
rect 9742 12752 9758 12816
rect 9822 12752 9860 12816
rect 9240 12736 9860 12752
rect 14840 12816 15460 12832
rect 14840 12752 14878 12816
rect 14942 12752 14958 12816
rect 15022 12752 15038 12816
rect 15102 12752 15118 12816
rect 15182 12752 15198 12816
rect 15262 12752 15278 12816
rect 15342 12752 15358 12816
rect 15422 12752 15460 12816
rect 14840 12736 15460 12752
rect 12341 12608 12407 12611
rect 13261 12608 13327 12611
rect 12341 12606 13327 12608
rect 12341 12550 12346 12606
rect 12402 12550 13266 12606
rect 13322 12550 13327 12606
rect 12341 12548 13327 12550
rect 12341 12545 12407 12548
rect 13261 12545 13327 12548
rect 15840 12367 15900 12914
rect 16757 12911 16823 12914
rect 20529 12974 20595 12977
rect 20529 12972 22524 12974
rect 20529 12916 20534 12972
rect 20590 12916 22524 12972
rect 20529 12914 22524 12916
rect 20529 12911 20595 12914
rect 20440 12816 21060 12832
rect 20440 12752 20478 12816
rect 20542 12752 20558 12816
rect 20622 12752 20638 12816
rect 20702 12752 20718 12816
rect 20782 12752 20798 12816
rect 20862 12752 20878 12816
rect 20942 12752 20958 12816
rect 21022 12752 21060 12816
rect 20440 12736 21060 12752
rect 22464 12730 22524 12914
rect 22464 12670 28796 12730
rect 16757 12608 16823 12611
rect 17493 12608 17559 12611
rect 16757 12606 17559 12608
rect 16757 12550 16762 12606
rect 16818 12550 17498 12606
rect 17554 12550 17559 12606
rect 16757 12548 17559 12550
rect 16757 12545 16823 12548
rect 17493 12545 17559 12548
rect 18597 12608 18663 12611
rect 20161 12608 20227 12611
rect 18597 12606 20227 12608
rect 18597 12550 18602 12606
rect 18658 12550 20166 12606
rect 20222 12550 20227 12606
rect 18597 12548 20227 12550
rect 18597 12545 18663 12548
rect 20161 12545 20227 12548
rect 21081 12486 21147 12489
rect 22737 12486 22803 12489
rect 21081 12484 22803 12486
rect 21081 12428 21086 12484
rect 21142 12428 22742 12484
rect 22798 12428 22803 12484
rect 21081 12426 22803 12428
rect 21081 12423 21147 12426
rect 22737 12423 22803 12426
rect 15837 12362 15903 12367
rect 15837 12306 15842 12362
rect 15898 12306 15903 12362
rect 15837 12301 15903 12306
rect 8000 12272 8620 12288
rect 8000 12208 8038 12272
rect 8102 12208 8118 12272
rect 8182 12208 8198 12272
rect 8262 12208 8278 12272
rect 8342 12208 8358 12272
rect 8422 12208 8438 12272
rect 8502 12208 8518 12272
rect 8582 12208 8620 12272
rect 8000 12192 8620 12208
rect 13600 12272 14220 12288
rect 13600 12208 13638 12272
rect 13702 12208 13718 12272
rect 13782 12208 13798 12272
rect 13862 12208 13878 12272
rect 13942 12208 13958 12272
rect 14022 12208 14038 12272
rect 14102 12208 14118 12272
rect 14182 12208 14220 12272
rect 13600 12192 14220 12208
rect 19200 12272 19820 12288
rect 19200 12208 19238 12272
rect 19302 12208 19318 12272
rect 19382 12208 19398 12272
rect 19462 12208 19478 12272
rect 19542 12208 19558 12272
rect 19622 12208 19638 12272
rect 19702 12208 19718 12272
rect 19782 12208 19820 12272
rect 19200 12192 19820 12208
rect 13997 11998 14063 12001
rect 15469 11998 15535 12001
rect 13997 11996 15535 11998
rect 13997 11940 14002 11996
rect 14058 11940 15474 11996
rect 15530 11940 15535 11996
rect 13997 11938 15535 11940
rect 13997 11935 14063 11938
rect 15469 11935 15535 11938
rect 21173 12000 21336 12001
rect 21173 11996 21266 12000
rect 21173 11940 21178 11996
rect 21234 11940 21266 11996
rect 21173 11936 21266 11940
rect 21330 11936 21336 12000
rect 21173 11935 21336 11936
rect 9240 11728 9860 11744
rect 9240 11664 9278 11728
rect 9342 11664 9358 11728
rect 9422 11664 9438 11728
rect 9502 11664 9518 11728
rect 9582 11664 9598 11728
rect 9662 11664 9678 11728
rect 9742 11664 9758 11728
rect 9822 11664 9860 11728
rect 9240 11648 9860 11664
rect 14840 11728 15460 11744
rect 14840 11664 14878 11728
rect 14942 11664 14958 11728
rect 15022 11664 15038 11728
rect 15102 11664 15118 11728
rect 15182 11664 15198 11728
rect 15262 11664 15278 11728
rect 15342 11664 15358 11728
rect 15422 11664 15460 11728
rect 14840 11648 15460 11664
rect 20440 11728 21060 11744
rect 20440 11664 20478 11728
rect 20542 11664 20558 11728
rect 20622 11664 20638 11728
rect 20702 11664 20718 11728
rect 20782 11664 20798 11728
rect 20862 11664 20878 11728
rect 20942 11664 20958 11728
rect 21022 11664 21060 11728
rect 20440 11648 21060 11664
rect 8000 11184 8620 11200
rect 8000 11120 8038 11184
rect 8102 11120 8118 11184
rect 8182 11120 8198 11184
rect 8262 11120 8278 11184
rect 8342 11120 8358 11184
rect 8422 11120 8438 11184
rect 8502 11120 8518 11184
rect 8582 11120 8620 11184
rect 8000 11104 8620 11120
rect 13600 11184 14220 11200
rect 13600 11120 13638 11184
rect 13702 11120 13718 11184
rect 13782 11120 13798 11184
rect 13862 11120 13878 11184
rect 13942 11120 13958 11184
rect 14022 11120 14038 11184
rect 14102 11120 14118 11184
rect 14182 11120 14220 11184
rect 13600 11104 14220 11120
rect 19200 11184 19820 11200
rect 19200 11120 19238 11184
rect 19302 11120 19318 11184
rect 19382 11120 19398 11184
rect 19462 11120 19478 11184
rect 19542 11120 19558 11184
rect 19622 11120 19638 11184
rect 19702 11120 19718 11184
rect 19782 11120 19820 11184
rect 19200 11104 19820 11120
rect 16849 10656 16915 10659
rect 18505 10656 18571 10659
rect 9240 10640 9860 10656
rect 9240 10576 9278 10640
rect 9342 10576 9358 10640
rect 9422 10576 9438 10640
rect 9502 10576 9518 10640
rect 9582 10576 9598 10640
rect 9662 10576 9678 10640
rect 9742 10576 9758 10640
rect 9822 10576 9860 10640
rect 9240 10560 9860 10576
rect 14840 10640 15460 10656
rect 14840 10576 14878 10640
rect 14942 10576 14958 10640
rect 15022 10576 15038 10640
rect 15102 10576 15118 10640
rect 15182 10576 15198 10640
rect 15262 10576 15278 10640
rect 15342 10576 15358 10640
rect 15422 10576 15460 10640
rect 16849 10654 18571 10656
rect 16849 10598 16854 10654
rect 16910 10598 18510 10654
rect 18566 10598 18571 10654
rect 16849 10596 18571 10598
rect 16849 10593 16915 10596
rect 18505 10593 18571 10596
rect 20440 10640 21060 10656
rect 14840 10560 15460 10576
rect 20440 10576 20478 10640
rect 20542 10576 20558 10640
rect 20622 10576 20638 10640
rect 20702 10576 20718 10640
rect 20782 10576 20798 10640
rect 20862 10576 20878 10640
rect 20942 10576 20958 10640
rect 21022 10576 21060 10640
rect 20440 10560 21060 10576
rect 15745 10412 15811 10415
rect 17953 10412 18019 10415
rect 15745 10410 18292 10412
rect 15745 10354 15750 10410
rect 15806 10354 17958 10410
rect 18014 10354 18292 10410
rect 15745 10352 18292 10354
rect 15745 10349 15811 10352
rect 17953 10349 18019 10352
rect 10041 10290 10107 10293
rect 18232 10290 18292 10352
rect 20345 10290 20411 10293
rect 10041 10288 14428 10290
rect 10041 10232 10046 10288
rect 10102 10232 14428 10288
rect 10041 10230 14428 10232
rect 18232 10288 20411 10290
rect 18232 10232 20350 10288
rect 20406 10232 20411 10288
rect 18232 10230 20411 10232
rect 10041 10227 10107 10230
rect 14368 10168 14428 10230
rect 20345 10227 20411 10230
rect 21817 10290 21883 10293
rect 21817 10288 28796 10290
rect 21817 10232 21822 10288
rect 21878 10232 28796 10288
rect 21817 10230 28796 10232
rect 21817 10227 21883 10230
rect 18137 10168 18203 10171
rect 14368 10166 18203 10168
rect 8000 10096 8620 10112
rect 8000 10032 8038 10096
rect 8102 10032 8118 10096
rect 8182 10032 8198 10096
rect 8262 10032 8278 10096
rect 8342 10032 8358 10096
rect 8422 10032 8438 10096
rect 8502 10032 8518 10096
rect 8582 10032 8620 10096
rect 8000 10016 8620 10032
rect 13600 10096 14220 10112
rect 14368 10110 18142 10166
rect 18198 10110 18203 10166
rect 14368 10108 18203 10110
rect 18137 10105 18203 10108
rect 13600 10032 13638 10096
rect 13702 10032 13718 10096
rect 13782 10032 13798 10096
rect 13862 10032 13878 10096
rect 13942 10032 13958 10096
rect 14022 10032 14038 10096
rect 14102 10032 14118 10096
rect 14182 10032 14220 10096
rect 13600 10016 14220 10032
rect 19200 10096 19820 10112
rect 19200 10032 19238 10096
rect 19302 10032 19318 10096
rect 19382 10032 19398 10096
rect 19462 10032 19478 10096
rect 19542 10032 19558 10096
rect 19622 10032 19638 10096
rect 19702 10032 19718 10096
rect 19782 10032 19820 10096
rect 19200 10016 19820 10032
rect 18045 9924 18111 9927
rect 21449 9924 21515 9927
rect 18045 9922 21515 9924
rect 18045 9866 18050 9922
rect 18106 9866 21454 9922
rect 21510 9866 21515 9922
rect 18045 9864 21515 9866
rect 18045 9861 18111 9864
rect 21449 9861 21515 9864
rect 16297 9680 16363 9683
rect 19149 9680 19215 9683
rect 16297 9678 19215 9680
rect 16297 9622 16302 9678
rect 16358 9622 19154 9678
rect 19210 9622 19215 9678
rect 16297 9620 19215 9622
rect 16297 9617 16363 9620
rect 9240 9552 9860 9568
rect 9240 9488 9278 9552
rect 9342 9488 9358 9552
rect 9422 9488 9438 9552
rect 9502 9488 9518 9552
rect 9582 9488 9598 9552
rect 9662 9488 9678 9552
rect 9742 9488 9758 9552
rect 9822 9488 9860 9552
rect 9240 9472 9860 9488
rect 14840 9552 15460 9568
rect 17128 9560 17188 9620
rect 19149 9617 19215 9620
rect 14840 9488 14878 9552
rect 14942 9488 14958 9552
rect 15022 9488 15038 9552
rect 15102 9488 15118 9552
rect 15182 9488 15198 9552
rect 15262 9488 15278 9552
rect 15342 9488 15358 9552
rect 15422 9488 15460 9552
rect 17120 9496 17126 9560
rect 17190 9496 17196 9560
rect 20440 9552 21060 9568
rect 14840 9472 15460 9488
rect 20440 9488 20478 9552
rect 20542 9488 20558 9552
rect 20622 9488 20638 9552
rect 20702 9488 20718 9552
rect 20782 9488 20798 9552
rect 20862 9488 20878 9552
rect 20942 9488 20958 9552
rect 21022 9488 21060 9552
rect 20440 9472 21060 9488
rect 15653 9436 15719 9439
rect 15653 9434 16636 9436
rect 15653 9378 15658 9434
rect 15714 9378 16636 9434
rect 15653 9376 16636 9378
rect 15653 9373 15719 9376
rect 16576 9314 16636 9376
rect 20161 9314 20227 9317
rect 16576 9312 20227 9314
rect 16576 9256 20166 9312
rect 20222 9256 20227 9312
rect 16576 9254 20227 9256
rect 20161 9251 20227 9254
rect 8000 9008 8620 9024
rect 8000 8944 8038 9008
rect 8102 8944 8118 9008
rect 8182 8944 8198 9008
rect 8262 8944 8278 9008
rect 8342 8944 8358 9008
rect 8422 8944 8438 9008
rect 8502 8944 8518 9008
rect 8582 8944 8620 9008
rect 8000 8928 8620 8944
rect 13600 9008 14220 9024
rect 13600 8944 13638 9008
rect 13702 8944 13718 9008
rect 13782 8944 13798 9008
rect 13862 8944 13878 9008
rect 13942 8944 13958 9008
rect 14022 8944 14038 9008
rect 14102 8944 14118 9008
rect 14182 8944 14220 9008
rect 13600 8928 14220 8944
rect 19200 9008 19820 9024
rect 19200 8944 19238 9008
rect 19302 8944 19318 9008
rect 19382 8944 19398 9008
rect 19462 8944 19478 9008
rect 19542 8944 19558 9008
rect 19622 8944 19638 9008
rect 19702 8944 19718 9008
rect 19782 8944 19820 9008
rect 19200 8928 19820 8944
rect 13445 8826 13511 8829
rect 15469 8826 15535 8829
rect 16021 8826 16087 8829
rect 18689 8826 18755 8829
rect 13445 8824 18755 8826
rect 13445 8768 13450 8824
rect 13506 8768 15474 8824
rect 15530 8768 16026 8824
rect 16082 8768 18694 8824
rect 18750 8768 18755 8824
rect 13445 8766 18755 8768
rect 13445 8763 13511 8766
rect 15469 8763 15535 8766
rect 16021 8763 16087 8766
rect 18689 8763 18755 8766
rect 16205 8582 16271 8585
rect 17033 8582 17099 8585
rect 20253 8582 20319 8585
rect 16205 8580 17464 8582
rect 16205 8524 16210 8580
rect 16266 8524 17038 8580
rect 17094 8524 17464 8580
rect 16205 8522 17464 8524
rect 16205 8519 16271 8522
rect 17033 8519 17099 8522
rect 9240 8464 9860 8480
rect 9240 8400 9278 8464
rect 9342 8400 9358 8464
rect 9422 8400 9438 8464
rect 9502 8400 9518 8464
rect 9582 8400 9598 8464
rect 9662 8400 9678 8464
rect 9742 8400 9758 8464
rect 9822 8400 9860 8464
rect 9240 8384 9860 8400
rect 14840 8464 15460 8480
rect 14840 8400 14878 8464
rect 14942 8400 14958 8464
rect 15022 8400 15038 8464
rect 15102 8400 15118 8464
rect 15182 8400 15198 8464
rect 15262 8400 15278 8464
rect 15342 8400 15358 8464
rect 15422 8400 15460 8464
rect 14840 8384 15460 8400
rect 17404 8338 17464 8522
rect 19980 8580 20319 8582
rect 19980 8524 20258 8580
rect 20314 8524 20319 8580
rect 19980 8522 20319 8524
rect 19980 8338 20040 8522
rect 20253 8519 20319 8522
rect 20440 8464 21060 8480
rect 20440 8400 20478 8464
rect 20542 8400 20558 8464
rect 20622 8400 20638 8464
rect 20702 8400 20718 8464
rect 20782 8400 20798 8464
rect 20862 8400 20878 8464
rect 20942 8400 20958 8464
rect 21022 8400 21060 8464
rect 20440 8384 21060 8400
rect 21265 8340 21331 8341
rect 21260 8338 21266 8340
rect 17404 8278 20040 8338
rect 21176 8278 21266 8338
rect 21260 8276 21266 8278
rect 21330 8276 21336 8340
rect 21265 8275 21331 8276
rect 20529 8094 20595 8097
rect 22737 8094 22803 8097
rect 28533 8094 28599 8097
rect 20529 8092 28599 8094
rect 20529 8036 20534 8092
rect 20590 8036 22742 8092
rect 22798 8036 28538 8092
rect 28594 8036 28599 8092
rect 20529 8034 28599 8036
rect 20529 8031 20595 8034
rect 22737 8031 22803 8034
rect 28533 8031 28599 8034
rect 17125 7974 17191 7975
rect 17120 7972 17126 7974
rect 8000 7920 8620 7936
rect 8000 7856 8038 7920
rect 8102 7856 8118 7920
rect 8182 7856 8198 7920
rect 8262 7856 8278 7920
rect 8342 7856 8358 7920
rect 8422 7856 8438 7920
rect 8502 7856 8518 7920
rect 8582 7856 8620 7920
rect 8000 7840 8620 7856
rect 13600 7920 14220 7936
rect 13600 7856 13638 7920
rect 13702 7856 13718 7920
rect 13782 7856 13798 7920
rect 13862 7856 13878 7920
rect 13942 7856 13958 7920
rect 14022 7856 14038 7920
rect 14102 7856 14118 7920
rect 14182 7856 14220 7920
rect 17036 7912 17126 7972
rect 17120 7910 17126 7912
rect 17190 7910 17196 7974
rect 19200 7920 19820 7936
rect 17125 7909 17191 7910
rect 13600 7840 14220 7856
rect 19200 7856 19238 7920
rect 19302 7856 19318 7920
rect 19382 7856 19398 7920
rect 19462 7856 19478 7920
rect 19542 7856 19558 7920
rect 19622 7856 19638 7920
rect 19702 7856 19718 7920
rect 19782 7856 19820 7920
rect 19200 7840 19820 7856
rect 9121 7728 9187 7731
rect 10685 7728 10751 7731
rect 12341 7728 12407 7731
rect 13629 7728 13695 7731
rect 14641 7728 14707 7731
rect 16205 7728 16271 7731
rect 18781 7728 18847 7731
rect 19241 7728 19307 7731
rect 19793 7728 19859 7731
rect 21357 7728 21423 7731
rect 9121 7726 21423 7728
rect 9121 7670 9126 7726
rect 9182 7670 10690 7726
rect 10746 7670 12346 7726
rect 12402 7670 13634 7726
rect 13690 7670 14646 7726
rect 14702 7670 16210 7726
rect 16266 7670 18786 7726
rect 18842 7670 19246 7726
rect 19302 7670 19798 7726
rect 19854 7670 21362 7726
rect 21418 7670 21423 7726
rect 9121 7668 21423 7670
rect 9121 7665 9187 7668
rect 10685 7665 10751 7668
rect 12341 7665 12407 7668
rect 13629 7665 13695 7668
rect 14641 7665 14707 7668
rect 16205 7665 16271 7668
rect 18781 7665 18847 7668
rect 19241 7665 19307 7668
rect 19793 7665 19859 7668
rect 21357 7665 21423 7668
rect 22001 7728 22067 7731
rect 22001 7726 28796 7728
rect 22001 7670 22006 7726
rect 22062 7670 28796 7726
rect 22001 7668 28796 7670
rect 22001 7665 22067 7668
rect 9240 7376 9860 7392
rect 9240 7312 9278 7376
rect 9342 7312 9358 7376
rect 9422 7312 9438 7376
rect 9502 7312 9518 7376
rect 9582 7312 9598 7376
rect 9662 7312 9678 7376
rect 9742 7312 9758 7376
rect 9822 7312 9860 7376
rect 9240 7296 9860 7312
rect 14840 7376 15460 7392
rect 14840 7312 14878 7376
rect 14942 7312 14958 7376
rect 15022 7312 15038 7376
rect 15102 7312 15118 7376
rect 15182 7312 15198 7376
rect 15262 7312 15278 7376
rect 15342 7312 15358 7376
rect 15422 7312 15460 7376
rect 14840 7296 15460 7312
rect 20440 7376 21060 7392
rect 20440 7312 20478 7376
rect 20542 7312 20558 7376
rect 20622 7312 20638 7376
rect 20702 7312 20718 7376
rect 20782 7312 20798 7376
rect 20862 7312 20878 7376
rect 20942 7312 20958 7376
rect 21022 7312 21060 7376
rect 20440 7296 21060 7312
rect 9305 6996 9371 6999
rect 18597 6996 18663 6999
rect 9305 6994 18663 6996
rect 9305 6938 9310 6994
rect 9366 6938 18602 6994
rect 18658 6938 18663 6994
rect 9305 6936 18663 6938
rect 9305 6933 9371 6936
rect 18597 6933 18663 6936
rect 8000 6832 8620 6848
rect 8000 6768 8038 6832
rect 8102 6768 8118 6832
rect 8182 6768 8198 6832
rect 8262 6768 8278 6832
rect 8342 6768 8358 6832
rect 8422 6768 8438 6832
rect 8502 6768 8518 6832
rect 8582 6768 8620 6832
rect 8000 6752 8620 6768
rect 13600 6832 14220 6848
rect 13600 6768 13638 6832
rect 13702 6768 13718 6832
rect 13782 6768 13798 6832
rect 13862 6768 13878 6832
rect 13942 6768 13958 6832
rect 14022 6768 14038 6832
rect 14102 6768 14118 6832
rect 14182 6768 14220 6832
rect 13600 6752 14220 6768
rect 19200 6832 19820 6848
rect 19200 6768 19238 6832
rect 19302 6768 19318 6832
rect 19382 6768 19398 6832
rect 19462 6768 19478 6832
rect 19542 6768 19558 6832
rect 19622 6768 19638 6832
rect 19702 6768 19718 6832
rect 19782 6768 19820 6832
rect 19200 6752 19820 6768
rect 7281 6630 7347 6633
rect 10225 6630 10291 6633
rect 7281 6628 10291 6630
rect 7281 6572 7286 6628
rect 7342 6572 10230 6628
rect 10286 6572 10291 6628
rect 7281 6570 10291 6572
rect 7281 6567 7347 6570
rect 8201 6386 8267 6389
rect 8480 6386 8540 6570
rect 10225 6567 10291 6570
rect 18781 6508 18847 6511
rect 21633 6508 21699 6511
rect 18781 6506 21699 6508
rect 18781 6450 18786 6506
rect 18842 6450 21638 6506
rect 21694 6450 21699 6506
rect 18781 6448 21699 6450
rect 18781 6445 18847 6448
rect 21633 6445 21699 6448
rect 8201 6384 8540 6386
rect 8201 6328 8206 6384
rect 8262 6328 8540 6384
rect 8201 6326 8540 6328
rect 8201 6323 8267 6326
rect 9240 6288 9860 6304
rect 9240 6224 9278 6288
rect 9342 6224 9358 6288
rect 9422 6224 9438 6288
rect 9502 6224 9518 6288
rect 9582 6224 9598 6288
rect 9662 6224 9678 6288
rect 9742 6224 9758 6288
rect 9822 6224 9860 6288
rect 9240 6208 9860 6224
rect 14840 6288 15460 6304
rect 14840 6224 14878 6288
rect 14942 6224 14958 6288
rect 15022 6224 15038 6288
rect 15102 6224 15118 6288
rect 15182 6224 15198 6288
rect 15262 6224 15278 6288
rect 15342 6224 15358 6288
rect 15422 6224 15460 6288
rect 14840 6208 15460 6224
rect 20440 6288 21060 6304
rect 20440 6224 20478 6288
rect 20542 6224 20558 6288
rect 20622 6224 20638 6288
rect 20702 6224 20718 6288
rect 20782 6224 20798 6288
rect 20862 6224 20878 6288
rect 20942 6224 20958 6288
rect 21022 6224 21060 6288
rect 20440 6208 21060 6224
rect 22461 6262 22527 6267
rect 22461 6206 22466 6262
rect 22522 6206 22527 6262
rect 22461 6201 22527 6206
rect 12249 6020 12315 6023
rect 13261 6020 13327 6023
rect 12249 6018 13327 6020
rect 12249 5962 12254 6018
rect 12310 5962 13266 6018
rect 13322 5962 13327 6018
rect 12249 5960 13327 5962
rect 12249 5957 12315 5960
rect 13261 5957 13327 5960
rect 16849 6020 16915 6023
rect 22464 6020 22524 6201
rect 16849 6018 22524 6020
rect 16849 5962 16854 6018
rect 16910 5962 22524 6018
rect 16849 5960 22524 5962
rect 16849 5957 16915 5960
rect 8000 5744 8620 5760
rect 8000 5680 8038 5744
rect 8102 5680 8118 5744
rect 8182 5680 8198 5744
rect 8262 5680 8278 5744
rect 8342 5680 8358 5744
rect 8422 5680 8438 5744
rect 8502 5680 8518 5744
rect 8582 5680 8620 5744
rect 8000 5664 8620 5680
rect 13600 5744 14220 5760
rect 13600 5680 13638 5744
rect 13702 5680 13718 5744
rect 13782 5680 13798 5744
rect 13862 5680 13878 5744
rect 13942 5680 13958 5744
rect 14022 5680 14038 5744
rect 14102 5680 14118 5744
rect 14182 5680 14220 5744
rect 13600 5664 14220 5680
rect 19200 5744 19820 5760
rect 19200 5680 19238 5744
rect 19302 5680 19318 5744
rect 19382 5680 19398 5744
rect 19462 5680 19478 5744
rect 19542 5680 19558 5744
rect 19622 5680 19638 5744
rect 19702 5680 19718 5744
rect 19782 5680 19820 5744
rect 19200 5664 19820 5680
rect 23197 5288 23263 5291
rect 23197 5286 28796 5288
rect 23197 5230 23202 5286
rect 23258 5230 28796 5286
rect 23197 5228 28796 5230
rect 23197 5225 23263 5228
rect 26233 2726 26299 2729
rect 26233 2724 28796 2726
rect 26233 2668 26238 2724
rect 26294 2668 28796 2724
rect 26233 2666 28796 2668
rect 26233 2663 26299 2666
rect 28717 408 28783 411
rect 28352 406 28783 408
rect 28352 350 28722 406
rect 28778 350 28783 406
rect 28352 348 28783 350
rect 14273 164 14339 167
rect 28352 164 28412 348
rect 28717 345 28783 348
rect 14273 162 28412 164
rect 14273 106 14278 162
rect 14334 106 28412 162
rect 14273 104 28412 106
rect 28533 164 28599 167
rect 28533 162 28796 164
rect 28533 106 28538 162
rect 28594 106 28796 162
rect 28533 104 28796 106
rect 14273 101 14339 104
rect 28533 101 28599 104
<< via3 >>
rect 8038 22060 8102 22064
rect 8038 22004 8042 22060
rect 8042 22004 8098 22060
rect 8098 22004 8102 22060
rect 8038 22000 8102 22004
rect 8118 22060 8182 22064
rect 8118 22004 8122 22060
rect 8122 22004 8178 22060
rect 8178 22004 8182 22060
rect 8118 22000 8182 22004
rect 8198 22060 8262 22064
rect 8198 22004 8202 22060
rect 8202 22004 8258 22060
rect 8258 22004 8262 22060
rect 8198 22000 8262 22004
rect 8278 22060 8342 22064
rect 8278 22004 8282 22060
rect 8282 22004 8338 22060
rect 8338 22004 8342 22060
rect 8278 22000 8342 22004
rect 8358 22060 8422 22064
rect 8358 22004 8362 22060
rect 8362 22004 8418 22060
rect 8418 22004 8422 22060
rect 8358 22000 8422 22004
rect 8438 22060 8502 22064
rect 8438 22004 8442 22060
rect 8442 22004 8498 22060
rect 8498 22004 8502 22060
rect 8438 22000 8502 22004
rect 8518 22060 8582 22064
rect 8518 22004 8522 22060
rect 8522 22004 8578 22060
rect 8578 22004 8582 22060
rect 8518 22000 8582 22004
rect 13638 22060 13702 22064
rect 13638 22004 13642 22060
rect 13642 22004 13698 22060
rect 13698 22004 13702 22060
rect 13638 22000 13702 22004
rect 13718 22060 13782 22064
rect 13718 22004 13722 22060
rect 13722 22004 13778 22060
rect 13778 22004 13782 22060
rect 13718 22000 13782 22004
rect 13798 22060 13862 22064
rect 13798 22004 13802 22060
rect 13802 22004 13858 22060
rect 13858 22004 13862 22060
rect 13798 22000 13862 22004
rect 13878 22060 13942 22064
rect 13878 22004 13882 22060
rect 13882 22004 13938 22060
rect 13938 22004 13942 22060
rect 13878 22000 13942 22004
rect 13958 22060 14022 22064
rect 13958 22004 13962 22060
rect 13962 22004 14018 22060
rect 14018 22004 14022 22060
rect 13958 22000 14022 22004
rect 14038 22060 14102 22064
rect 14038 22004 14042 22060
rect 14042 22004 14098 22060
rect 14098 22004 14102 22060
rect 14038 22000 14102 22004
rect 14118 22060 14182 22064
rect 14118 22004 14122 22060
rect 14122 22004 14178 22060
rect 14178 22004 14182 22060
rect 14118 22000 14182 22004
rect 19238 22060 19302 22064
rect 19238 22004 19242 22060
rect 19242 22004 19298 22060
rect 19298 22004 19302 22060
rect 19238 22000 19302 22004
rect 19318 22060 19382 22064
rect 19318 22004 19322 22060
rect 19322 22004 19378 22060
rect 19378 22004 19382 22060
rect 19318 22000 19382 22004
rect 19398 22060 19462 22064
rect 19398 22004 19402 22060
rect 19402 22004 19458 22060
rect 19458 22004 19462 22060
rect 19398 22000 19462 22004
rect 19478 22060 19542 22064
rect 19478 22004 19482 22060
rect 19482 22004 19538 22060
rect 19538 22004 19542 22060
rect 19478 22000 19542 22004
rect 19558 22060 19622 22064
rect 19558 22004 19562 22060
rect 19562 22004 19618 22060
rect 19618 22004 19622 22060
rect 19558 22000 19622 22004
rect 19638 22060 19702 22064
rect 19638 22004 19642 22060
rect 19642 22004 19698 22060
rect 19698 22004 19702 22060
rect 19638 22000 19702 22004
rect 19718 22060 19782 22064
rect 19718 22004 19722 22060
rect 19722 22004 19778 22060
rect 19778 22004 19782 22060
rect 19718 22000 19782 22004
rect 9278 21516 9342 21520
rect 9278 21460 9282 21516
rect 9282 21460 9338 21516
rect 9338 21460 9342 21516
rect 9278 21456 9342 21460
rect 9358 21516 9422 21520
rect 9358 21460 9362 21516
rect 9362 21460 9418 21516
rect 9418 21460 9422 21516
rect 9358 21456 9422 21460
rect 9438 21516 9502 21520
rect 9438 21460 9442 21516
rect 9442 21460 9498 21516
rect 9498 21460 9502 21516
rect 9438 21456 9502 21460
rect 9518 21516 9582 21520
rect 9518 21460 9522 21516
rect 9522 21460 9578 21516
rect 9578 21460 9582 21516
rect 9518 21456 9582 21460
rect 9598 21516 9662 21520
rect 9598 21460 9602 21516
rect 9602 21460 9658 21516
rect 9658 21460 9662 21516
rect 9598 21456 9662 21460
rect 9678 21516 9742 21520
rect 9678 21460 9682 21516
rect 9682 21460 9738 21516
rect 9738 21460 9742 21516
rect 9678 21456 9742 21460
rect 9758 21516 9822 21520
rect 9758 21460 9762 21516
rect 9762 21460 9818 21516
rect 9818 21460 9822 21516
rect 9758 21456 9822 21460
rect 14878 21516 14942 21520
rect 14878 21460 14882 21516
rect 14882 21460 14938 21516
rect 14938 21460 14942 21516
rect 14878 21456 14942 21460
rect 14958 21516 15022 21520
rect 14958 21460 14962 21516
rect 14962 21460 15018 21516
rect 15018 21460 15022 21516
rect 14958 21456 15022 21460
rect 15038 21516 15102 21520
rect 15038 21460 15042 21516
rect 15042 21460 15098 21516
rect 15098 21460 15102 21516
rect 15038 21456 15102 21460
rect 15118 21516 15182 21520
rect 15118 21460 15122 21516
rect 15122 21460 15178 21516
rect 15178 21460 15182 21516
rect 15118 21456 15182 21460
rect 15198 21516 15262 21520
rect 15198 21460 15202 21516
rect 15202 21460 15258 21516
rect 15258 21460 15262 21516
rect 15198 21456 15262 21460
rect 15278 21516 15342 21520
rect 15278 21460 15282 21516
rect 15282 21460 15338 21516
rect 15338 21460 15342 21516
rect 15278 21456 15342 21460
rect 15358 21516 15422 21520
rect 15358 21460 15362 21516
rect 15362 21460 15418 21516
rect 15418 21460 15422 21516
rect 15358 21456 15422 21460
rect 20478 21516 20542 21520
rect 20478 21460 20482 21516
rect 20482 21460 20538 21516
rect 20538 21460 20542 21516
rect 20478 21456 20542 21460
rect 20558 21516 20622 21520
rect 20558 21460 20562 21516
rect 20562 21460 20618 21516
rect 20618 21460 20622 21516
rect 20558 21456 20622 21460
rect 20638 21516 20702 21520
rect 20638 21460 20642 21516
rect 20642 21460 20698 21516
rect 20698 21460 20702 21516
rect 20638 21456 20702 21460
rect 20718 21516 20782 21520
rect 20718 21460 20722 21516
rect 20722 21460 20778 21516
rect 20778 21460 20782 21516
rect 20718 21456 20782 21460
rect 20798 21516 20862 21520
rect 20798 21460 20802 21516
rect 20802 21460 20858 21516
rect 20858 21460 20862 21516
rect 20798 21456 20862 21460
rect 20878 21516 20942 21520
rect 20878 21460 20882 21516
rect 20882 21460 20938 21516
rect 20938 21460 20942 21516
rect 20878 21456 20942 21460
rect 20958 21516 21022 21520
rect 20958 21460 20962 21516
rect 20962 21460 21018 21516
rect 21018 21460 21022 21516
rect 20958 21456 21022 21460
rect 8038 20972 8102 20976
rect 8038 20916 8042 20972
rect 8042 20916 8098 20972
rect 8098 20916 8102 20972
rect 8038 20912 8102 20916
rect 8118 20972 8182 20976
rect 8118 20916 8122 20972
rect 8122 20916 8178 20972
rect 8178 20916 8182 20972
rect 8118 20912 8182 20916
rect 8198 20972 8262 20976
rect 8198 20916 8202 20972
rect 8202 20916 8258 20972
rect 8258 20916 8262 20972
rect 8198 20912 8262 20916
rect 8278 20972 8342 20976
rect 8278 20916 8282 20972
rect 8282 20916 8338 20972
rect 8338 20916 8342 20972
rect 8278 20912 8342 20916
rect 8358 20972 8422 20976
rect 8358 20916 8362 20972
rect 8362 20916 8418 20972
rect 8418 20916 8422 20972
rect 8358 20912 8422 20916
rect 8438 20972 8502 20976
rect 8438 20916 8442 20972
rect 8442 20916 8498 20972
rect 8498 20916 8502 20972
rect 8438 20912 8502 20916
rect 8518 20972 8582 20976
rect 8518 20916 8522 20972
rect 8522 20916 8578 20972
rect 8578 20916 8582 20972
rect 8518 20912 8582 20916
rect 13638 20972 13702 20976
rect 13638 20916 13642 20972
rect 13642 20916 13698 20972
rect 13698 20916 13702 20972
rect 13638 20912 13702 20916
rect 13718 20972 13782 20976
rect 13718 20916 13722 20972
rect 13722 20916 13778 20972
rect 13778 20916 13782 20972
rect 13718 20912 13782 20916
rect 13798 20972 13862 20976
rect 13798 20916 13802 20972
rect 13802 20916 13858 20972
rect 13858 20916 13862 20972
rect 13798 20912 13862 20916
rect 13878 20972 13942 20976
rect 13878 20916 13882 20972
rect 13882 20916 13938 20972
rect 13938 20916 13942 20972
rect 13878 20912 13942 20916
rect 13958 20972 14022 20976
rect 13958 20916 13962 20972
rect 13962 20916 14018 20972
rect 14018 20916 14022 20972
rect 13958 20912 14022 20916
rect 14038 20972 14102 20976
rect 14038 20916 14042 20972
rect 14042 20916 14098 20972
rect 14098 20916 14102 20972
rect 14038 20912 14102 20916
rect 14118 20972 14182 20976
rect 14118 20916 14122 20972
rect 14122 20916 14178 20972
rect 14178 20916 14182 20972
rect 14118 20912 14182 20916
rect 19238 20972 19302 20976
rect 19238 20916 19242 20972
rect 19242 20916 19298 20972
rect 19298 20916 19302 20972
rect 19238 20912 19302 20916
rect 19318 20972 19382 20976
rect 19318 20916 19322 20972
rect 19322 20916 19378 20972
rect 19378 20916 19382 20972
rect 19318 20912 19382 20916
rect 19398 20972 19462 20976
rect 19398 20916 19402 20972
rect 19402 20916 19458 20972
rect 19458 20916 19462 20972
rect 19398 20912 19462 20916
rect 19478 20972 19542 20976
rect 19478 20916 19482 20972
rect 19482 20916 19538 20972
rect 19538 20916 19542 20972
rect 19478 20912 19542 20916
rect 19558 20972 19622 20976
rect 19558 20916 19562 20972
rect 19562 20916 19618 20972
rect 19618 20916 19622 20972
rect 19558 20912 19622 20916
rect 19638 20972 19702 20976
rect 19638 20916 19642 20972
rect 19642 20916 19698 20972
rect 19698 20916 19702 20972
rect 19638 20912 19702 20916
rect 19718 20972 19782 20976
rect 19718 20916 19722 20972
rect 19722 20916 19778 20972
rect 19778 20916 19782 20972
rect 19718 20912 19782 20916
rect 9278 20428 9342 20432
rect 9278 20372 9282 20428
rect 9282 20372 9338 20428
rect 9338 20372 9342 20428
rect 9278 20368 9342 20372
rect 9358 20428 9422 20432
rect 9358 20372 9362 20428
rect 9362 20372 9418 20428
rect 9418 20372 9422 20428
rect 9358 20368 9422 20372
rect 9438 20428 9502 20432
rect 9438 20372 9442 20428
rect 9442 20372 9498 20428
rect 9498 20372 9502 20428
rect 9438 20368 9502 20372
rect 9518 20428 9582 20432
rect 9518 20372 9522 20428
rect 9522 20372 9578 20428
rect 9578 20372 9582 20428
rect 9518 20368 9582 20372
rect 9598 20428 9662 20432
rect 9598 20372 9602 20428
rect 9602 20372 9658 20428
rect 9658 20372 9662 20428
rect 9598 20368 9662 20372
rect 9678 20428 9742 20432
rect 9678 20372 9682 20428
rect 9682 20372 9738 20428
rect 9738 20372 9742 20428
rect 9678 20368 9742 20372
rect 9758 20428 9822 20432
rect 9758 20372 9762 20428
rect 9762 20372 9818 20428
rect 9818 20372 9822 20428
rect 9758 20368 9822 20372
rect 14878 20428 14942 20432
rect 14878 20372 14882 20428
rect 14882 20372 14938 20428
rect 14938 20372 14942 20428
rect 14878 20368 14942 20372
rect 14958 20428 15022 20432
rect 14958 20372 14962 20428
rect 14962 20372 15018 20428
rect 15018 20372 15022 20428
rect 14958 20368 15022 20372
rect 15038 20428 15102 20432
rect 15038 20372 15042 20428
rect 15042 20372 15098 20428
rect 15098 20372 15102 20428
rect 15038 20368 15102 20372
rect 15118 20428 15182 20432
rect 15118 20372 15122 20428
rect 15122 20372 15178 20428
rect 15178 20372 15182 20428
rect 15118 20368 15182 20372
rect 15198 20428 15262 20432
rect 15198 20372 15202 20428
rect 15202 20372 15258 20428
rect 15258 20372 15262 20428
rect 15198 20368 15262 20372
rect 15278 20428 15342 20432
rect 15278 20372 15282 20428
rect 15282 20372 15338 20428
rect 15338 20372 15342 20428
rect 15278 20368 15342 20372
rect 15358 20428 15422 20432
rect 15358 20372 15362 20428
rect 15362 20372 15418 20428
rect 15418 20372 15422 20428
rect 15358 20368 15422 20372
rect 20478 20428 20542 20432
rect 20478 20372 20482 20428
rect 20482 20372 20538 20428
rect 20538 20372 20542 20428
rect 20478 20368 20542 20372
rect 20558 20428 20622 20432
rect 20558 20372 20562 20428
rect 20562 20372 20618 20428
rect 20618 20372 20622 20428
rect 20558 20368 20622 20372
rect 20638 20428 20702 20432
rect 20638 20372 20642 20428
rect 20642 20372 20698 20428
rect 20698 20372 20702 20428
rect 20638 20368 20702 20372
rect 20718 20428 20782 20432
rect 20718 20372 20722 20428
rect 20722 20372 20778 20428
rect 20778 20372 20782 20428
rect 20718 20368 20782 20372
rect 20798 20428 20862 20432
rect 20798 20372 20802 20428
rect 20802 20372 20858 20428
rect 20858 20372 20862 20428
rect 20798 20368 20862 20372
rect 20878 20428 20942 20432
rect 20878 20372 20882 20428
rect 20882 20372 20938 20428
rect 20938 20372 20942 20428
rect 20878 20368 20942 20372
rect 20958 20428 21022 20432
rect 20958 20372 20962 20428
rect 20962 20372 21018 20428
rect 21018 20372 21022 20428
rect 20958 20368 21022 20372
rect 8038 19884 8102 19888
rect 8038 19828 8042 19884
rect 8042 19828 8098 19884
rect 8098 19828 8102 19884
rect 8038 19824 8102 19828
rect 8118 19884 8182 19888
rect 8118 19828 8122 19884
rect 8122 19828 8178 19884
rect 8178 19828 8182 19884
rect 8118 19824 8182 19828
rect 8198 19884 8262 19888
rect 8198 19828 8202 19884
rect 8202 19828 8258 19884
rect 8258 19828 8262 19884
rect 8198 19824 8262 19828
rect 8278 19884 8342 19888
rect 8278 19828 8282 19884
rect 8282 19828 8338 19884
rect 8338 19828 8342 19884
rect 8278 19824 8342 19828
rect 8358 19884 8422 19888
rect 8358 19828 8362 19884
rect 8362 19828 8418 19884
rect 8418 19828 8422 19884
rect 8358 19824 8422 19828
rect 8438 19884 8502 19888
rect 8438 19828 8442 19884
rect 8442 19828 8498 19884
rect 8498 19828 8502 19884
rect 8438 19824 8502 19828
rect 8518 19884 8582 19888
rect 8518 19828 8522 19884
rect 8522 19828 8578 19884
rect 8578 19828 8582 19884
rect 8518 19824 8582 19828
rect 13638 19884 13702 19888
rect 13638 19828 13642 19884
rect 13642 19828 13698 19884
rect 13698 19828 13702 19884
rect 13638 19824 13702 19828
rect 13718 19884 13782 19888
rect 13718 19828 13722 19884
rect 13722 19828 13778 19884
rect 13778 19828 13782 19884
rect 13718 19824 13782 19828
rect 13798 19884 13862 19888
rect 13798 19828 13802 19884
rect 13802 19828 13858 19884
rect 13858 19828 13862 19884
rect 13798 19824 13862 19828
rect 13878 19884 13942 19888
rect 13878 19828 13882 19884
rect 13882 19828 13938 19884
rect 13938 19828 13942 19884
rect 13878 19824 13942 19828
rect 13958 19884 14022 19888
rect 13958 19828 13962 19884
rect 13962 19828 14018 19884
rect 14018 19828 14022 19884
rect 13958 19824 14022 19828
rect 14038 19884 14102 19888
rect 14038 19828 14042 19884
rect 14042 19828 14098 19884
rect 14098 19828 14102 19884
rect 14038 19824 14102 19828
rect 14118 19884 14182 19888
rect 14118 19828 14122 19884
rect 14122 19828 14178 19884
rect 14178 19828 14182 19884
rect 14118 19824 14182 19828
rect 19238 19884 19302 19888
rect 19238 19828 19242 19884
rect 19242 19828 19298 19884
rect 19298 19828 19302 19884
rect 19238 19824 19302 19828
rect 19318 19884 19382 19888
rect 19318 19828 19322 19884
rect 19322 19828 19378 19884
rect 19378 19828 19382 19884
rect 19318 19824 19382 19828
rect 19398 19884 19462 19888
rect 19398 19828 19402 19884
rect 19402 19828 19458 19884
rect 19458 19828 19462 19884
rect 19398 19824 19462 19828
rect 19478 19884 19542 19888
rect 19478 19828 19482 19884
rect 19482 19828 19538 19884
rect 19538 19828 19542 19884
rect 19478 19824 19542 19828
rect 19558 19884 19622 19888
rect 19558 19828 19562 19884
rect 19562 19828 19618 19884
rect 19618 19828 19622 19884
rect 19558 19824 19622 19828
rect 19638 19884 19702 19888
rect 19638 19828 19642 19884
rect 19642 19828 19698 19884
rect 19698 19828 19702 19884
rect 19638 19824 19702 19828
rect 19718 19884 19782 19888
rect 19718 19828 19722 19884
rect 19722 19828 19778 19884
rect 19778 19828 19782 19884
rect 19718 19824 19782 19828
rect 9278 19340 9342 19344
rect 9278 19284 9282 19340
rect 9282 19284 9338 19340
rect 9338 19284 9342 19340
rect 9278 19280 9342 19284
rect 9358 19340 9422 19344
rect 9358 19284 9362 19340
rect 9362 19284 9418 19340
rect 9418 19284 9422 19340
rect 9358 19280 9422 19284
rect 9438 19340 9502 19344
rect 9438 19284 9442 19340
rect 9442 19284 9498 19340
rect 9498 19284 9502 19340
rect 9438 19280 9502 19284
rect 9518 19340 9582 19344
rect 9518 19284 9522 19340
rect 9522 19284 9578 19340
rect 9578 19284 9582 19340
rect 9518 19280 9582 19284
rect 9598 19340 9662 19344
rect 9598 19284 9602 19340
rect 9602 19284 9658 19340
rect 9658 19284 9662 19340
rect 9598 19280 9662 19284
rect 9678 19340 9742 19344
rect 9678 19284 9682 19340
rect 9682 19284 9738 19340
rect 9738 19284 9742 19340
rect 9678 19280 9742 19284
rect 9758 19340 9822 19344
rect 9758 19284 9762 19340
rect 9762 19284 9818 19340
rect 9818 19284 9822 19340
rect 9758 19280 9822 19284
rect 14878 19340 14942 19344
rect 14878 19284 14882 19340
rect 14882 19284 14938 19340
rect 14938 19284 14942 19340
rect 14878 19280 14942 19284
rect 14958 19340 15022 19344
rect 14958 19284 14962 19340
rect 14962 19284 15018 19340
rect 15018 19284 15022 19340
rect 14958 19280 15022 19284
rect 15038 19340 15102 19344
rect 15038 19284 15042 19340
rect 15042 19284 15098 19340
rect 15098 19284 15102 19340
rect 15038 19280 15102 19284
rect 15118 19340 15182 19344
rect 15118 19284 15122 19340
rect 15122 19284 15178 19340
rect 15178 19284 15182 19340
rect 15118 19280 15182 19284
rect 15198 19340 15262 19344
rect 15198 19284 15202 19340
rect 15202 19284 15258 19340
rect 15258 19284 15262 19340
rect 15198 19280 15262 19284
rect 15278 19340 15342 19344
rect 15278 19284 15282 19340
rect 15282 19284 15338 19340
rect 15338 19284 15342 19340
rect 15278 19280 15342 19284
rect 15358 19340 15422 19344
rect 15358 19284 15362 19340
rect 15362 19284 15418 19340
rect 15418 19284 15422 19340
rect 15358 19280 15422 19284
rect 20478 19340 20542 19344
rect 20478 19284 20482 19340
rect 20482 19284 20538 19340
rect 20538 19284 20542 19340
rect 20478 19280 20542 19284
rect 20558 19340 20622 19344
rect 20558 19284 20562 19340
rect 20562 19284 20618 19340
rect 20618 19284 20622 19340
rect 20558 19280 20622 19284
rect 20638 19340 20702 19344
rect 20638 19284 20642 19340
rect 20642 19284 20698 19340
rect 20698 19284 20702 19340
rect 20638 19280 20702 19284
rect 20718 19340 20782 19344
rect 20718 19284 20722 19340
rect 20722 19284 20778 19340
rect 20778 19284 20782 19340
rect 20718 19280 20782 19284
rect 20798 19340 20862 19344
rect 20798 19284 20802 19340
rect 20802 19284 20858 19340
rect 20858 19284 20862 19340
rect 20798 19280 20862 19284
rect 20878 19340 20942 19344
rect 20878 19284 20882 19340
rect 20882 19284 20938 19340
rect 20938 19284 20942 19340
rect 20878 19280 20942 19284
rect 20958 19340 21022 19344
rect 20958 19284 20962 19340
rect 20962 19284 21018 19340
rect 21018 19284 21022 19340
rect 20958 19280 21022 19284
rect 8038 18796 8102 18800
rect 8038 18740 8042 18796
rect 8042 18740 8098 18796
rect 8098 18740 8102 18796
rect 8038 18736 8102 18740
rect 8118 18796 8182 18800
rect 8118 18740 8122 18796
rect 8122 18740 8178 18796
rect 8178 18740 8182 18796
rect 8118 18736 8182 18740
rect 8198 18796 8262 18800
rect 8198 18740 8202 18796
rect 8202 18740 8258 18796
rect 8258 18740 8262 18796
rect 8198 18736 8262 18740
rect 8278 18796 8342 18800
rect 8278 18740 8282 18796
rect 8282 18740 8338 18796
rect 8338 18740 8342 18796
rect 8278 18736 8342 18740
rect 8358 18796 8422 18800
rect 8358 18740 8362 18796
rect 8362 18740 8418 18796
rect 8418 18740 8422 18796
rect 8358 18736 8422 18740
rect 8438 18796 8502 18800
rect 8438 18740 8442 18796
rect 8442 18740 8498 18796
rect 8498 18740 8502 18796
rect 8438 18736 8502 18740
rect 8518 18796 8582 18800
rect 8518 18740 8522 18796
rect 8522 18740 8578 18796
rect 8578 18740 8582 18796
rect 8518 18736 8582 18740
rect 13638 18796 13702 18800
rect 13638 18740 13642 18796
rect 13642 18740 13698 18796
rect 13698 18740 13702 18796
rect 13638 18736 13702 18740
rect 13718 18796 13782 18800
rect 13718 18740 13722 18796
rect 13722 18740 13778 18796
rect 13778 18740 13782 18796
rect 13718 18736 13782 18740
rect 13798 18796 13862 18800
rect 13798 18740 13802 18796
rect 13802 18740 13858 18796
rect 13858 18740 13862 18796
rect 13798 18736 13862 18740
rect 13878 18796 13942 18800
rect 13878 18740 13882 18796
rect 13882 18740 13938 18796
rect 13938 18740 13942 18796
rect 13878 18736 13942 18740
rect 13958 18796 14022 18800
rect 13958 18740 13962 18796
rect 13962 18740 14018 18796
rect 14018 18740 14022 18796
rect 13958 18736 14022 18740
rect 14038 18796 14102 18800
rect 14038 18740 14042 18796
rect 14042 18740 14098 18796
rect 14098 18740 14102 18796
rect 14038 18736 14102 18740
rect 14118 18796 14182 18800
rect 14118 18740 14122 18796
rect 14122 18740 14178 18796
rect 14178 18740 14182 18796
rect 14118 18736 14182 18740
rect 19238 18796 19302 18800
rect 19238 18740 19242 18796
rect 19242 18740 19298 18796
rect 19298 18740 19302 18796
rect 19238 18736 19302 18740
rect 19318 18796 19382 18800
rect 19318 18740 19322 18796
rect 19322 18740 19378 18796
rect 19378 18740 19382 18796
rect 19318 18736 19382 18740
rect 19398 18796 19462 18800
rect 19398 18740 19402 18796
rect 19402 18740 19458 18796
rect 19458 18740 19462 18796
rect 19398 18736 19462 18740
rect 19478 18796 19542 18800
rect 19478 18740 19482 18796
rect 19482 18740 19538 18796
rect 19538 18740 19542 18796
rect 19478 18736 19542 18740
rect 19558 18796 19622 18800
rect 19558 18740 19562 18796
rect 19562 18740 19618 18796
rect 19618 18740 19622 18796
rect 19558 18736 19622 18740
rect 19638 18796 19702 18800
rect 19638 18740 19642 18796
rect 19642 18740 19698 18796
rect 19698 18740 19702 18796
rect 19638 18736 19702 18740
rect 19718 18796 19782 18800
rect 19718 18740 19722 18796
rect 19722 18740 19778 18796
rect 19778 18740 19782 18796
rect 19718 18736 19782 18740
rect 9278 18252 9342 18256
rect 9278 18196 9282 18252
rect 9282 18196 9338 18252
rect 9338 18196 9342 18252
rect 9278 18192 9342 18196
rect 9358 18252 9422 18256
rect 9358 18196 9362 18252
rect 9362 18196 9418 18252
rect 9418 18196 9422 18252
rect 9358 18192 9422 18196
rect 9438 18252 9502 18256
rect 9438 18196 9442 18252
rect 9442 18196 9498 18252
rect 9498 18196 9502 18252
rect 9438 18192 9502 18196
rect 9518 18252 9582 18256
rect 9518 18196 9522 18252
rect 9522 18196 9578 18252
rect 9578 18196 9582 18252
rect 9518 18192 9582 18196
rect 9598 18252 9662 18256
rect 9598 18196 9602 18252
rect 9602 18196 9658 18252
rect 9658 18196 9662 18252
rect 9598 18192 9662 18196
rect 9678 18252 9742 18256
rect 9678 18196 9682 18252
rect 9682 18196 9738 18252
rect 9738 18196 9742 18252
rect 9678 18192 9742 18196
rect 9758 18252 9822 18256
rect 9758 18196 9762 18252
rect 9762 18196 9818 18252
rect 9818 18196 9822 18252
rect 9758 18192 9822 18196
rect 14878 18252 14942 18256
rect 14878 18196 14882 18252
rect 14882 18196 14938 18252
rect 14938 18196 14942 18252
rect 14878 18192 14942 18196
rect 14958 18252 15022 18256
rect 14958 18196 14962 18252
rect 14962 18196 15018 18252
rect 15018 18196 15022 18252
rect 14958 18192 15022 18196
rect 15038 18252 15102 18256
rect 15038 18196 15042 18252
rect 15042 18196 15098 18252
rect 15098 18196 15102 18252
rect 15038 18192 15102 18196
rect 15118 18252 15182 18256
rect 15118 18196 15122 18252
rect 15122 18196 15178 18252
rect 15178 18196 15182 18252
rect 15118 18192 15182 18196
rect 15198 18252 15262 18256
rect 15198 18196 15202 18252
rect 15202 18196 15258 18252
rect 15258 18196 15262 18252
rect 15198 18192 15262 18196
rect 15278 18252 15342 18256
rect 15278 18196 15282 18252
rect 15282 18196 15338 18252
rect 15338 18196 15342 18252
rect 15278 18192 15342 18196
rect 15358 18252 15422 18256
rect 15358 18196 15362 18252
rect 15362 18196 15418 18252
rect 15418 18196 15422 18252
rect 15358 18192 15422 18196
rect 20478 18252 20542 18256
rect 20478 18196 20482 18252
rect 20482 18196 20538 18252
rect 20538 18196 20542 18252
rect 20478 18192 20542 18196
rect 20558 18252 20622 18256
rect 20558 18196 20562 18252
rect 20562 18196 20618 18252
rect 20618 18196 20622 18252
rect 20558 18192 20622 18196
rect 20638 18252 20702 18256
rect 20638 18196 20642 18252
rect 20642 18196 20698 18252
rect 20698 18196 20702 18252
rect 20638 18192 20702 18196
rect 20718 18252 20782 18256
rect 20718 18196 20722 18252
rect 20722 18196 20778 18252
rect 20778 18196 20782 18252
rect 20718 18192 20782 18196
rect 20798 18252 20862 18256
rect 20798 18196 20802 18252
rect 20802 18196 20858 18252
rect 20858 18196 20862 18252
rect 20798 18192 20862 18196
rect 20878 18252 20942 18256
rect 20878 18196 20882 18252
rect 20882 18196 20938 18252
rect 20938 18196 20942 18252
rect 20878 18192 20942 18196
rect 20958 18252 21022 18256
rect 20958 18196 20962 18252
rect 20962 18196 21018 18252
rect 21018 18196 21022 18252
rect 20958 18192 21022 18196
rect 8038 17708 8102 17712
rect 8038 17652 8042 17708
rect 8042 17652 8098 17708
rect 8098 17652 8102 17708
rect 8038 17648 8102 17652
rect 8118 17708 8182 17712
rect 8118 17652 8122 17708
rect 8122 17652 8178 17708
rect 8178 17652 8182 17708
rect 8118 17648 8182 17652
rect 8198 17708 8262 17712
rect 8198 17652 8202 17708
rect 8202 17652 8258 17708
rect 8258 17652 8262 17708
rect 8198 17648 8262 17652
rect 8278 17708 8342 17712
rect 8278 17652 8282 17708
rect 8282 17652 8338 17708
rect 8338 17652 8342 17708
rect 8278 17648 8342 17652
rect 8358 17708 8422 17712
rect 8358 17652 8362 17708
rect 8362 17652 8418 17708
rect 8418 17652 8422 17708
rect 8358 17648 8422 17652
rect 8438 17708 8502 17712
rect 8438 17652 8442 17708
rect 8442 17652 8498 17708
rect 8498 17652 8502 17708
rect 8438 17648 8502 17652
rect 8518 17708 8582 17712
rect 8518 17652 8522 17708
rect 8522 17652 8578 17708
rect 8578 17652 8582 17708
rect 8518 17648 8582 17652
rect 13638 17708 13702 17712
rect 13638 17652 13642 17708
rect 13642 17652 13698 17708
rect 13698 17652 13702 17708
rect 13638 17648 13702 17652
rect 13718 17708 13782 17712
rect 13718 17652 13722 17708
rect 13722 17652 13778 17708
rect 13778 17652 13782 17708
rect 13718 17648 13782 17652
rect 13798 17708 13862 17712
rect 13798 17652 13802 17708
rect 13802 17652 13858 17708
rect 13858 17652 13862 17708
rect 13798 17648 13862 17652
rect 13878 17708 13942 17712
rect 13878 17652 13882 17708
rect 13882 17652 13938 17708
rect 13938 17652 13942 17708
rect 13878 17648 13942 17652
rect 13958 17708 14022 17712
rect 13958 17652 13962 17708
rect 13962 17652 14018 17708
rect 14018 17652 14022 17708
rect 13958 17648 14022 17652
rect 14038 17708 14102 17712
rect 14038 17652 14042 17708
rect 14042 17652 14098 17708
rect 14098 17652 14102 17708
rect 14038 17648 14102 17652
rect 14118 17708 14182 17712
rect 14118 17652 14122 17708
rect 14122 17652 14178 17708
rect 14178 17652 14182 17708
rect 14118 17648 14182 17652
rect 19238 17708 19302 17712
rect 19238 17652 19242 17708
rect 19242 17652 19298 17708
rect 19298 17652 19302 17708
rect 19238 17648 19302 17652
rect 19318 17708 19382 17712
rect 19318 17652 19322 17708
rect 19322 17652 19378 17708
rect 19378 17652 19382 17708
rect 19318 17648 19382 17652
rect 19398 17708 19462 17712
rect 19398 17652 19402 17708
rect 19402 17652 19458 17708
rect 19458 17652 19462 17708
rect 19398 17648 19462 17652
rect 19478 17708 19542 17712
rect 19478 17652 19482 17708
rect 19482 17652 19538 17708
rect 19538 17652 19542 17708
rect 19478 17648 19542 17652
rect 19558 17708 19622 17712
rect 19558 17652 19562 17708
rect 19562 17652 19618 17708
rect 19618 17652 19622 17708
rect 19558 17648 19622 17652
rect 19638 17708 19702 17712
rect 19638 17652 19642 17708
rect 19642 17652 19698 17708
rect 19698 17652 19702 17708
rect 19638 17648 19702 17652
rect 19718 17708 19782 17712
rect 19718 17652 19722 17708
rect 19722 17652 19778 17708
rect 19778 17652 19782 17708
rect 19718 17648 19782 17652
rect 9278 17164 9342 17168
rect 9278 17108 9282 17164
rect 9282 17108 9338 17164
rect 9338 17108 9342 17164
rect 9278 17104 9342 17108
rect 9358 17164 9422 17168
rect 9358 17108 9362 17164
rect 9362 17108 9418 17164
rect 9418 17108 9422 17164
rect 9358 17104 9422 17108
rect 9438 17164 9502 17168
rect 9438 17108 9442 17164
rect 9442 17108 9498 17164
rect 9498 17108 9502 17164
rect 9438 17104 9502 17108
rect 9518 17164 9582 17168
rect 9518 17108 9522 17164
rect 9522 17108 9578 17164
rect 9578 17108 9582 17164
rect 9518 17104 9582 17108
rect 9598 17164 9662 17168
rect 9598 17108 9602 17164
rect 9602 17108 9658 17164
rect 9658 17108 9662 17164
rect 9598 17104 9662 17108
rect 9678 17164 9742 17168
rect 9678 17108 9682 17164
rect 9682 17108 9738 17164
rect 9738 17108 9742 17164
rect 9678 17104 9742 17108
rect 9758 17164 9822 17168
rect 9758 17108 9762 17164
rect 9762 17108 9818 17164
rect 9818 17108 9822 17164
rect 9758 17104 9822 17108
rect 14878 17164 14942 17168
rect 14878 17108 14882 17164
rect 14882 17108 14938 17164
rect 14938 17108 14942 17164
rect 14878 17104 14942 17108
rect 14958 17164 15022 17168
rect 14958 17108 14962 17164
rect 14962 17108 15018 17164
rect 15018 17108 15022 17164
rect 14958 17104 15022 17108
rect 15038 17164 15102 17168
rect 15038 17108 15042 17164
rect 15042 17108 15098 17164
rect 15098 17108 15102 17164
rect 15038 17104 15102 17108
rect 15118 17164 15182 17168
rect 15118 17108 15122 17164
rect 15122 17108 15178 17164
rect 15178 17108 15182 17164
rect 15118 17104 15182 17108
rect 15198 17164 15262 17168
rect 15198 17108 15202 17164
rect 15202 17108 15258 17164
rect 15258 17108 15262 17164
rect 15198 17104 15262 17108
rect 15278 17164 15342 17168
rect 15278 17108 15282 17164
rect 15282 17108 15338 17164
rect 15338 17108 15342 17164
rect 15278 17104 15342 17108
rect 15358 17164 15422 17168
rect 15358 17108 15362 17164
rect 15362 17108 15418 17164
rect 15418 17108 15422 17164
rect 15358 17104 15422 17108
rect 20478 17164 20542 17168
rect 20478 17108 20482 17164
rect 20482 17108 20538 17164
rect 20538 17108 20542 17164
rect 20478 17104 20542 17108
rect 20558 17164 20622 17168
rect 20558 17108 20562 17164
rect 20562 17108 20618 17164
rect 20618 17108 20622 17164
rect 20558 17104 20622 17108
rect 20638 17164 20702 17168
rect 20638 17108 20642 17164
rect 20642 17108 20698 17164
rect 20698 17108 20702 17164
rect 20638 17104 20702 17108
rect 20718 17164 20782 17168
rect 20718 17108 20722 17164
rect 20722 17108 20778 17164
rect 20778 17108 20782 17164
rect 20718 17104 20782 17108
rect 20798 17164 20862 17168
rect 20798 17108 20802 17164
rect 20802 17108 20858 17164
rect 20858 17108 20862 17164
rect 20798 17104 20862 17108
rect 20878 17164 20942 17168
rect 20878 17108 20882 17164
rect 20882 17108 20938 17164
rect 20938 17108 20942 17164
rect 20878 17104 20942 17108
rect 20958 17164 21022 17168
rect 20958 17108 20962 17164
rect 20962 17108 21018 17164
rect 21018 17108 21022 17164
rect 20958 17104 21022 17108
rect 8038 16620 8102 16624
rect 8038 16564 8042 16620
rect 8042 16564 8098 16620
rect 8098 16564 8102 16620
rect 8038 16560 8102 16564
rect 8118 16620 8182 16624
rect 8118 16564 8122 16620
rect 8122 16564 8178 16620
rect 8178 16564 8182 16620
rect 8118 16560 8182 16564
rect 8198 16620 8262 16624
rect 8198 16564 8202 16620
rect 8202 16564 8258 16620
rect 8258 16564 8262 16620
rect 8198 16560 8262 16564
rect 8278 16620 8342 16624
rect 8278 16564 8282 16620
rect 8282 16564 8338 16620
rect 8338 16564 8342 16620
rect 8278 16560 8342 16564
rect 8358 16620 8422 16624
rect 8358 16564 8362 16620
rect 8362 16564 8418 16620
rect 8418 16564 8422 16620
rect 8358 16560 8422 16564
rect 8438 16620 8502 16624
rect 8438 16564 8442 16620
rect 8442 16564 8498 16620
rect 8498 16564 8502 16620
rect 8438 16560 8502 16564
rect 8518 16620 8582 16624
rect 8518 16564 8522 16620
rect 8522 16564 8578 16620
rect 8578 16564 8582 16620
rect 8518 16560 8582 16564
rect 13638 16620 13702 16624
rect 13638 16564 13642 16620
rect 13642 16564 13698 16620
rect 13698 16564 13702 16620
rect 13638 16560 13702 16564
rect 13718 16620 13782 16624
rect 13718 16564 13722 16620
rect 13722 16564 13778 16620
rect 13778 16564 13782 16620
rect 13718 16560 13782 16564
rect 13798 16620 13862 16624
rect 13798 16564 13802 16620
rect 13802 16564 13858 16620
rect 13858 16564 13862 16620
rect 13798 16560 13862 16564
rect 13878 16620 13942 16624
rect 13878 16564 13882 16620
rect 13882 16564 13938 16620
rect 13938 16564 13942 16620
rect 13878 16560 13942 16564
rect 13958 16620 14022 16624
rect 13958 16564 13962 16620
rect 13962 16564 14018 16620
rect 14018 16564 14022 16620
rect 13958 16560 14022 16564
rect 14038 16620 14102 16624
rect 14038 16564 14042 16620
rect 14042 16564 14098 16620
rect 14098 16564 14102 16620
rect 14038 16560 14102 16564
rect 14118 16620 14182 16624
rect 14118 16564 14122 16620
rect 14122 16564 14178 16620
rect 14178 16564 14182 16620
rect 14118 16560 14182 16564
rect 19238 16620 19302 16624
rect 19238 16564 19242 16620
rect 19242 16564 19298 16620
rect 19298 16564 19302 16620
rect 19238 16560 19302 16564
rect 19318 16620 19382 16624
rect 19318 16564 19322 16620
rect 19322 16564 19378 16620
rect 19378 16564 19382 16620
rect 19318 16560 19382 16564
rect 19398 16620 19462 16624
rect 19398 16564 19402 16620
rect 19402 16564 19458 16620
rect 19458 16564 19462 16620
rect 19398 16560 19462 16564
rect 19478 16620 19542 16624
rect 19478 16564 19482 16620
rect 19482 16564 19538 16620
rect 19538 16564 19542 16620
rect 19478 16560 19542 16564
rect 19558 16620 19622 16624
rect 19558 16564 19562 16620
rect 19562 16564 19618 16620
rect 19618 16564 19622 16620
rect 19558 16560 19622 16564
rect 19638 16620 19702 16624
rect 19638 16564 19642 16620
rect 19642 16564 19698 16620
rect 19698 16564 19702 16620
rect 19638 16560 19702 16564
rect 19718 16620 19782 16624
rect 19718 16564 19722 16620
rect 19722 16564 19778 16620
rect 19778 16564 19782 16620
rect 19718 16560 19782 16564
rect 21266 16388 21330 16392
rect 21266 16332 21270 16388
rect 21270 16332 21326 16388
rect 21326 16332 21330 16388
rect 21266 16328 21330 16332
rect 9278 16076 9342 16080
rect 9278 16020 9282 16076
rect 9282 16020 9338 16076
rect 9338 16020 9342 16076
rect 9278 16016 9342 16020
rect 9358 16076 9422 16080
rect 9358 16020 9362 16076
rect 9362 16020 9418 16076
rect 9418 16020 9422 16076
rect 9358 16016 9422 16020
rect 9438 16076 9502 16080
rect 9438 16020 9442 16076
rect 9442 16020 9498 16076
rect 9498 16020 9502 16076
rect 9438 16016 9502 16020
rect 9518 16076 9582 16080
rect 9518 16020 9522 16076
rect 9522 16020 9578 16076
rect 9578 16020 9582 16076
rect 9518 16016 9582 16020
rect 9598 16076 9662 16080
rect 9598 16020 9602 16076
rect 9602 16020 9658 16076
rect 9658 16020 9662 16076
rect 9598 16016 9662 16020
rect 9678 16076 9742 16080
rect 9678 16020 9682 16076
rect 9682 16020 9738 16076
rect 9738 16020 9742 16076
rect 9678 16016 9742 16020
rect 9758 16076 9822 16080
rect 9758 16020 9762 16076
rect 9762 16020 9818 16076
rect 9818 16020 9822 16076
rect 9758 16016 9822 16020
rect 14878 16076 14942 16080
rect 14878 16020 14882 16076
rect 14882 16020 14938 16076
rect 14938 16020 14942 16076
rect 14878 16016 14942 16020
rect 14958 16076 15022 16080
rect 14958 16020 14962 16076
rect 14962 16020 15018 16076
rect 15018 16020 15022 16076
rect 14958 16016 15022 16020
rect 15038 16076 15102 16080
rect 15038 16020 15042 16076
rect 15042 16020 15098 16076
rect 15098 16020 15102 16076
rect 15038 16016 15102 16020
rect 15118 16076 15182 16080
rect 15118 16020 15122 16076
rect 15122 16020 15178 16076
rect 15178 16020 15182 16076
rect 15118 16016 15182 16020
rect 15198 16076 15262 16080
rect 15198 16020 15202 16076
rect 15202 16020 15258 16076
rect 15258 16020 15262 16076
rect 15198 16016 15262 16020
rect 15278 16076 15342 16080
rect 15278 16020 15282 16076
rect 15282 16020 15338 16076
rect 15338 16020 15342 16076
rect 15278 16016 15342 16020
rect 15358 16076 15422 16080
rect 15358 16020 15362 16076
rect 15362 16020 15418 16076
rect 15418 16020 15422 16076
rect 15358 16016 15422 16020
rect 20478 16076 20542 16080
rect 20478 16020 20482 16076
rect 20482 16020 20538 16076
rect 20538 16020 20542 16076
rect 20478 16016 20542 16020
rect 20558 16076 20622 16080
rect 20558 16020 20562 16076
rect 20562 16020 20618 16076
rect 20618 16020 20622 16076
rect 20558 16016 20622 16020
rect 20638 16076 20702 16080
rect 20638 16020 20642 16076
rect 20642 16020 20698 16076
rect 20698 16020 20702 16076
rect 20638 16016 20702 16020
rect 20718 16076 20782 16080
rect 20718 16020 20722 16076
rect 20722 16020 20778 16076
rect 20778 16020 20782 16076
rect 20718 16016 20782 16020
rect 20798 16076 20862 16080
rect 20798 16020 20802 16076
rect 20802 16020 20858 16076
rect 20858 16020 20862 16076
rect 20798 16016 20862 16020
rect 20878 16076 20942 16080
rect 20878 16020 20882 16076
rect 20882 16020 20938 16076
rect 20938 16020 20942 16076
rect 20878 16016 20942 16020
rect 20958 16076 21022 16080
rect 20958 16020 20962 16076
rect 20962 16020 21018 16076
rect 21018 16020 21022 16076
rect 20958 16016 21022 16020
rect 8038 15532 8102 15536
rect 8038 15476 8042 15532
rect 8042 15476 8098 15532
rect 8098 15476 8102 15532
rect 8038 15472 8102 15476
rect 8118 15532 8182 15536
rect 8118 15476 8122 15532
rect 8122 15476 8178 15532
rect 8178 15476 8182 15532
rect 8118 15472 8182 15476
rect 8198 15532 8262 15536
rect 8198 15476 8202 15532
rect 8202 15476 8258 15532
rect 8258 15476 8262 15532
rect 8198 15472 8262 15476
rect 8278 15532 8342 15536
rect 8278 15476 8282 15532
rect 8282 15476 8338 15532
rect 8338 15476 8342 15532
rect 8278 15472 8342 15476
rect 8358 15532 8422 15536
rect 8358 15476 8362 15532
rect 8362 15476 8418 15532
rect 8418 15476 8422 15532
rect 8358 15472 8422 15476
rect 8438 15532 8502 15536
rect 8438 15476 8442 15532
rect 8442 15476 8498 15532
rect 8498 15476 8502 15532
rect 8438 15472 8502 15476
rect 8518 15532 8582 15536
rect 8518 15476 8522 15532
rect 8522 15476 8578 15532
rect 8578 15476 8582 15532
rect 8518 15472 8582 15476
rect 13638 15532 13702 15536
rect 13638 15476 13642 15532
rect 13642 15476 13698 15532
rect 13698 15476 13702 15532
rect 13638 15472 13702 15476
rect 13718 15532 13782 15536
rect 13718 15476 13722 15532
rect 13722 15476 13778 15532
rect 13778 15476 13782 15532
rect 13718 15472 13782 15476
rect 13798 15532 13862 15536
rect 13798 15476 13802 15532
rect 13802 15476 13858 15532
rect 13858 15476 13862 15532
rect 13798 15472 13862 15476
rect 13878 15532 13942 15536
rect 13878 15476 13882 15532
rect 13882 15476 13938 15532
rect 13938 15476 13942 15532
rect 13878 15472 13942 15476
rect 13958 15532 14022 15536
rect 13958 15476 13962 15532
rect 13962 15476 14018 15532
rect 14018 15476 14022 15532
rect 13958 15472 14022 15476
rect 14038 15532 14102 15536
rect 14038 15476 14042 15532
rect 14042 15476 14098 15532
rect 14098 15476 14102 15532
rect 14038 15472 14102 15476
rect 14118 15532 14182 15536
rect 14118 15476 14122 15532
rect 14122 15476 14178 15532
rect 14178 15476 14182 15532
rect 14118 15472 14182 15476
rect 19238 15532 19302 15536
rect 19238 15476 19242 15532
rect 19242 15476 19298 15532
rect 19298 15476 19302 15532
rect 19238 15472 19302 15476
rect 19318 15532 19382 15536
rect 19318 15476 19322 15532
rect 19322 15476 19378 15532
rect 19378 15476 19382 15532
rect 19318 15472 19382 15476
rect 19398 15532 19462 15536
rect 19398 15476 19402 15532
rect 19402 15476 19458 15532
rect 19458 15476 19462 15532
rect 19398 15472 19462 15476
rect 19478 15532 19542 15536
rect 19478 15476 19482 15532
rect 19482 15476 19538 15532
rect 19538 15476 19542 15532
rect 19478 15472 19542 15476
rect 19558 15532 19622 15536
rect 19558 15476 19562 15532
rect 19562 15476 19618 15532
rect 19618 15476 19622 15532
rect 19558 15472 19622 15476
rect 19638 15532 19702 15536
rect 19638 15476 19642 15532
rect 19642 15476 19698 15532
rect 19698 15476 19702 15532
rect 19638 15472 19702 15476
rect 19718 15532 19782 15536
rect 19718 15476 19722 15532
rect 19722 15476 19778 15532
rect 19778 15476 19782 15532
rect 19718 15472 19782 15476
rect 9278 14988 9342 14992
rect 9278 14932 9282 14988
rect 9282 14932 9338 14988
rect 9338 14932 9342 14988
rect 9278 14928 9342 14932
rect 9358 14988 9422 14992
rect 9358 14932 9362 14988
rect 9362 14932 9418 14988
rect 9418 14932 9422 14988
rect 9358 14928 9422 14932
rect 9438 14988 9502 14992
rect 9438 14932 9442 14988
rect 9442 14932 9498 14988
rect 9498 14932 9502 14988
rect 9438 14928 9502 14932
rect 9518 14988 9582 14992
rect 9518 14932 9522 14988
rect 9522 14932 9578 14988
rect 9578 14932 9582 14988
rect 9518 14928 9582 14932
rect 9598 14988 9662 14992
rect 9598 14932 9602 14988
rect 9602 14932 9658 14988
rect 9658 14932 9662 14988
rect 9598 14928 9662 14932
rect 9678 14988 9742 14992
rect 9678 14932 9682 14988
rect 9682 14932 9738 14988
rect 9738 14932 9742 14988
rect 9678 14928 9742 14932
rect 9758 14988 9822 14992
rect 9758 14932 9762 14988
rect 9762 14932 9818 14988
rect 9818 14932 9822 14988
rect 9758 14928 9822 14932
rect 14878 14988 14942 14992
rect 14878 14932 14882 14988
rect 14882 14932 14938 14988
rect 14938 14932 14942 14988
rect 14878 14928 14942 14932
rect 14958 14988 15022 14992
rect 14958 14932 14962 14988
rect 14962 14932 15018 14988
rect 15018 14932 15022 14988
rect 14958 14928 15022 14932
rect 15038 14988 15102 14992
rect 15038 14932 15042 14988
rect 15042 14932 15098 14988
rect 15098 14932 15102 14988
rect 15038 14928 15102 14932
rect 15118 14988 15182 14992
rect 15118 14932 15122 14988
rect 15122 14932 15178 14988
rect 15178 14932 15182 14988
rect 15118 14928 15182 14932
rect 15198 14988 15262 14992
rect 15198 14932 15202 14988
rect 15202 14932 15258 14988
rect 15258 14932 15262 14988
rect 15198 14928 15262 14932
rect 15278 14988 15342 14992
rect 15278 14932 15282 14988
rect 15282 14932 15338 14988
rect 15338 14932 15342 14988
rect 15278 14928 15342 14932
rect 15358 14988 15422 14992
rect 15358 14932 15362 14988
rect 15362 14932 15418 14988
rect 15418 14932 15422 14988
rect 15358 14928 15422 14932
rect 20478 14988 20542 14992
rect 20478 14932 20482 14988
rect 20482 14932 20538 14988
rect 20538 14932 20542 14988
rect 20478 14928 20542 14932
rect 20558 14988 20622 14992
rect 20558 14932 20562 14988
rect 20562 14932 20618 14988
rect 20618 14932 20622 14988
rect 20558 14928 20622 14932
rect 20638 14988 20702 14992
rect 20638 14932 20642 14988
rect 20642 14932 20698 14988
rect 20698 14932 20702 14988
rect 20638 14928 20702 14932
rect 20718 14988 20782 14992
rect 20718 14932 20722 14988
rect 20722 14932 20778 14988
rect 20778 14932 20782 14988
rect 20718 14928 20782 14932
rect 20798 14988 20862 14992
rect 20798 14932 20802 14988
rect 20802 14932 20858 14988
rect 20858 14932 20862 14988
rect 20798 14928 20862 14932
rect 20878 14988 20942 14992
rect 20878 14932 20882 14988
rect 20882 14932 20938 14988
rect 20938 14932 20942 14988
rect 20878 14928 20942 14932
rect 20958 14988 21022 14992
rect 20958 14932 20962 14988
rect 20962 14932 21018 14988
rect 21018 14932 21022 14988
rect 20958 14928 21022 14932
rect 8038 14444 8102 14448
rect 8038 14388 8042 14444
rect 8042 14388 8098 14444
rect 8098 14388 8102 14444
rect 8038 14384 8102 14388
rect 8118 14444 8182 14448
rect 8118 14388 8122 14444
rect 8122 14388 8178 14444
rect 8178 14388 8182 14444
rect 8118 14384 8182 14388
rect 8198 14444 8262 14448
rect 8198 14388 8202 14444
rect 8202 14388 8258 14444
rect 8258 14388 8262 14444
rect 8198 14384 8262 14388
rect 8278 14444 8342 14448
rect 8278 14388 8282 14444
rect 8282 14388 8338 14444
rect 8338 14388 8342 14444
rect 8278 14384 8342 14388
rect 8358 14444 8422 14448
rect 8358 14388 8362 14444
rect 8362 14388 8418 14444
rect 8418 14388 8422 14444
rect 8358 14384 8422 14388
rect 8438 14444 8502 14448
rect 8438 14388 8442 14444
rect 8442 14388 8498 14444
rect 8498 14388 8502 14444
rect 8438 14384 8502 14388
rect 8518 14444 8582 14448
rect 8518 14388 8522 14444
rect 8522 14388 8578 14444
rect 8578 14388 8582 14444
rect 8518 14384 8582 14388
rect 13638 14444 13702 14448
rect 13638 14388 13642 14444
rect 13642 14388 13698 14444
rect 13698 14388 13702 14444
rect 13638 14384 13702 14388
rect 13718 14444 13782 14448
rect 13718 14388 13722 14444
rect 13722 14388 13778 14444
rect 13778 14388 13782 14444
rect 13718 14384 13782 14388
rect 13798 14444 13862 14448
rect 13798 14388 13802 14444
rect 13802 14388 13858 14444
rect 13858 14388 13862 14444
rect 13798 14384 13862 14388
rect 13878 14444 13942 14448
rect 13878 14388 13882 14444
rect 13882 14388 13938 14444
rect 13938 14388 13942 14444
rect 13878 14384 13942 14388
rect 13958 14444 14022 14448
rect 13958 14388 13962 14444
rect 13962 14388 14018 14444
rect 14018 14388 14022 14444
rect 13958 14384 14022 14388
rect 14038 14444 14102 14448
rect 14038 14388 14042 14444
rect 14042 14388 14098 14444
rect 14098 14388 14102 14444
rect 14038 14384 14102 14388
rect 14118 14444 14182 14448
rect 14118 14388 14122 14444
rect 14122 14388 14178 14444
rect 14178 14388 14182 14444
rect 14118 14384 14182 14388
rect 19238 14444 19302 14448
rect 19238 14388 19242 14444
rect 19242 14388 19298 14444
rect 19298 14388 19302 14444
rect 19238 14384 19302 14388
rect 19318 14444 19382 14448
rect 19318 14388 19322 14444
rect 19322 14388 19378 14444
rect 19378 14388 19382 14444
rect 19318 14384 19382 14388
rect 19398 14444 19462 14448
rect 19398 14388 19402 14444
rect 19402 14388 19458 14444
rect 19458 14388 19462 14444
rect 19398 14384 19462 14388
rect 19478 14444 19542 14448
rect 19478 14388 19482 14444
rect 19482 14388 19538 14444
rect 19538 14388 19542 14444
rect 19478 14384 19542 14388
rect 19558 14444 19622 14448
rect 19558 14388 19562 14444
rect 19562 14388 19618 14444
rect 19618 14388 19622 14444
rect 19558 14384 19622 14388
rect 19638 14444 19702 14448
rect 19638 14388 19642 14444
rect 19642 14388 19698 14444
rect 19698 14388 19702 14444
rect 19638 14384 19702 14388
rect 19718 14444 19782 14448
rect 19718 14388 19722 14444
rect 19722 14388 19778 14444
rect 19778 14388 19782 14444
rect 19718 14384 19782 14388
rect 9278 13900 9342 13904
rect 9278 13844 9282 13900
rect 9282 13844 9338 13900
rect 9338 13844 9342 13900
rect 9278 13840 9342 13844
rect 9358 13900 9422 13904
rect 9358 13844 9362 13900
rect 9362 13844 9418 13900
rect 9418 13844 9422 13900
rect 9358 13840 9422 13844
rect 9438 13900 9502 13904
rect 9438 13844 9442 13900
rect 9442 13844 9498 13900
rect 9498 13844 9502 13900
rect 9438 13840 9502 13844
rect 9518 13900 9582 13904
rect 9518 13844 9522 13900
rect 9522 13844 9578 13900
rect 9578 13844 9582 13900
rect 9518 13840 9582 13844
rect 9598 13900 9662 13904
rect 9598 13844 9602 13900
rect 9602 13844 9658 13900
rect 9658 13844 9662 13900
rect 9598 13840 9662 13844
rect 9678 13900 9742 13904
rect 9678 13844 9682 13900
rect 9682 13844 9738 13900
rect 9738 13844 9742 13900
rect 9678 13840 9742 13844
rect 9758 13900 9822 13904
rect 9758 13844 9762 13900
rect 9762 13844 9818 13900
rect 9818 13844 9822 13900
rect 9758 13840 9822 13844
rect 14878 13900 14942 13904
rect 14878 13844 14882 13900
rect 14882 13844 14938 13900
rect 14938 13844 14942 13900
rect 14878 13840 14942 13844
rect 14958 13900 15022 13904
rect 14958 13844 14962 13900
rect 14962 13844 15018 13900
rect 15018 13844 15022 13900
rect 14958 13840 15022 13844
rect 15038 13900 15102 13904
rect 15038 13844 15042 13900
rect 15042 13844 15098 13900
rect 15098 13844 15102 13900
rect 15038 13840 15102 13844
rect 15118 13900 15182 13904
rect 15118 13844 15122 13900
rect 15122 13844 15178 13900
rect 15178 13844 15182 13900
rect 15118 13840 15182 13844
rect 15198 13900 15262 13904
rect 15198 13844 15202 13900
rect 15202 13844 15258 13900
rect 15258 13844 15262 13900
rect 15198 13840 15262 13844
rect 15278 13900 15342 13904
rect 15278 13844 15282 13900
rect 15282 13844 15338 13900
rect 15338 13844 15342 13900
rect 15278 13840 15342 13844
rect 15358 13900 15422 13904
rect 15358 13844 15362 13900
rect 15362 13844 15418 13900
rect 15418 13844 15422 13900
rect 15358 13840 15422 13844
rect 20478 13900 20542 13904
rect 20478 13844 20482 13900
rect 20482 13844 20538 13900
rect 20538 13844 20542 13900
rect 20478 13840 20542 13844
rect 20558 13900 20622 13904
rect 20558 13844 20562 13900
rect 20562 13844 20618 13900
rect 20618 13844 20622 13900
rect 20558 13840 20622 13844
rect 20638 13900 20702 13904
rect 20638 13844 20642 13900
rect 20642 13844 20698 13900
rect 20698 13844 20702 13900
rect 20638 13840 20702 13844
rect 20718 13900 20782 13904
rect 20718 13844 20722 13900
rect 20722 13844 20778 13900
rect 20778 13844 20782 13900
rect 20718 13840 20782 13844
rect 20798 13900 20862 13904
rect 20798 13844 20802 13900
rect 20802 13844 20858 13900
rect 20858 13844 20862 13900
rect 20798 13840 20862 13844
rect 20878 13900 20942 13904
rect 20878 13844 20882 13900
rect 20882 13844 20938 13900
rect 20938 13844 20942 13900
rect 20878 13840 20942 13844
rect 20958 13900 21022 13904
rect 20958 13844 20962 13900
rect 20962 13844 21018 13900
rect 21018 13844 21022 13900
rect 20958 13840 21022 13844
rect 8038 13356 8102 13360
rect 8038 13300 8042 13356
rect 8042 13300 8098 13356
rect 8098 13300 8102 13356
rect 8038 13296 8102 13300
rect 8118 13356 8182 13360
rect 8118 13300 8122 13356
rect 8122 13300 8178 13356
rect 8178 13300 8182 13356
rect 8118 13296 8182 13300
rect 8198 13356 8262 13360
rect 8198 13300 8202 13356
rect 8202 13300 8258 13356
rect 8258 13300 8262 13356
rect 8198 13296 8262 13300
rect 8278 13356 8342 13360
rect 8278 13300 8282 13356
rect 8282 13300 8338 13356
rect 8338 13300 8342 13356
rect 8278 13296 8342 13300
rect 8358 13356 8422 13360
rect 8358 13300 8362 13356
rect 8362 13300 8418 13356
rect 8418 13300 8422 13356
rect 8358 13296 8422 13300
rect 8438 13356 8502 13360
rect 8438 13300 8442 13356
rect 8442 13300 8498 13356
rect 8498 13300 8502 13356
rect 8438 13296 8502 13300
rect 8518 13356 8582 13360
rect 8518 13300 8522 13356
rect 8522 13300 8578 13356
rect 8578 13300 8582 13356
rect 8518 13296 8582 13300
rect 13638 13356 13702 13360
rect 13638 13300 13642 13356
rect 13642 13300 13698 13356
rect 13698 13300 13702 13356
rect 13638 13296 13702 13300
rect 13718 13356 13782 13360
rect 13718 13300 13722 13356
rect 13722 13300 13778 13356
rect 13778 13300 13782 13356
rect 13718 13296 13782 13300
rect 13798 13356 13862 13360
rect 13798 13300 13802 13356
rect 13802 13300 13858 13356
rect 13858 13300 13862 13356
rect 13798 13296 13862 13300
rect 13878 13356 13942 13360
rect 13878 13300 13882 13356
rect 13882 13300 13938 13356
rect 13938 13300 13942 13356
rect 13878 13296 13942 13300
rect 13958 13356 14022 13360
rect 13958 13300 13962 13356
rect 13962 13300 14018 13356
rect 14018 13300 14022 13356
rect 13958 13296 14022 13300
rect 14038 13356 14102 13360
rect 14038 13300 14042 13356
rect 14042 13300 14098 13356
rect 14098 13300 14102 13356
rect 14038 13296 14102 13300
rect 14118 13356 14182 13360
rect 14118 13300 14122 13356
rect 14122 13300 14178 13356
rect 14178 13300 14182 13356
rect 14118 13296 14182 13300
rect 19238 13356 19302 13360
rect 19238 13300 19242 13356
rect 19242 13300 19298 13356
rect 19298 13300 19302 13356
rect 19238 13296 19302 13300
rect 19318 13356 19382 13360
rect 19318 13300 19322 13356
rect 19322 13300 19378 13356
rect 19378 13300 19382 13356
rect 19318 13296 19382 13300
rect 19398 13356 19462 13360
rect 19398 13300 19402 13356
rect 19402 13300 19458 13356
rect 19458 13300 19462 13356
rect 19398 13296 19462 13300
rect 19478 13356 19542 13360
rect 19478 13300 19482 13356
rect 19482 13300 19538 13356
rect 19538 13300 19542 13356
rect 19478 13296 19542 13300
rect 19558 13356 19622 13360
rect 19558 13300 19562 13356
rect 19562 13300 19618 13356
rect 19618 13300 19622 13356
rect 19558 13296 19622 13300
rect 19638 13356 19702 13360
rect 19638 13300 19642 13356
rect 19642 13300 19698 13356
rect 19698 13300 19702 13356
rect 19638 13296 19702 13300
rect 19718 13356 19782 13360
rect 19718 13300 19722 13356
rect 19722 13300 19778 13356
rect 19778 13300 19782 13356
rect 19718 13296 19782 13300
rect 9278 12812 9342 12816
rect 9278 12756 9282 12812
rect 9282 12756 9338 12812
rect 9338 12756 9342 12812
rect 9278 12752 9342 12756
rect 9358 12812 9422 12816
rect 9358 12756 9362 12812
rect 9362 12756 9418 12812
rect 9418 12756 9422 12812
rect 9358 12752 9422 12756
rect 9438 12812 9502 12816
rect 9438 12756 9442 12812
rect 9442 12756 9498 12812
rect 9498 12756 9502 12812
rect 9438 12752 9502 12756
rect 9518 12812 9582 12816
rect 9518 12756 9522 12812
rect 9522 12756 9578 12812
rect 9578 12756 9582 12812
rect 9518 12752 9582 12756
rect 9598 12812 9662 12816
rect 9598 12756 9602 12812
rect 9602 12756 9658 12812
rect 9658 12756 9662 12812
rect 9598 12752 9662 12756
rect 9678 12812 9742 12816
rect 9678 12756 9682 12812
rect 9682 12756 9738 12812
rect 9738 12756 9742 12812
rect 9678 12752 9742 12756
rect 9758 12812 9822 12816
rect 9758 12756 9762 12812
rect 9762 12756 9818 12812
rect 9818 12756 9822 12812
rect 9758 12752 9822 12756
rect 14878 12812 14942 12816
rect 14878 12756 14882 12812
rect 14882 12756 14938 12812
rect 14938 12756 14942 12812
rect 14878 12752 14942 12756
rect 14958 12812 15022 12816
rect 14958 12756 14962 12812
rect 14962 12756 15018 12812
rect 15018 12756 15022 12812
rect 14958 12752 15022 12756
rect 15038 12812 15102 12816
rect 15038 12756 15042 12812
rect 15042 12756 15098 12812
rect 15098 12756 15102 12812
rect 15038 12752 15102 12756
rect 15118 12812 15182 12816
rect 15118 12756 15122 12812
rect 15122 12756 15178 12812
rect 15178 12756 15182 12812
rect 15118 12752 15182 12756
rect 15198 12812 15262 12816
rect 15198 12756 15202 12812
rect 15202 12756 15258 12812
rect 15258 12756 15262 12812
rect 15198 12752 15262 12756
rect 15278 12812 15342 12816
rect 15278 12756 15282 12812
rect 15282 12756 15338 12812
rect 15338 12756 15342 12812
rect 15278 12752 15342 12756
rect 15358 12812 15422 12816
rect 15358 12756 15362 12812
rect 15362 12756 15418 12812
rect 15418 12756 15422 12812
rect 15358 12752 15422 12756
rect 20478 12812 20542 12816
rect 20478 12756 20482 12812
rect 20482 12756 20538 12812
rect 20538 12756 20542 12812
rect 20478 12752 20542 12756
rect 20558 12812 20622 12816
rect 20558 12756 20562 12812
rect 20562 12756 20618 12812
rect 20618 12756 20622 12812
rect 20558 12752 20622 12756
rect 20638 12812 20702 12816
rect 20638 12756 20642 12812
rect 20642 12756 20698 12812
rect 20698 12756 20702 12812
rect 20638 12752 20702 12756
rect 20718 12812 20782 12816
rect 20718 12756 20722 12812
rect 20722 12756 20778 12812
rect 20778 12756 20782 12812
rect 20718 12752 20782 12756
rect 20798 12812 20862 12816
rect 20798 12756 20802 12812
rect 20802 12756 20858 12812
rect 20858 12756 20862 12812
rect 20798 12752 20862 12756
rect 20878 12812 20942 12816
rect 20878 12756 20882 12812
rect 20882 12756 20938 12812
rect 20938 12756 20942 12812
rect 20878 12752 20942 12756
rect 20958 12812 21022 12816
rect 20958 12756 20962 12812
rect 20962 12756 21018 12812
rect 21018 12756 21022 12812
rect 20958 12752 21022 12756
rect 8038 12268 8102 12272
rect 8038 12212 8042 12268
rect 8042 12212 8098 12268
rect 8098 12212 8102 12268
rect 8038 12208 8102 12212
rect 8118 12268 8182 12272
rect 8118 12212 8122 12268
rect 8122 12212 8178 12268
rect 8178 12212 8182 12268
rect 8118 12208 8182 12212
rect 8198 12268 8262 12272
rect 8198 12212 8202 12268
rect 8202 12212 8258 12268
rect 8258 12212 8262 12268
rect 8198 12208 8262 12212
rect 8278 12268 8342 12272
rect 8278 12212 8282 12268
rect 8282 12212 8338 12268
rect 8338 12212 8342 12268
rect 8278 12208 8342 12212
rect 8358 12268 8422 12272
rect 8358 12212 8362 12268
rect 8362 12212 8418 12268
rect 8418 12212 8422 12268
rect 8358 12208 8422 12212
rect 8438 12268 8502 12272
rect 8438 12212 8442 12268
rect 8442 12212 8498 12268
rect 8498 12212 8502 12268
rect 8438 12208 8502 12212
rect 8518 12268 8582 12272
rect 8518 12212 8522 12268
rect 8522 12212 8578 12268
rect 8578 12212 8582 12268
rect 8518 12208 8582 12212
rect 13638 12268 13702 12272
rect 13638 12212 13642 12268
rect 13642 12212 13698 12268
rect 13698 12212 13702 12268
rect 13638 12208 13702 12212
rect 13718 12268 13782 12272
rect 13718 12212 13722 12268
rect 13722 12212 13778 12268
rect 13778 12212 13782 12268
rect 13718 12208 13782 12212
rect 13798 12268 13862 12272
rect 13798 12212 13802 12268
rect 13802 12212 13858 12268
rect 13858 12212 13862 12268
rect 13798 12208 13862 12212
rect 13878 12268 13942 12272
rect 13878 12212 13882 12268
rect 13882 12212 13938 12268
rect 13938 12212 13942 12268
rect 13878 12208 13942 12212
rect 13958 12268 14022 12272
rect 13958 12212 13962 12268
rect 13962 12212 14018 12268
rect 14018 12212 14022 12268
rect 13958 12208 14022 12212
rect 14038 12268 14102 12272
rect 14038 12212 14042 12268
rect 14042 12212 14098 12268
rect 14098 12212 14102 12268
rect 14038 12208 14102 12212
rect 14118 12268 14182 12272
rect 14118 12212 14122 12268
rect 14122 12212 14178 12268
rect 14178 12212 14182 12268
rect 14118 12208 14182 12212
rect 19238 12268 19302 12272
rect 19238 12212 19242 12268
rect 19242 12212 19298 12268
rect 19298 12212 19302 12268
rect 19238 12208 19302 12212
rect 19318 12268 19382 12272
rect 19318 12212 19322 12268
rect 19322 12212 19378 12268
rect 19378 12212 19382 12268
rect 19318 12208 19382 12212
rect 19398 12268 19462 12272
rect 19398 12212 19402 12268
rect 19402 12212 19458 12268
rect 19458 12212 19462 12268
rect 19398 12208 19462 12212
rect 19478 12268 19542 12272
rect 19478 12212 19482 12268
rect 19482 12212 19538 12268
rect 19538 12212 19542 12268
rect 19478 12208 19542 12212
rect 19558 12268 19622 12272
rect 19558 12212 19562 12268
rect 19562 12212 19618 12268
rect 19618 12212 19622 12268
rect 19558 12208 19622 12212
rect 19638 12268 19702 12272
rect 19638 12212 19642 12268
rect 19642 12212 19698 12268
rect 19698 12212 19702 12268
rect 19638 12208 19702 12212
rect 19718 12268 19782 12272
rect 19718 12212 19722 12268
rect 19722 12212 19778 12268
rect 19778 12212 19782 12268
rect 19718 12208 19782 12212
rect 21266 11936 21330 12000
rect 9278 11724 9342 11728
rect 9278 11668 9282 11724
rect 9282 11668 9338 11724
rect 9338 11668 9342 11724
rect 9278 11664 9342 11668
rect 9358 11724 9422 11728
rect 9358 11668 9362 11724
rect 9362 11668 9418 11724
rect 9418 11668 9422 11724
rect 9358 11664 9422 11668
rect 9438 11724 9502 11728
rect 9438 11668 9442 11724
rect 9442 11668 9498 11724
rect 9498 11668 9502 11724
rect 9438 11664 9502 11668
rect 9518 11724 9582 11728
rect 9518 11668 9522 11724
rect 9522 11668 9578 11724
rect 9578 11668 9582 11724
rect 9518 11664 9582 11668
rect 9598 11724 9662 11728
rect 9598 11668 9602 11724
rect 9602 11668 9658 11724
rect 9658 11668 9662 11724
rect 9598 11664 9662 11668
rect 9678 11724 9742 11728
rect 9678 11668 9682 11724
rect 9682 11668 9738 11724
rect 9738 11668 9742 11724
rect 9678 11664 9742 11668
rect 9758 11724 9822 11728
rect 9758 11668 9762 11724
rect 9762 11668 9818 11724
rect 9818 11668 9822 11724
rect 9758 11664 9822 11668
rect 14878 11724 14942 11728
rect 14878 11668 14882 11724
rect 14882 11668 14938 11724
rect 14938 11668 14942 11724
rect 14878 11664 14942 11668
rect 14958 11724 15022 11728
rect 14958 11668 14962 11724
rect 14962 11668 15018 11724
rect 15018 11668 15022 11724
rect 14958 11664 15022 11668
rect 15038 11724 15102 11728
rect 15038 11668 15042 11724
rect 15042 11668 15098 11724
rect 15098 11668 15102 11724
rect 15038 11664 15102 11668
rect 15118 11724 15182 11728
rect 15118 11668 15122 11724
rect 15122 11668 15178 11724
rect 15178 11668 15182 11724
rect 15118 11664 15182 11668
rect 15198 11724 15262 11728
rect 15198 11668 15202 11724
rect 15202 11668 15258 11724
rect 15258 11668 15262 11724
rect 15198 11664 15262 11668
rect 15278 11724 15342 11728
rect 15278 11668 15282 11724
rect 15282 11668 15338 11724
rect 15338 11668 15342 11724
rect 15278 11664 15342 11668
rect 15358 11724 15422 11728
rect 15358 11668 15362 11724
rect 15362 11668 15418 11724
rect 15418 11668 15422 11724
rect 15358 11664 15422 11668
rect 20478 11724 20542 11728
rect 20478 11668 20482 11724
rect 20482 11668 20538 11724
rect 20538 11668 20542 11724
rect 20478 11664 20542 11668
rect 20558 11724 20622 11728
rect 20558 11668 20562 11724
rect 20562 11668 20618 11724
rect 20618 11668 20622 11724
rect 20558 11664 20622 11668
rect 20638 11724 20702 11728
rect 20638 11668 20642 11724
rect 20642 11668 20698 11724
rect 20698 11668 20702 11724
rect 20638 11664 20702 11668
rect 20718 11724 20782 11728
rect 20718 11668 20722 11724
rect 20722 11668 20778 11724
rect 20778 11668 20782 11724
rect 20718 11664 20782 11668
rect 20798 11724 20862 11728
rect 20798 11668 20802 11724
rect 20802 11668 20858 11724
rect 20858 11668 20862 11724
rect 20798 11664 20862 11668
rect 20878 11724 20942 11728
rect 20878 11668 20882 11724
rect 20882 11668 20938 11724
rect 20938 11668 20942 11724
rect 20878 11664 20942 11668
rect 20958 11724 21022 11728
rect 20958 11668 20962 11724
rect 20962 11668 21018 11724
rect 21018 11668 21022 11724
rect 20958 11664 21022 11668
rect 8038 11180 8102 11184
rect 8038 11124 8042 11180
rect 8042 11124 8098 11180
rect 8098 11124 8102 11180
rect 8038 11120 8102 11124
rect 8118 11180 8182 11184
rect 8118 11124 8122 11180
rect 8122 11124 8178 11180
rect 8178 11124 8182 11180
rect 8118 11120 8182 11124
rect 8198 11180 8262 11184
rect 8198 11124 8202 11180
rect 8202 11124 8258 11180
rect 8258 11124 8262 11180
rect 8198 11120 8262 11124
rect 8278 11180 8342 11184
rect 8278 11124 8282 11180
rect 8282 11124 8338 11180
rect 8338 11124 8342 11180
rect 8278 11120 8342 11124
rect 8358 11180 8422 11184
rect 8358 11124 8362 11180
rect 8362 11124 8418 11180
rect 8418 11124 8422 11180
rect 8358 11120 8422 11124
rect 8438 11180 8502 11184
rect 8438 11124 8442 11180
rect 8442 11124 8498 11180
rect 8498 11124 8502 11180
rect 8438 11120 8502 11124
rect 8518 11180 8582 11184
rect 8518 11124 8522 11180
rect 8522 11124 8578 11180
rect 8578 11124 8582 11180
rect 8518 11120 8582 11124
rect 13638 11180 13702 11184
rect 13638 11124 13642 11180
rect 13642 11124 13698 11180
rect 13698 11124 13702 11180
rect 13638 11120 13702 11124
rect 13718 11180 13782 11184
rect 13718 11124 13722 11180
rect 13722 11124 13778 11180
rect 13778 11124 13782 11180
rect 13718 11120 13782 11124
rect 13798 11180 13862 11184
rect 13798 11124 13802 11180
rect 13802 11124 13858 11180
rect 13858 11124 13862 11180
rect 13798 11120 13862 11124
rect 13878 11180 13942 11184
rect 13878 11124 13882 11180
rect 13882 11124 13938 11180
rect 13938 11124 13942 11180
rect 13878 11120 13942 11124
rect 13958 11180 14022 11184
rect 13958 11124 13962 11180
rect 13962 11124 14018 11180
rect 14018 11124 14022 11180
rect 13958 11120 14022 11124
rect 14038 11180 14102 11184
rect 14038 11124 14042 11180
rect 14042 11124 14098 11180
rect 14098 11124 14102 11180
rect 14038 11120 14102 11124
rect 14118 11180 14182 11184
rect 14118 11124 14122 11180
rect 14122 11124 14178 11180
rect 14178 11124 14182 11180
rect 14118 11120 14182 11124
rect 19238 11180 19302 11184
rect 19238 11124 19242 11180
rect 19242 11124 19298 11180
rect 19298 11124 19302 11180
rect 19238 11120 19302 11124
rect 19318 11180 19382 11184
rect 19318 11124 19322 11180
rect 19322 11124 19378 11180
rect 19378 11124 19382 11180
rect 19318 11120 19382 11124
rect 19398 11180 19462 11184
rect 19398 11124 19402 11180
rect 19402 11124 19458 11180
rect 19458 11124 19462 11180
rect 19398 11120 19462 11124
rect 19478 11180 19542 11184
rect 19478 11124 19482 11180
rect 19482 11124 19538 11180
rect 19538 11124 19542 11180
rect 19478 11120 19542 11124
rect 19558 11180 19622 11184
rect 19558 11124 19562 11180
rect 19562 11124 19618 11180
rect 19618 11124 19622 11180
rect 19558 11120 19622 11124
rect 19638 11180 19702 11184
rect 19638 11124 19642 11180
rect 19642 11124 19698 11180
rect 19698 11124 19702 11180
rect 19638 11120 19702 11124
rect 19718 11180 19782 11184
rect 19718 11124 19722 11180
rect 19722 11124 19778 11180
rect 19778 11124 19782 11180
rect 19718 11120 19782 11124
rect 9278 10636 9342 10640
rect 9278 10580 9282 10636
rect 9282 10580 9338 10636
rect 9338 10580 9342 10636
rect 9278 10576 9342 10580
rect 9358 10636 9422 10640
rect 9358 10580 9362 10636
rect 9362 10580 9418 10636
rect 9418 10580 9422 10636
rect 9358 10576 9422 10580
rect 9438 10636 9502 10640
rect 9438 10580 9442 10636
rect 9442 10580 9498 10636
rect 9498 10580 9502 10636
rect 9438 10576 9502 10580
rect 9518 10636 9582 10640
rect 9518 10580 9522 10636
rect 9522 10580 9578 10636
rect 9578 10580 9582 10636
rect 9518 10576 9582 10580
rect 9598 10636 9662 10640
rect 9598 10580 9602 10636
rect 9602 10580 9658 10636
rect 9658 10580 9662 10636
rect 9598 10576 9662 10580
rect 9678 10636 9742 10640
rect 9678 10580 9682 10636
rect 9682 10580 9738 10636
rect 9738 10580 9742 10636
rect 9678 10576 9742 10580
rect 9758 10636 9822 10640
rect 9758 10580 9762 10636
rect 9762 10580 9818 10636
rect 9818 10580 9822 10636
rect 9758 10576 9822 10580
rect 14878 10636 14942 10640
rect 14878 10580 14882 10636
rect 14882 10580 14938 10636
rect 14938 10580 14942 10636
rect 14878 10576 14942 10580
rect 14958 10636 15022 10640
rect 14958 10580 14962 10636
rect 14962 10580 15018 10636
rect 15018 10580 15022 10636
rect 14958 10576 15022 10580
rect 15038 10636 15102 10640
rect 15038 10580 15042 10636
rect 15042 10580 15098 10636
rect 15098 10580 15102 10636
rect 15038 10576 15102 10580
rect 15118 10636 15182 10640
rect 15118 10580 15122 10636
rect 15122 10580 15178 10636
rect 15178 10580 15182 10636
rect 15118 10576 15182 10580
rect 15198 10636 15262 10640
rect 15198 10580 15202 10636
rect 15202 10580 15258 10636
rect 15258 10580 15262 10636
rect 15198 10576 15262 10580
rect 15278 10636 15342 10640
rect 15278 10580 15282 10636
rect 15282 10580 15338 10636
rect 15338 10580 15342 10636
rect 15278 10576 15342 10580
rect 15358 10636 15422 10640
rect 15358 10580 15362 10636
rect 15362 10580 15418 10636
rect 15418 10580 15422 10636
rect 15358 10576 15422 10580
rect 20478 10636 20542 10640
rect 20478 10580 20482 10636
rect 20482 10580 20538 10636
rect 20538 10580 20542 10636
rect 20478 10576 20542 10580
rect 20558 10636 20622 10640
rect 20558 10580 20562 10636
rect 20562 10580 20618 10636
rect 20618 10580 20622 10636
rect 20558 10576 20622 10580
rect 20638 10636 20702 10640
rect 20638 10580 20642 10636
rect 20642 10580 20698 10636
rect 20698 10580 20702 10636
rect 20638 10576 20702 10580
rect 20718 10636 20782 10640
rect 20718 10580 20722 10636
rect 20722 10580 20778 10636
rect 20778 10580 20782 10636
rect 20718 10576 20782 10580
rect 20798 10636 20862 10640
rect 20798 10580 20802 10636
rect 20802 10580 20858 10636
rect 20858 10580 20862 10636
rect 20798 10576 20862 10580
rect 20878 10636 20942 10640
rect 20878 10580 20882 10636
rect 20882 10580 20938 10636
rect 20938 10580 20942 10636
rect 20878 10576 20942 10580
rect 20958 10636 21022 10640
rect 20958 10580 20962 10636
rect 20962 10580 21018 10636
rect 21018 10580 21022 10636
rect 20958 10576 21022 10580
rect 8038 10092 8102 10096
rect 8038 10036 8042 10092
rect 8042 10036 8098 10092
rect 8098 10036 8102 10092
rect 8038 10032 8102 10036
rect 8118 10092 8182 10096
rect 8118 10036 8122 10092
rect 8122 10036 8178 10092
rect 8178 10036 8182 10092
rect 8118 10032 8182 10036
rect 8198 10092 8262 10096
rect 8198 10036 8202 10092
rect 8202 10036 8258 10092
rect 8258 10036 8262 10092
rect 8198 10032 8262 10036
rect 8278 10092 8342 10096
rect 8278 10036 8282 10092
rect 8282 10036 8338 10092
rect 8338 10036 8342 10092
rect 8278 10032 8342 10036
rect 8358 10092 8422 10096
rect 8358 10036 8362 10092
rect 8362 10036 8418 10092
rect 8418 10036 8422 10092
rect 8358 10032 8422 10036
rect 8438 10092 8502 10096
rect 8438 10036 8442 10092
rect 8442 10036 8498 10092
rect 8498 10036 8502 10092
rect 8438 10032 8502 10036
rect 8518 10092 8582 10096
rect 8518 10036 8522 10092
rect 8522 10036 8578 10092
rect 8578 10036 8582 10092
rect 8518 10032 8582 10036
rect 13638 10092 13702 10096
rect 13638 10036 13642 10092
rect 13642 10036 13698 10092
rect 13698 10036 13702 10092
rect 13638 10032 13702 10036
rect 13718 10092 13782 10096
rect 13718 10036 13722 10092
rect 13722 10036 13778 10092
rect 13778 10036 13782 10092
rect 13718 10032 13782 10036
rect 13798 10092 13862 10096
rect 13798 10036 13802 10092
rect 13802 10036 13858 10092
rect 13858 10036 13862 10092
rect 13798 10032 13862 10036
rect 13878 10092 13942 10096
rect 13878 10036 13882 10092
rect 13882 10036 13938 10092
rect 13938 10036 13942 10092
rect 13878 10032 13942 10036
rect 13958 10092 14022 10096
rect 13958 10036 13962 10092
rect 13962 10036 14018 10092
rect 14018 10036 14022 10092
rect 13958 10032 14022 10036
rect 14038 10092 14102 10096
rect 14038 10036 14042 10092
rect 14042 10036 14098 10092
rect 14098 10036 14102 10092
rect 14038 10032 14102 10036
rect 14118 10092 14182 10096
rect 14118 10036 14122 10092
rect 14122 10036 14178 10092
rect 14178 10036 14182 10092
rect 14118 10032 14182 10036
rect 19238 10092 19302 10096
rect 19238 10036 19242 10092
rect 19242 10036 19298 10092
rect 19298 10036 19302 10092
rect 19238 10032 19302 10036
rect 19318 10092 19382 10096
rect 19318 10036 19322 10092
rect 19322 10036 19378 10092
rect 19378 10036 19382 10092
rect 19318 10032 19382 10036
rect 19398 10092 19462 10096
rect 19398 10036 19402 10092
rect 19402 10036 19458 10092
rect 19458 10036 19462 10092
rect 19398 10032 19462 10036
rect 19478 10092 19542 10096
rect 19478 10036 19482 10092
rect 19482 10036 19538 10092
rect 19538 10036 19542 10092
rect 19478 10032 19542 10036
rect 19558 10092 19622 10096
rect 19558 10036 19562 10092
rect 19562 10036 19618 10092
rect 19618 10036 19622 10092
rect 19558 10032 19622 10036
rect 19638 10092 19702 10096
rect 19638 10036 19642 10092
rect 19642 10036 19698 10092
rect 19698 10036 19702 10092
rect 19638 10032 19702 10036
rect 19718 10092 19782 10096
rect 19718 10036 19722 10092
rect 19722 10036 19778 10092
rect 19778 10036 19782 10092
rect 19718 10032 19782 10036
rect 9278 9548 9342 9552
rect 9278 9492 9282 9548
rect 9282 9492 9338 9548
rect 9338 9492 9342 9548
rect 9278 9488 9342 9492
rect 9358 9548 9422 9552
rect 9358 9492 9362 9548
rect 9362 9492 9418 9548
rect 9418 9492 9422 9548
rect 9358 9488 9422 9492
rect 9438 9548 9502 9552
rect 9438 9492 9442 9548
rect 9442 9492 9498 9548
rect 9498 9492 9502 9548
rect 9438 9488 9502 9492
rect 9518 9548 9582 9552
rect 9518 9492 9522 9548
rect 9522 9492 9578 9548
rect 9578 9492 9582 9548
rect 9518 9488 9582 9492
rect 9598 9548 9662 9552
rect 9598 9492 9602 9548
rect 9602 9492 9658 9548
rect 9658 9492 9662 9548
rect 9598 9488 9662 9492
rect 9678 9548 9742 9552
rect 9678 9492 9682 9548
rect 9682 9492 9738 9548
rect 9738 9492 9742 9548
rect 9678 9488 9742 9492
rect 9758 9548 9822 9552
rect 9758 9492 9762 9548
rect 9762 9492 9818 9548
rect 9818 9492 9822 9548
rect 9758 9488 9822 9492
rect 14878 9548 14942 9552
rect 14878 9492 14882 9548
rect 14882 9492 14938 9548
rect 14938 9492 14942 9548
rect 14878 9488 14942 9492
rect 14958 9548 15022 9552
rect 14958 9492 14962 9548
rect 14962 9492 15018 9548
rect 15018 9492 15022 9548
rect 14958 9488 15022 9492
rect 15038 9548 15102 9552
rect 15038 9492 15042 9548
rect 15042 9492 15098 9548
rect 15098 9492 15102 9548
rect 15038 9488 15102 9492
rect 15118 9548 15182 9552
rect 15118 9492 15122 9548
rect 15122 9492 15178 9548
rect 15178 9492 15182 9548
rect 15118 9488 15182 9492
rect 15198 9548 15262 9552
rect 15198 9492 15202 9548
rect 15202 9492 15258 9548
rect 15258 9492 15262 9548
rect 15198 9488 15262 9492
rect 15278 9548 15342 9552
rect 15278 9492 15282 9548
rect 15282 9492 15338 9548
rect 15338 9492 15342 9548
rect 15278 9488 15342 9492
rect 15358 9548 15422 9552
rect 15358 9492 15362 9548
rect 15362 9492 15418 9548
rect 15418 9492 15422 9548
rect 15358 9488 15422 9492
rect 17126 9496 17190 9560
rect 20478 9548 20542 9552
rect 20478 9492 20482 9548
rect 20482 9492 20538 9548
rect 20538 9492 20542 9548
rect 20478 9488 20542 9492
rect 20558 9548 20622 9552
rect 20558 9492 20562 9548
rect 20562 9492 20618 9548
rect 20618 9492 20622 9548
rect 20558 9488 20622 9492
rect 20638 9548 20702 9552
rect 20638 9492 20642 9548
rect 20642 9492 20698 9548
rect 20698 9492 20702 9548
rect 20638 9488 20702 9492
rect 20718 9548 20782 9552
rect 20718 9492 20722 9548
rect 20722 9492 20778 9548
rect 20778 9492 20782 9548
rect 20718 9488 20782 9492
rect 20798 9548 20862 9552
rect 20798 9492 20802 9548
rect 20802 9492 20858 9548
rect 20858 9492 20862 9548
rect 20798 9488 20862 9492
rect 20878 9548 20942 9552
rect 20878 9492 20882 9548
rect 20882 9492 20938 9548
rect 20938 9492 20942 9548
rect 20878 9488 20942 9492
rect 20958 9548 21022 9552
rect 20958 9492 20962 9548
rect 20962 9492 21018 9548
rect 21018 9492 21022 9548
rect 20958 9488 21022 9492
rect 8038 9004 8102 9008
rect 8038 8948 8042 9004
rect 8042 8948 8098 9004
rect 8098 8948 8102 9004
rect 8038 8944 8102 8948
rect 8118 9004 8182 9008
rect 8118 8948 8122 9004
rect 8122 8948 8178 9004
rect 8178 8948 8182 9004
rect 8118 8944 8182 8948
rect 8198 9004 8262 9008
rect 8198 8948 8202 9004
rect 8202 8948 8258 9004
rect 8258 8948 8262 9004
rect 8198 8944 8262 8948
rect 8278 9004 8342 9008
rect 8278 8948 8282 9004
rect 8282 8948 8338 9004
rect 8338 8948 8342 9004
rect 8278 8944 8342 8948
rect 8358 9004 8422 9008
rect 8358 8948 8362 9004
rect 8362 8948 8418 9004
rect 8418 8948 8422 9004
rect 8358 8944 8422 8948
rect 8438 9004 8502 9008
rect 8438 8948 8442 9004
rect 8442 8948 8498 9004
rect 8498 8948 8502 9004
rect 8438 8944 8502 8948
rect 8518 9004 8582 9008
rect 8518 8948 8522 9004
rect 8522 8948 8578 9004
rect 8578 8948 8582 9004
rect 8518 8944 8582 8948
rect 13638 9004 13702 9008
rect 13638 8948 13642 9004
rect 13642 8948 13698 9004
rect 13698 8948 13702 9004
rect 13638 8944 13702 8948
rect 13718 9004 13782 9008
rect 13718 8948 13722 9004
rect 13722 8948 13778 9004
rect 13778 8948 13782 9004
rect 13718 8944 13782 8948
rect 13798 9004 13862 9008
rect 13798 8948 13802 9004
rect 13802 8948 13858 9004
rect 13858 8948 13862 9004
rect 13798 8944 13862 8948
rect 13878 9004 13942 9008
rect 13878 8948 13882 9004
rect 13882 8948 13938 9004
rect 13938 8948 13942 9004
rect 13878 8944 13942 8948
rect 13958 9004 14022 9008
rect 13958 8948 13962 9004
rect 13962 8948 14018 9004
rect 14018 8948 14022 9004
rect 13958 8944 14022 8948
rect 14038 9004 14102 9008
rect 14038 8948 14042 9004
rect 14042 8948 14098 9004
rect 14098 8948 14102 9004
rect 14038 8944 14102 8948
rect 14118 9004 14182 9008
rect 14118 8948 14122 9004
rect 14122 8948 14178 9004
rect 14178 8948 14182 9004
rect 14118 8944 14182 8948
rect 19238 9004 19302 9008
rect 19238 8948 19242 9004
rect 19242 8948 19298 9004
rect 19298 8948 19302 9004
rect 19238 8944 19302 8948
rect 19318 9004 19382 9008
rect 19318 8948 19322 9004
rect 19322 8948 19378 9004
rect 19378 8948 19382 9004
rect 19318 8944 19382 8948
rect 19398 9004 19462 9008
rect 19398 8948 19402 9004
rect 19402 8948 19458 9004
rect 19458 8948 19462 9004
rect 19398 8944 19462 8948
rect 19478 9004 19542 9008
rect 19478 8948 19482 9004
rect 19482 8948 19538 9004
rect 19538 8948 19542 9004
rect 19478 8944 19542 8948
rect 19558 9004 19622 9008
rect 19558 8948 19562 9004
rect 19562 8948 19618 9004
rect 19618 8948 19622 9004
rect 19558 8944 19622 8948
rect 19638 9004 19702 9008
rect 19638 8948 19642 9004
rect 19642 8948 19698 9004
rect 19698 8948 19702 9004
rect 19638 8944 19702 8948
rect 19718 9004 19782 9008
rect 19718 8948 19722 9004
rect 19722 8948 19778 9004
rect 19778 8948 19782 9004
rect 19718 8944 19782 8948
rect 9278 8460 9342 8464
rect 9278 8404 9282 8460
rect 9282 8404 9338 8460
rect 9338 8404 9342 8460
rect 9278 8400 9342 8404
rect 9358 8460 9422 8464
rect 9358 8404 9362 8460
rect 9362 8404 9418 8460
rect 9418 8404 9422 8460
rect 9358 8400 9422 8404
rect 9438 8460 9502 8464
rect 9438 8404 9442 8460
rect 9442 8404 9498 8460
rect 9498 8404 9502 8460
rect 9438 8400 9502 8404
rect 9518 8460 9582 8464
rect 9518 8404 9522 8460
rect 9522 8404 9578 8460
rect 9578 8404 9582 8460
rect 9518 8400 9582 8404
rect 9598 8460 9662 8464
rect 9598 8404 9602 8460
rect 9602 8404 9658 8460
rect 9658 8404 9662 8460
rect 9598 8400 9662 8404
rect 9678 8460 9742 8464
rect 9678 8404 9682 8460
rect 9682 8404 9738 8460
rect 9738 8404 9742 8460
rect 9678 8400 9742 8404
rect 9758 8460 9822 8464
rect 9758 8404 9762 8460
rect 9762 8404 9818 8460
rect 9818 8404 9822 8460
rect 9758 8400 9822 8404
rect 14878 8460 14942 8464
rect 14878 8404 14882 8460
rect 14882 8404 14938 8460
rect 14938 8404 14942 8460
rect 14878 8400 14942 8404
rect 14958 8460 15022 8464
rect 14958 8404 14962 8460
rect 14962 8404 15018 8460
rect 15018 8404 15022 8460
rect 14958 8400 15022 8404
rect 15038 8460 15102 8464
rect 15038 8404 15042 8460
rect 15042 8404 15098 8460
rect 15098 8404 15102 8460
rect 15038 8400 15102 8404
rect 15118 8460 15182 8464
rect 15118 8404 15122 8460
rect 15122 8404 15178 8460
rect 15178 8404 15182 8460
rect 15118 8400 15182 8404
rect 15198 8460 15262 8464
rect 15198 8404 15202 8460
rect 15202 8404 15258 8460
rect 15258 8404 15262 8460
rect 15198 8400 15262 8404
rect 15278 8460 15342 8464
rect 15278 8404 15282 8460
rect 15282 8404 15338 8460
rect 15338 8404 15342 8460
rect 15278 8400 15342 8404
rect 15358 8460 15422 8464
rect 15358 8404 15362 8460
rect 15362 8404 15418 8460
rect 15418 8404 15422 8460
rect 15358 8400 15422 8404
rect 20478 8460 20542 8464
rect 20478 8404 20482 8460
rect 20482 8404 20538 8460
rect 20538 8404 20542 8460
rect 20478 8400 20542 8404
rect 20558 8460 20622 8464
rect 20558 8404 20562 8460
rect 20562 8404 20618 8460
rect 20618 8404 20622 8460
rect 20558 8400 20622 8404
rect 20638 8460 20702 8464
rect 20638 8404 20642 8460
rect 20642 8404 20698 8460
rect 20698 8404 20702 8460
rect 20638 8400 20702 8404
rect 20718 8460 20782 8464
rect 20718 8404 20722 8460
rect 20722 8404 20778 8460
rect 20778 8404 20782 8460
rect 20718 8400 20782 8404
rect 20798 8460 20862 8464
rect 20798 8404 20802 8460
rect 20802 8404 20858 8460
rect 20858 8404 20862 8460
rect 20798 8400 20862 8404
rect 20878 8460 20942 8464
rect 20878 8404 20882 8460
rect 20882 8404 20938 8460
rect 20938 8404 20942 8460
rect 20878 8400 20942 8404
rect 20958 8460 21022 8464
rect 20958 8404 20962 8460
rect 20962 8404 21018 8460
rect 21018 8404 21022 8460
rect 20958 8400 21022 8404
rect 21266 8336 21330 8340
rect 21266 8280 21270 8336
rect 21270 8280 21326 8336
rect 21326 8280 21330 8336
rect 21266 8276 21330 8280
rect 8038 7916 8102 7920
rect 8038 7860 8042 7916
rect 8042 7860 8098 7916
rect 8098 7860 8102 7916
rect 8038 7856 8102 7860
rect 8118 7916 8182 7920
rect 8118 7860 8122 7916
rect 8122 7860 8178 7916
rect 8178 7860 8182 7916
rect 8118 7856 8182 7860
rect 8198 7916 8262 7920
rect 8198 7860 8202 7916
rect 8202 7860 8258 7916
rect 8258 7860 8262 7916
rect 8198 7856 8262 7860
rect 8278 7916 8342 7920
rect 8278 7860 8282 7916
rect 8282 7860 8338 7916
rect 8338 7860 8342 7916
rect 8278 7856 8342 7860
rect 8358 7916 8422 7920
rect 8358 7860 8362 7916
rect 8362 7860 8418 7916
rect 8418 7860 8422 7916
rect 8358 7856 8422 7860
rect 8438 7916 8502 7920
rect 8438 7860 8442 7916
rect 8442 7860 8498 7916
rect 8498 7860 8502 7916
rect 8438 7856 8502 7860
rect 8518 7916 8582 7920
rect 8518 7860 8522 7916
rect 8522 7860 8578 7916
rect 8578 7860 8582 7916
rect 8518 7856 8582 7860
rect 13638 7916 13702 7920
rect 13638 7860 13642 7916
rect 13642 7860 13698 7916
rect 13698 7860 13702 7916
rect 13638 7856 13702 7860
rect 13718 7916 13782 7920
rect 13718 7860 13722 7916
rect 13722 7860 13778 7916
rect 13778 7860 13782 7916
rect 13718 7856 13782 7860
rect 13798 7916 13862 7920
rect 13798 7860 13802 7916
rect 13802 7860 13858 7916
rect 13858 7860 13862 7916
rect 13798 7856 13862 7860
rect 13878 7916 13942 7920
rect 13878 7860 13882 7916
rect 13882 7860 13938 7916
rect 13938 7860 13942 7916
rect 13878 7856 13942 7860
rect 13958 7916 14022 7920
rect 13958 7860 13962 7916
rect 13962 7860 14018 7916
rect 14018 7860 14022 7916
rect 13958 7856 14022 7860
rect 14038 7916 14102 7920
rect 14038 7860 14042 7916
rect 14042 7860 14098 7916
rect 14098 7860 14102 7916
rect 14038 7856 14102 7860
rect 14118 7916 14182 7920
rect 14118 7860 14122 7916
rect 14122 7860 14178 7916
rect 14178 7860 14182 7916
rect 14118 7856 14182 7860
rect 17126 7970 17190 7974
rect 17126 7914 17130 7970
rect 17130 7914 17186 7970
rect 17186 7914 17190 7970
rect 17126 7910 17190 7914
rect 19238 7916 19302 7920
rect 19238 7860 19242 7916
rect 19242 7860 19298 7916
rect 19298 7860 19302 7916
rect 19238 7856 19302 7860
rect 19318 7916 19382 7920
rect 19318 7860 19322 7916
rect 19322 7860 19378 7916
rect 19378 7860 19382 7916
rect 19318 7856 19382 7860
rect 19398 7916 19462 7920
rect 19398 7860 19402 7916
rect 19402 7860 19458 7916
rect 19458 7860 19462 7916
rect 19398 7856 19462 7860
rect 19478 7916 19542 7920
rect 19478 7860 19482 7916
rect 19482 7860 19538 7916
rect 19538 7860 19542 7916
rect 19478 7856 19542 7860
rect 19558 7916 19622 7920
rect 19558 7860 19562 7916
rect 19562 7860 19618 7916
rect 19618 7860 19622 7916
rect 19558 7856 19622 7860
rect 19638 7916 19702 7920
rect 19638 7860 19642 7916
rect 19642 7860 19698 7916
rect 19698 7860 19702 7916
rect 19638 7856 19702 7860
rect 19718 7916 19782 7920
rect 19718 7860 19722 7916
rect 19722 7860 19778 7916
rect 19778 7860 19782 7916
rect 19718 7856 19782 7860
rect 9278 7372 9342 7376
rect 9278 7316 9282 7372
rect 9282 7316 9338 7372
rect 9338 7316 9342 7372
rect 9278 7312 9342 7316
rect 9358 7372 9422 7376
rect 9358 7316 9362 7372
rect 9362 7316 9418 7372
rect 9418 7316 9422 7372
rect 9358 7312 9422 7316
rect 9438 7372 9502 7376
rect 9438 7316 9442 7372
rect 9442 7316 9498 7372
rect 9498 7316 9502 7372
rect 9438 7312 9502 7316
rect 9518 7372 9582 7376
rect 9518 7316 9522 7372
rect 9522 7316 9578 7372
rect 9578 7316 9582 7372
rect 9518 7312 9582 7316
rect 9598 7372 9662 7376
rect 9598 7316 9602 7372
rect 9602 7316 9658 7372
rect 9658 7316 9662 7372
rect 9598 7312 9662 7316
rect 9678 7372 9742 7376
rect 9678 7316 9682 7372
rect 9682 7316 9738 7372
rect 9738 7316 9742 7372
rect 9678 7312 9742 7316
rect 9758 7372 9822 7376
rect 9758 7316 9762 7372
rect 9762 7316 9818 7372
rect 9818 7316 9822 7372
rect 9758 7312 9822 7316
rect 14878 7372 14942 7376
rect 14878 7316 14882 7372
rect 14882 7316 14938 7372
rect 14938 7316 14942 7372
rect 14878 7312 14942 7316
rect 14958 7372 15022 7376
rect 14958 7316 14962 7372
rect 14962 7316 15018 7372
rect 15018 7316 15022 7372
rect 14958 7312 15022 7316
rect 15038 7372 15102 7376
rect 15038 7316 15042 7372
rect 15042 7316 15098 7372
rect 15098 7316 15102 7372
rect 15038 7312 15102 7316
rect 15118 7372 15182 7376
rect 15118 7316 15122 7372
rect 15122 7316 15178 7372
rect 15178 7316 15182 7372
rect 15118 7312 15182 7316
rect 15198 7372 15262 7376
rect 15198 7316 15202 7372
rect 15202 7316 15258 7372
rect 15258 7316 15262 7372
rect 15198 7312 15262 7316
rect 15278 7372 15342 7376
rect 15278 7316 15282 7372
rect 15282 7316 15338 7372
rect 15338 7316 15342 7372
rect 15278 7312 15342 7316
rect 15358 7372 15422 7376
rect 15358 7316 15362 7372
rect 15362 7316 15418 7372
rect 15418 7316 15422 7372
rect 15358 7312 15422 7316
rect 20478 7372 20542 7376
rect 20478 7316 20482 7372
rect 20482 7316 20538 7372
rect 20538 7316 20542 7372
rect 20478 7312 20542 7316
rect 20558 7372 20622 7376
rect 20558 7316 20562 7372
rect 20562 7316 20618 7372
rect 20618 7316 20622 7372
rect 20558 7312 20622 7316
rect 20638 7372 20702 7376
rect 20638 7316 20642 7372
rect 20642 7316 20698 7372
rect 20698 7316 20702 7372
rect 20638 7312 20702 7316
rect 20718 7372 20782 7376
rect 20718 7316 20722 7372
rect 20722 7316 20778 7372
rect 20778 7316 20782 7372
rect 20718 7312 20782 7316
rect 20798 7372 20862 7376
rect 20798 7316 20802 7372
rect 20802 7316 20858 7372
rect 20858 7316 20862 7372
rect 20798 7312 20862 7316
rect 20878 7372 20942 7376
rect 20878 7316 20882 7372
rect 20882 7316 20938 7372
rect 20938 7316 20942 7372
rect 20878 7312 20942 7316
rect 20958 7372 21022 7376
rect 20958 7316 20962 7372
rect 20962 7316 21018 7372
rect 21018 7316 21022 7372
rect 20958 7312 21022 7316
rect 8038 6828 8102 6832
rect 8038 6772 8042 6828
rect 8042 6772 8098 6828
rect 8098 6772 8102 6828
rect 8038 6768 8102 6772
rect 8118 6828 8182 6832
rect 8118 6772 8122 6828
rect 8122 6772 8178 6828
rect 8178 6772 8182 6828
rect 8118 6768 8182 6772
rect 8198 6828 8262 6832
rect 8198 6772 8202 6828
rect 8202 6772 8258 6828
rect 8258 6772 8262 6828
rect 8198 6768 8262 6772
rect 8278 6828 8342 6832
rect 8278 6772 8282 6828
rect 8282 6772 8338 6828
rect 8338 6772 8342 6828
rect 8278 6768 8342 6772
rect 8358 6828 8422 6832
rect 8358 6772 8362 6828
rect 8362 6772 8418 6828
rect 8418 6772 8422 6828
rect 8358 6768 8422 6772
rect 8438 6828 8502 6832
rect 8438 6772 8442 6828
rect 8442 6772 8498 6828
rect 8498 6772 8502 6828
rect 8438 6768 8502 6772
rect 8518 6828 8582 6832
rect 8518 6772 8522 6828
rect 8522 6772 8578 6828
rect 8578 6772 8582 6828
rect 8518 6768 8582 6772
rect 13638 6828 13702 6832
rect 13638 6772 13642 6828
rect 13642 6772 13698 6828
rect 13698 6772 13702 6828
rect 13638 6768 13702 6772
rect 13718 6828 13782 6832
rect 13718 6772 13722 6828
rect 13722 6772 13778 6828
rect 13778 6772 13782 6828
rect 13718 6768 13782 6772
rect 13798 6828 13862 6832
rect 13798 6772 13802 6828
rect 13802 6772 13858 6828
rect 13858 6772 13862 6828
rect 13798 6768 13862 6772
rect 13878 6828 13942 6832
rect 13878 6772 13882 6828
rect 13882 6772 13938 6828
rect 13938 6772 13942 6828
rect 13878 6768 13942 6772
rect 13958 6828 14022 6832
rect 13958 6772 13962 6828
rect 13962 6772 14018 6828
rect 14018 6772 14022 6828
rect 13958 6768 14022 6772
rect 14038 6828 14102 6832
rect 14038 6772 14042 6828
rect 14042 6772 14098 6828
rect 14098 6772 14102 6828
rect 14038 6768 14102 6772
rect 14118 6828 14182 6832
rect 14118 6772 14122 6828
rect 14122 6772 14178 6828
rect 14178 6772 14182 6828
rect 14118 6768 14182 6772
rect 19238 6828 19302 6832
rect 19238 6772 19242 6828
rect 19242 6772 19298 6828
rect 19298 6772 19302 6828
rect 19238 6768 19302 6772
rect 19318 6828 19382 6832
rect 19318 6772 19322 6828
rect 19322 6772 19378 6828
rect 19378 6772 19382 6828
rect 19318 6768 19382 6772
rect 19398 6828 19462 6832
rect 19398 6772 19402 6828
rect 19402 6772 19458 6828
rect 19458 6772 19462 6828
rect 19398 6768 19462 6772
rect 19478 6828 19542 6832
rect 19478 6772 19482 6828
rect 19482 6772 19538 6828
rect 19538 6772 19542 6828
rect 19478 6768 19542 6772
rect 19558 6828 19622 6832
rect 19558 6772 19562 6828
rect 19562 6772 19618 6828
rect 19618 6772 19622 6828
rect 19558 6768 19622 6772
rect 19638 6828 19702 6832
rect 19638 6772 19642 6828
rect 19642 6772 19698 6828
rect 19698 6772 19702 6828
rect 19638 6768 19702 6772
rect 19718 6828 19782 6832
rect 19718 6772 19722 6828
rect 19722 6772 19778 6828
rect 19778 6772 19782 6828
rect 19718 6768 19782 6772
rect 9278 6284 9342 6288
rect 9278 6228 9282 6284
rect 9282 6228 9338 6284
rect 9338 6228 9342 6284
rect 9278 6224 9342 6228
rect 9358 6284 9422 6288
rect 9358 6228 9362 6284
rect 9362 6228 9418 6284
rect 9418 6228 9422 6284
rect 9358 6224 9422 6228
rect 9438 6284 9502 6288
rect 9438 6228 9442 6284
rect 9442 6228 9498 6284
rect 9498 6228 9502 6284
rect 9438 6224 9502 6228
rect 9518 6284 9582 6288
rect 9518 6228 9522 6284
rect 9522 6228 9578 6284
rect 9578 6228 9582 6284
rect 9518 6224 9582 6228
rect 9598 6284 9662 6288
rect 9598 6228 9602 6284
rect 9602 6228 9658 6284
rect 9658 6228 9662 6284
rect 9598 6224 9662 6228
rect 9678 6284 9742 6288
rect 9678 6228 9682 6284
rect 9682 6228 9738 6284
rect 9738 6228 9742 6284
rect 9678 6224 9742 6228
rect 9758 6284 9822 6288
rect 9758 6228 9762 6284
rect 9762 6228 9818 6284
rect 9818 6228 9822 6284
rect 9758 6224 9822 6228
rect 14878 6284 14942 6288
rect 14878 6228 14882 6284
rect 14882 6228 14938 6284
rect 14938 6228 14942 6284
rect 14878 6224 14942 6228
rect 14958 6284 15022 6288
rect 14958 6228 14962 6284
rect 14962 6228 15018 6284
rect 15018 6228 15022 6284
rect 14958 6224 15022 6228
rect 15038 6284 15102 6288
rect 15038 6228 15042 6284
rect 15042 6228 15098 6284
rect 15098 6228 15102 6284
rect 15038 6224 15102 6228
rect 15118 6284 15182 6288
rect 15118 6228 15122 6284
rect 15122 6228 15178 6284
rect 15178 6228 15182 6284
rect 15118 6224 15182 6228
rect 15198 6284 15262 6288
rect 15198 6228 15202 6284
rect 15202 6228 15258 6284
rect 15258 6228 15262 6284
rect 15198 6224 15262 6228
rect 15278 6284 15342 6288
rect 15278 6228 15282 6284
rect 15282 6228 15338 6284
rect 15338 6228 15342 6284
rect 15278 6224 15342 6228
rect 15358 6284 15422 6288
rect 15358 6228 15362 6284
rect 15362 6228 15418 6284
rect 15418 6228 15422 6284
rect 15358 6224 15422 6228
rect 20478 6284 20542 6288
rect 20478 6228 20482 6284
rect 20482 6228 20538 6284
rect 20538 6228 20542 6284
rect 20478 6224 20542 6228
rect 20558 6284 20622 6288
rect 20558 6228 20562 6284
rect 20562 6228 20618 6284
rect 20618 6228 20622 6284
rect 20558 6224 20622 6228
rect 20638 6284 20702 6288
rect 20638 6228 20642 6284
rect 20642 6228 20698 6284
rect 20698 6228 20702 6284
rect 20638 6224 20702 6228
rect 20718 6284 20782 6288
rect 20718 6228 20722 6284
rect 20722 6228 20778 6284
rect 20778 6228 20782 6284
rect 20718 6224 20782 6228
rect 20798 6284 20862 6288
rect 20798 6228 20802 6284
rect 20802 6228 20858 6284
rect 20858 6228 20862 6284
rect 20798 6224 20862 6228
rect 20878 6284 20942 6288
rect 20878 6228 20882 6284
rect 20882 6228 20938 6284
rect 20938 6228 20942 6284
rect 20878 6224 20942 6228
rect 20958 6284 21022 6288
rect 20958 6228 20962 6284
rect 20962 6228 21018 6284
rect 21018 6228 21022 6284
rect 20958 6224 21022 6228
rect 8038 5740 8102 5744
rect 8038 5684 8042 5740
rect 8042 5684 8098 5740
rect 8098 5684 8102 5740
rect 8038 5680 8102 5684
rect 8118 5740 8182 5744
rect 8118 5684 8122 5740
rect 8122 5684 8178 5740
rect 8178 5684 8182 5740
rect 8118 5680 8182 5684
rect 8198 5740 8262 5744
rect 8198 5684 8202 5740
rect 8202 5684 8258 5740
rect 8258 5684 8262 5740
rect 8198 5680 8262 5684
rect 8278 5740 8342 5744
rect 8278 5684 8282 5740
rect 8282 5684 8338 5740
rect 8338 5684 8342 5740
rect 8278 5680 8342 5684
rect 8358 5740 8422 5744
rect 8358 5684 8362 5740
rect 8362 5684 8418 5740
rect 8418 5684 8422 5740
rect 8358 5680 8422 5684
rect 8438 5740 8502 5744
rect 8438 5684 8442 5740
rect 8442 5684 8498 5740
rect 8498 5684 8502 5740
rect 8438 5680 8502 5684
rect 8518 5740 8582 5744
rect 8518 5684 8522 5740
rect 8522 5684 8578 5740
rect 8578 5684 8582 5740
rect 8518 5680 8582 5684
rect 13638 5740 13702 5744
rect 13638 5684 13642 5740
rect 13642 5684 13698 5740
rect 13698 5684 13702 5740
rect 13638 5680 13702 5684
rect 13718 5740 13782 5744
rect 13718 5684 13722 5740
rect 13722 5684 13778 5740
rect 13778 5684 13782 5740
rect 13718 5680 13782 5684
rect 13798 5740 13862 5744
rect 13798 5684 13802 5740
rect 13802 5684 13858 5740
rect 13858 5684 13862 5740
rect 13798 5680 13862 5684
rect 13878 5740 13942 5744
rect 13878 5684 13882 5740
rect 13882 5684 13938 5740
rect 13938 5684 13942 5740
rect 13878 5680 13942 5684
rect 13958 5740 14022 5744
rect 13958 5684 13962 5740
rect 13962 5684 14018 5740
rect 14018 5684 14022 5740
rect 13958 5680 14022 5684
rect 14038 5740 14102 5744
rect 14038 5684 14042 5740
rect 14042 5684 14098 5740
rect 14098 5684 14102 5740
rect 14038 5680 14102 5684
rect 14118 5740 14182 5744
rect 14118 5684 14122 5740
rect 14122 5684 14178 5740
rect 14178 5684 14182 5740
rect 14118 5680 14182 5684
rect 19238 5740 19302 5744
rect 19238 5684 19242 5740
rect 19242 5684 19298 5740
rect 19298 5684 19302 5740
rect 19238 5680 19302 5684
rect 19318 5740 19382 5744
rect 19318 5684 19322 5740
rect 19322 5684 19378 5740
rect 19378 5684 19382 5740
rect 19318 5680 19382 5684
rect 19398 5740 19462 5744
rect 19398 5684 19402 5740
rect 19402 5684 19458 5740
rect 19458 5684 19462 5740
rect 19398 5680 19462 5684
rect 19478 5740 19542 5744
rect 19478 5684 19482 5740
rect 19482 5684 19538 5740
rect 19538 5684 19542 5740
rect 19478 5680 19542 5684
rect 19558 5740 19622 5744
rect 19558 5684 19562 5740
rect 19562 5684 19618 5740
rect 19618 5684 19622 5740
rect 19558 5680 19622 5684
rect 19638 5740 19702 5744
rect 19638 5684 19642 5740
rect 19642 5684 19698 5740
rect 19698 5684 19702 5740
rect 19638 5680 19702 5684
rect 19718 5740 19782 5744
rect 19718 5684 19722 5740
rect 19722 5684 19778 5740
rect 19778 5684 19782 5740
rect 19718 5680 19782 5684
<< metal4 >>
rect 3936 23860 4556 27744
rect 3936 23304 3968 23860
rect 4524 23304 4556 23860
rect 3936 4440 4556 23304
rect 3936 3884 3968 4440
rect 4524 3884 4556 4440
rect 3936 0 4556 3884
rect 5176 22620 5796 27744
rect 5176 22064 5208 22620
rect 5764 22064 5796 22620
rect 5176 5680 5796 22064
rect 5176 5124 5208 5680
rect 5764 5124 5796 5680
rect 5176 0 5796 5124
rect 8000 23860 8620 23892
rect 8000 23304 8032 23860
rect 8588 23304 8620 23860
rect 8000 22064 8620 23304
rect 13600 23860 14220 23892
rect 13600 23304 13632 23860
rect 14188 23304 14220 23860
rect 8000 22000 8038 22064
rect 8102 22000 8118 22064
rect 8182 22000 8198 22064
rect 8262 22000 8278 22064
rect 8342 22000 8358 22064
rect 8422 22000 8438 22064
rect 8502 22000 8518 22064
rect 8582 22000 8620 22064
rect 8000 20976 8620 22000
rect 8000 20912 8038 20976
rect 8102 20912 8118 20976
rect 8182 20912 8198 20976
rect 8262 20912 8278 20976
rect 8342 20912 8358 20976
rect 8422 20912 8438 20976
rect 8502 20912 8518 20976
rect 8582 20912 8620 20976
rect 8000 19888 8620 20912
rect 8000 19824 8038 19888
rect 8102 19824 8118 19888
rect 8182 19824 8198 19888
rect 8262 19824 8278 19888
rect 8342 19824 8358 19888
rect 8422 19824 8438 19888
rect 8502 19824 8518 19888
rect 8582 19824 8620 19888
rect 8000 18800 8620 19824
rect 8000 18736 8038 18800
rect 8102 18736 8118 18800
rect 8182 18736 8198 18800
rect 8262 18736 8278 18800
rect 8342 18736 8358 18800
rect 8422 18736 8438 18800
rect 8502 18736 8518 18800
rect 8582 18736 8620 18800
rect 8000 17712 8620 18736
rect 8000 17648 8038 17712
rect 8102 17648 8118 17712
rect 8182 17648 8198 17712
rect 8262 17648 8278 17712
rect 8342 17648 8358 17712
rect 8422 17648 8438 17712
rect 8502 17648 8518 17712
rect 8582 17648 8620 17712
rect 8000 16624 8620 17648
rect 8000 16560 8038 16624
rect 8102 16560 8118 16624
rect 8182 16560 8198 16624
rect 8262 16560 8278 16624
rect 8342 16560 8358 16624
rect 8422 16560 8438 16624
rect 8502 16560 8518 16624
rect 8582 16560 8620 16624
rect 8000 15536 8620 16560
rect 8000 15472 8038 15536
rect 8102 15472 8118 15536
rect 8182 15472 8198 15536
rect 8262 15472 8278 15536
rect 8342 15472 8358 15536
rect 8422 15472 8438 15536
rect 8502 15472 8518 15536
rect 8582 15472 8620 15536
rect 8000 14448 8620 15472
rect 8000 14384 8038 14448
rect 8102 14384 8118 14448
rect 8182 14384 8198 14448
rect 8262 14384 8278 14448
rect 8342 14384 8358 14448
rect 8422 14384 8438 14448
rect 8502 14384 8518 14448
rect 8582 14384 8620 14448
rect 8000 13360 8620 14384
rect 8000 13296 8038 13360
rect 8102 13296 8118 13360
rect 8182 13296 8198 13360
rect 8262 13296 8278 13360
rect 8342 13296 8358 13360
rect 8422 13296 8438 13360
rect 8502 13296 8518 13360
rect 8582 13296 8620 13360
rect 8000 12272 8620 13296
rect 8000 12208 8038 12272
rect 8102 12208 8118 12272
rect 8182 12208 8198 12272
rect 8262 12208 8278 12272
rect 8342 12208 8358 12272
rect 8422 12208 8438 12272
rect 8502 12208 8518 12272
rect 8582 12208 8620 12272
rect 8000 11184 8620 12208
rect 8000 11120 8038 11184
rect 8102 11120 8118 11184
rect 8182 11120 8198 11184
rect 8262 11120 8278 11184
rect 8342 11120 8358 11184
rect 8422 11120 8438 11184
rect 8502 11120 8518 11184
rect 8582 11120 8620 11184
rect 8000 10096 8620 11120
rect 8000 10032 8038 10096
rect 8102 10032 8118 10096
rect 8182 10032 8198 10096
rect 8262 10032 8278 10096
rect 8342 10032 8358 10096
rect 8422 10032 8438 10096
rect 8502 10032 8518 10096
rect 8582 10032 8620 10096
rect 8000 9008 8620 10032
rect 8000 8944 8038 9008
rect 8102 8944 8118 9008
rect 8182 8944 8198 9008
rect 8262 8944 8278 9008
rect 8342 8944 8358 9008
rect 8422 8944 8438 9008
rect 8502 8944 8518 9008
rect 8582 8944 8620 9008
rect 8000 7920 8620 8944
rect 8000 7856 8038 7920
rect 8102 7856 8118 7920
rect 8182 7856 8198 7920
rect 8262 7856 8278 7920
rect 8342 7856 8358 7920
rect 8422 7856 8438 7920
rect 8502 7856 8518 7920
rect 8582 7856 8620 7920
rect 8000 6832 8620 7856
rect 8000 6768 8038 6832
rect 8102 6768 8118 6832
rect 8182 6768 8198 6832
rect 8262 6768 8278 6832
rect 8342 6768 8358 6832
rect 8422 6768 8438 6832
rect 8502 6768 8518 6832
rect 8582 6768 8620 6832
rect 8000 5744 8620 6768
rect 8000 5680 8038 5744
rect 8102 5680 8118 5744
rect 8182 5680 8198 5744
rect 8262 5680 8278 5744
rect 8342 5680 8358 5744
rect 8422 5680 8438 5744
rect 8502 5680 8518 5744
rect 8582 5680 8620 5744
rect 8000 4440 8620 5680
rect 9240 22620 9860 22652
rect 9240 22064 9272 22620
rect 9828 22064 9860 22620
rect 9240 21520 9860 22064
rect 9240 21456 9278 21520
rect 9342 21456 9358 21520
rect 9422 21456 9438 21520
rect 9502 21456 9518 21520
rect 9582 21456 9598 21520
rect 9662 21456 9678 21520
rect 9742 21456 9758 21520
rect 9822 21456 9860 21520
rect 9240 20432 9860 21456
rect 9240 20368 9278 20432
rect 9342 20368 9358 20432
rect 9422 20368 9438 20432
rect 9502 20368 9518 20432
rect 9582 20368 9598 20432
rect 9662 20368 9678 20432
rect 9742 20368 9758 20432
rect 9822 20368 9860 20432
rect 9240 19344 9860 20368
rect 9240 19280 9278 19344
rect 9342 19280 9358 19344
rect 9422 19280 9438 19344
rect 9502 19280 9518 19344
rect 9582 19280 9598 19344
rect 9662 19280 9678 19344
rect 9742 19280 9758 19344
rect 9822 19280 9860 19344
rect 9240 18256 9860 19280
rect 9240 18192 9278 18256
rect 9342 18192 9358 18256
rect 9422 18192 9438 18256
rect 9502 18192 9518 18256
rect 9582 18192 9598 18256
rect 9662 18192 9678 18256
rect 9742 18192 9758 18256
rect 9822 18192 9860 18256
rect 9240 17168 9860 18192
rect 9240 17104 9278 17168
rect 9342 17104 9358 17168
rect 9422 17104 9438 17168
rect 9502 17104 9518 17168
rect 9582 17104 9598 17168
rect 9662 17104 9678 17168
rect 9742 17104 9758 17168
rect 9822 17104 9860 17168
rect 9240 16080 9860 17104
rect 9240 16016 9278 16080
rect 9342 16016 9358 16080
rect 9422 16016 9438 16080
rect 9502 16016 9518 16080
rect 9582 16016 9598 16080
rect 9662 16016 9678 16080
rect 9742 16016 9758 16080
rect 9822 16016 9860 16080
rect 9240 14992 9860 16016
rect 9240 14928 9278 14992
rect 9342 14928 9358 14992
rect 9422 14928 9438 14992
rect 9502 14928 9518 14992
rect 9582 14928 9598 14992
rect 9662 14928 9678 14992
rect 9742 14928 9758 14992
rect 9822 14928 9860 14992
rect 9240 13904 9860 14928
rect 9240 13840 9278 13904
rect 9342 13840 9358 13904
rect 9422 13840 9438 13904
rect 9502 13840 9518 13904
rect 9582 13840 9598 13904
rect 9662 13840 9678 13904
rect 9742 13840 9758 13904
rect 9822 13840 9860 13904
rect 9240 12816 9860 13840
rect 9240 12752 9278 12816
rect 9342 12752 9358 12816
rect 9422 12752 9438 12816
rect 9502 12752 9518 12816
rect 9582 12752 9598 12816
rect 9662 12752 9678 12816
rect 9742 12752 9758 12816
rect 9822 12752 9860 12816
rect 9240 11728 9860 12752
rect 9240 11664 9278 11728
rect 9342 11664 9358 11728
rect 9422 11664 9438 11728
rect 9502 11664 9518 11728
rect 9582 11664 9598 11728
rect 9662 11664 9678 11728
rect 9742 11664 9758 11728
rect 9822 11664 9860 11728
rect 9240 10640 9860 11664
rect 9240 10576 9278 10640
rect 9342 10576 9358 10640
rect 9422 10576 9438 10640
rect 9502 10576 9518 10640
rect 9582 10576 9598 10640
rect 9662 10576 9678 10640
rect 9742 10576 9758 10640
rect 9822 10576 9860 10640
rect 9240 9552 9860 10576
rect 9240 9488 9278 9552
rect 9342 9488 9358 9552
rect 9422 9488 9438 9552
rect 9502 9488 9518 9552
rect 9582 9488 9598 9552
rect 9662 9488 9678 9552
rect 9742 9488 9758 9552
rect 9822 9488 9860 9552
rect 9240 8464 9860 9488
rect 9240 8400 9278 8464
rect 9342 8400 9358 8464
rect 9422 8400 9438 8464
rect 9502 8400 9518 8464
rect 9582 8400 9598 8464
rect 9662 8400 9678 8464
rect 9742 8400 9758 8464
rect 9822 8400 9860 8464
rect 9240 7376 9860 8400
rect 9240 7312 9278 7376
rect 9342 7312 9358 7376
rect 9422 7312 9438 7376
rect 9502 7312 9518 7376
rect 9582 7312 9598 7376
rect 9662 7312 9678 7376
rect 9742 7312 9758 7376
rect 9822 7312 9860 7376
rect 9240 6288 9860 7312
rect 9240 6224 9278 6288
rect 9342 6224 9358 6288
rect 9422 6224 9438 6288
rect 9502 6224 9518 6288
rect 9582 6224 9598 6288
rect 9662 6224 9678 6288
rect 9742 6224 9758 6288
rect 9822 6224 9860 6288
rect 9240 5680 9860 6224
rect 9240 5124 9272 5680
rect 9828 5124 9860 5680
rect 9240 5092 9860 5124
rect 13600 22064 14220 23304
rect 19200 23860 19820 23892
rect 19200 23304 19232 23860
rect 19788 23304 19820 23860
rect 13600 22000 13638 22064
rect 13702 22000 13718 22064
rect 13782 22000 13798 22064
rect 13862 22000 13878 22064
rect 13942 22000 13958 22064
rect 14022 22000 14038 22064
rect 14102 22000 14118 22064
rect 14182 22000 14220 22064
rect 13600 20976 14220 22000
rect 13600 20912 13638 20976
rect 13702 20912 13718 20976
rect 13782 20912 13798 20976
rect 13862 20912 13878 20976
rect 13942 20912 13958 20976
rect 14022 20912 14038 20976
rect 14102 20912 14118 20976
rect 14182 20912 14220 20976
rect 13600 19888 14220 20912
rect 13600 19824 13638 19888
rect 13702 19824 13718 19888
rect 13782 19824 13798 19888
rect 13862 19824 13878 19888
rect 13942 19824 13958 19888
rect 14022 19824 14038 19888
rect 14102 19824 14118 19888
rect 14182 19824 14220 19888
rect 13600 18800 14220 19824
rect 13600 18736 13638 18800
rect 13702 18736 13718 18800
rect 13782 18736 13798 18800
rect 13862 18736 13878 18800
rect 13942 18736 13958 18800
rect 14022 18736 14038 18800
rect 14102 18736 14118 18800
rect 14182 18736 14220 18800
rect 13600 17712 14220 18736
rect 13600 17648 13638 17712
rect 13702 17648 13718 17712
rect 13782 17648 13798 17712
rect 13862 17648 13878 17712
rect 13942 17648 13958 17712
rect 14022 17648 14038 17712
rect 14102 17648 14118 17712
rect 14182 17648 14220 17712
rect 13600 16624 14220 17648
rect 13600 16560 13638 16624
rect 13702 16560 13718 16624
rect 13782 16560 13798 16624
rect 13862 16560 13878 16624
rect 13942 16560 13958 16624
rect 14022 16560 14038 16624
rect 14102 16560 14118 16624
rect 14182 16560 14220 16624
rect 13600 15536 14220 16560
rect 13600 15472 13638 15536
rect 13702 15472 13718 15536
rect 13782 15472 13798 15536
rect 13862 15472 13878 15536
rect 13942 15472 13958 15536
rect 14022 15472 14038 15536
rect 14102 15472 14118 15536
rect 14182 15472 14220 15536
rect 13600 14448 14220 15472
rect 13600 14384 13638 14448
rect 13702 14384 13718 14448
rect 13782 14384 13798 14448
rect 13862 14384 13878 14448
rect 13942 14384 13958 14448
rect 14022 14384 14038 14448
rect 14102 14384 14118 14448
rect 14182 14384 14220 14448
rect 13600 13360 14220 14384
rect 13600 13296 13638 13360
rect 13702 13296 13718 13360
rect 13782 13296 13798 13360
rect 13862 13296 13878 13360
rect 13942 13296 13958 13360
rect 14022 13296 14038 13360
rect 14102 13296 14118 13360
rect 14182 13296 14220 13360
rect 13600 12272 14220 13296
rect 13600 12208 13638 12272
rect 13702 12208 13718 12272
rect 13782 12208 13798 12272
rect 13862 12208 13878 12272
rect 13942 12208 13958 12272
rect 14022 12208 14038 12272
rect 14102 12208 14118 12272
rect 14182 12208 14220 12272
rect 13600 11184 14220 12208
rect 13600 11120 13638 11184
rect 13702 11120 13718 11184
rect 13782 11120 13798 11184
rect 13862 11120 13878 11184
rect 13942 11120 13958 11184
rect 14022 11120 14038 11184
rect 14102 11120 14118 11184
rect 14182 11120 14220 11184
rect 13600 10096 14220 11120
rect 13600 10032 13638 10096
rect 13702 10032 13718 10096
rect 13782 10032 13798 10096
rect 13862 10032 13878 10096
rect 13942 10032 13958 10096
rect 14022 10032 14038 10096
rect 14102 10032 14118 10096
rect 14182 10032 14220 10096
rect 13600 9008 14220 10032
rect 13600 8944 13638 9008
rect 13702 8944 13718 9008
rect 13782 8944 13798 9008
rect 13862 8944 13878 9008
rect 13942 8944 13958 9008
rect 14022 8944 14038 9008
rect 14102 8944 14118 9008
rect 14182 8944 14220 9008
rect 13600 7920 14220 8944
rect 13600 7856 13638 7920
rect 13702 7856 13718 7920
rect 13782 7856 13798 7920
rect 13862 7856 13878 7920
rect 13942 7856 13958 7920
rect 14022 7856 14038 7920
rect 14102 7856 14118 7920
rect 14182 7856 14220 7920
rect 13600 6832 14220 7856
rect 13600 6768 13638 6832
rect 13702 6768 13718 6832
rect 13782 6768 13798 6832
rect 13862 6768 13878 6832
rect 13942 6768 13958 6832
rect 14022 6768 14038 6832
rect 14102 6768 14118 6832
rect 14182 6768 14220 6832
rect 13600 5744 14220 6768
rect 13600 5680 13638 5744
rect 13702 5680 13718 5744
rect 13782 5680 13798 5744
rect 13862 5680 13878 5744
rect 13942 5680 13958 5744
rect 14022 5680 14038 5744
rect 14102 5680 14118 5744
rect 14182 5680 14220 5744
rect 8000 3884 8032 4440
rect 8588 3884 8620 4440
rect 8000 3852 8620 3884
rect 13600 4440 14220 5680
rect 14840 22620 15460 22652
rect 14840 22064 14872 22620
rect 15428 22064 15460 22620
rect 14840 21520 15460 22064
rect 14840 21456 14878 21520
rect 14942 21456 14958 21520
rect 15022 21456 15038 21520
rect 15102 21456 15118 21520
rect 15182 21456 15198 21520
rect 15262 21456 15278 21520
rect 15342 21456 15358 21520
rect 15422 21456 15460 21520
rect 14840 20432 15460 21456
rect 14840 20368 14878 20432
rect 14942 20368 14958 20432
rect 15022 20368 15038 20432
rect 15102 20368 15118 20432
rect 15182 20368 15198 20432
rect 15262 20368 15278 20432
rect 15342 20368 15358 20432
rect 15422 20368 15460 20432
rect 14840 19344 15460 20368
rect 14840 19280 14878 19344
rect 14942 19280 14958 19344
rect 15022 19280 15038 19344
rect 15102 19280 15118 19344
rect 15182 19280 15198 19344
rect 15262 19280 15278 19344
rect 15342 19280 15358 19344
rect 15422 19280 15460 19344
rect 14840 18256 15460 19280
rect 14840 18192 14878 18256
rect 14942 18192 14958 18256
rect 15022 18192 15038 18256
rect 15102 18192 15118 18256
rect 15182 18192 15198 18256
rect 15262 18192 15278 18256
rect 15342 18192 15358 18256
rect 15422 18192 15460 18256
rect 14840 17168 15460 18192
rect 14840 17104 14878 17168
rect 14942 17104 14958 17168
rect 15022 17104 15038 17168
rect 15102 17104 15118 17168
rect 15182 17104 15198 17168
rect 15262 17104 15278 17168
rect 15342 17104 15358 17168
rect 15422 17104 15460 17168
rect 14840 16080 15460 17104
rect 14840 16016 14878 16080
rect 14942 16016 14958 16080
rect 15022 16016 15038 16080
rect 15102 16016 15118 16080
rect 15182 16016 15198 16080
rect 15262 16016 15278 16080
rect 15342 16016 15358 16080
rect 15422 16016 15460 16080
rect 14840 14992 15460 16016
rect 14840 14928 14878 14992
rect 14942 14928 14958 14992
rect 15022 14928 15038 14992
rect 15102 14928 15118 14992
rect 15182 14928 15198 14992
rect 15262 14928 15278 14992
rect 15342 14928 15358 14992
rect 15422 14928 15460 14992
rect 14840 13904 15460 14928
rect 14840 13840 14878 13904
rect 14942 13840 14958 13904
rect 15022 13840 15038 13904
rect 15102 13840 15118 13904
rect 15182 13840 15198 13904
rect 15262 13840 15278 13904
rect 15342 13840 15358 13904
rect 15422 13840 15460 13904
rect 14840 12816 15460 13840
rect 14840 12752 14878 12816
rect 14942 12752 14958 12816
rect 15022 12752 15038 12816
rect 15102 12752 15118 12816
rect 15182 12752 15198 12816
rect 15262 12752 15278 12816
rect 15342 12752 15358 12816
rect 15422 12752 15460 12816
rect 14840 11728 15460 12752
rect 14840 11664 14878 11728
rect 14942 11664 14958 11728
rect 15022 11664 15038 11728
rect 15102 11664 15118 11728
rect 15182 11664 15198 11728
rect 15262 11664 15278 11728
rect 15342 11664 15358 11728
rect 15422 11664 15460 11728
rect 14840 10640 15460 11664
rect 14840 10576 14878 10640
rect 14942 10576 14958 10640
rect 15022 10576 15038 10640
rect 15102 10576 15118 10640
rect 15182 10576 15198 10640
rect 15262 10576 15278 10640
rect 15342 10576 15358 10640
rect 15422 10576 15460 10640
rect 14840 9552 15460 10576
rect 19200 22064 19820 23304
rect 19200 22000 19238 22064
rect 19302 22000 19318 22064
rect 19382 22000 19398 22064
rect 19462 22000 19478 22064
rect 19542 22000 19558 22064
rect 19622 22000 19638 22064
rect 19702 22000 19718 22064
rect 19782 22000 19820 22064
rect 19200 20976 19820 22000
rect 19200 20912 19238 20976
rect 19302 20912 19318 20976
rect 19382 20912 19398 20976
rect 19462 20912 19478 20976
rect 19542 20912 19558 20976
rect 19622 20912 19638 20976
rect 19702 20912 19718 20976
rect 19782 20912 19820 20976
rect 19200 19888 19820 20912
rect 19200 19824 19238 19888
rect 19302 19824 19318 19888
rect 19382 19824 19398 19888
rect 19462 19824 19478 19888
rect 19542 19824 19558 19888
rect 19622 19824 19638 19888
rect 19702 19824 19718 19888
rect 19782 19824 19820 19888
rect 19200 18800 19820 19824
rect 19200 18736 19238 18800
rect 19302 18736 19318 18800
rect 19382 18736 19398 18800
rect 19462 18736 19478 18800
rect 19542 18736 19558 18800
rect 19622 18736 19638 18800
rect 19702 18736 19718 18800
rect 19782 18736 19820 18800
rect 19200 17712 19820 18736
rect 19200 17648 19238 17712
rect 19302 17648 19318 17712
rect 19382 17648 19398 17712
rect 19462 17648 19478 17712
rect 19542 17648 19558 17712
rect 19622 17648 19638 17712
rect 19702 17648 19718 17712
rect 19782 17648 19820 17712
rect 19200 16624 19820 17648
rect 19200 16560 19238 16624
rect 19302 16560 19318 16624
rect 19382 16560 19398 16624
rect 19462 16560 19478 16624
rect 19542 16560 19558 16624
rect 19622 16560 19638 16624
rect 19702 16560 19718 16624
rect 19782 16560 19820 16624
rect 19200 15536 19820 16560
rect 19200 15472 19238 15536
rect 19302 15472 19318 15536
rect 19382 15472 19398 15536
rect 19462 15472 19478 15536
rect 19542 15472 19558 15536
rect 19622 15472 19638 15536
rect 19702 15472 19718 15536
rect 19782 15472 19820 15536
rect 19200 14448 19820 15472
rect 19200 14384 19238 14448
rect 19302 14384 19318 14448
rect 19382 14384 19398 14448
rect 19462 14384 19478 14448
rect 19542 14384 19558 14448
rect 19622 14384 19638 14448
rect 19702 14384 19718 14448
rect 19782 14384 19820 14448
rect 19200 13360 19820 14384
rect 19200 13296 19238 13360
rect 19302 13296 19318 13360
rect 19382 13296 19398 13360
rect 19462 13296 19478 13360
rect 19542 13296 19558 13360
rect 19622 13296 19638 13360
rect 19702 13296 19718 13360
rect 19782 13296 19820 13360
rect 19200 12272 19820 13296
rect 19200 12208 19238 12272
rect 19302 12208 19318 12272
rect 19382 12208 19398 12272
rect 19462 12208 19478 12272
rect 19542 12208 19558 12272
rect 19622 12208 19638 12272
rect 19702 12208 19718 12272
rect 19782 12208 19820 12272
rect 19200 11184 19820 12208
rect 19200 11120 19238 11184
rect 19302 11120 19318 11184
rect 19382 11120 19398 11184
rect 19462 11120 19478 11184
rect 19542 11120 19558 11184
rect 19622 11120 19638 11184
rect 19702 11120 19718 11184
rect 19782 11120 19820 11184
rect 19200 10096 19820 11120
rect 19200 10032 19238 10096
rect 19302 10032 19318 10096
rect 19382 10032 19398 10096
rect 19462 10032 19478 10096
rect 19542 10032 19558 10096
rect 19622 10032 19638 10096
rect 19702 10032 19718 10096
rect 19782 10032 19820 10096
rect 14840 9488 14878 9552
rect 14942 9488 14958 9552
rect 15022 9488 15038 9552
rect 15102 9488 15118 9552
rect 15182 9488 15198 9552
rect 15262 9488 15278 9552
rect 15342 9488 15358 9552
rect 15422 9488 15460 9552
rect 17125 9560 17191 9561
rect 17125 9496 17126 9560
rect 17190 9496 17191 9560
rect 17125 9495 17191 9496
rect 14840 8464 15460 9488
rect 14840 8400 14878 8464
rect 14942 8400 14958 8464
rect 15022 8400 15038 8464
rect 15102 8400 15118 8464
rect 15182 8400 15198 8464
rect 15262 8400 15278 8464
rect 15342 8400 15358 8464
rect 15422 8400 15460 8464
rect 14840 7376 15460 8400
rect 17128 7975 17188 9495
rect 19200 9008 19820 10032
rect 19200 8944 19238 9008
rect 19302 8944 19318 9008
rect 19382 8944 19398 9008
rect 19462 8944 19478 9008
rect 19542 8944 19558 9008
rect 19622 8944 19638 9008
rect 19702 8944 19718 9008
rect 19782 8944 19820 9008
rect 17125 7974 17191 7975
rect 17125 7910 17126 7974
rect 17190 7910 17191 7974
rect 17125 7909 17191 7910
rect 19200 7920 19820 8944
rect 14840 7312 14878 7376
rect 14942 7312 14958 7376
rect 15022 7312 15038 7376
rect 15102 7312 15118 7376
rect 15182 7312 15198 7376
rect 15262 7312 15278 7376
rect 15342 7312 15358 7376
rect 15422 7312 15460 7376
rect 14840 6288 15460 7312
rect 14840 6224 14878 6288
rect 14942 6224 14958 6288
rect 15022 6224 15038 6288
rect 15102 6224 15118 6288
rect 15182 6224 15198 6288
rect 15262 6224 15278 6288
rect 15342 6224 15358 6288
rect 15422 6224 15460 6288
rect 14840 5680 15460 6224
rect 14840 5124 14872 5680
rect 15428 5124 15460 5680
rect 14840 5092 15460 5124
rect 19200 7856 19238 7920
rect 19302 7856 19318 7920
rect 19382 7856 19398 7920
rect 19462 7856 19478 7920
rect 19542 7856 19558 7920
rect 19622 7856 19638 7920
rect 19702 7856 19718 7920
rect 19782 7856 19820 7920
rect 19200 6832 19820 7856
rect 19200 6768 19238 6832
rect 19302 6768 19318 6832
rect 19382 6768 19398 6832
rect 19462 6768 19478 6832
rect 19542 6768 19558 6832
rect 19622 6768 19638 6832
rect 19702 6768 19718 6832
rect 19782 6768 19820 6832
rect 19200 5744 19820 6768
rect 19200 5680 19238 5744
rect 19302 5680 19318 5744
rect 19382 5680 19398 5744
rect 19462 5680 19478 5744
rect 19542 5680 19558 5744
rect 19622 5680 19638 5744
rect 19702 5680 19718 5744
rect 19782 5680 19820 5744
rect 13600 3884 13632 4440
rect 14188 3884 14220 4440
rect 13600 3852 14220 3884
rect 19200 4440 19820 5680
rect 20440 22620 21060 22652
rect 20440 22064 20472 22620
rect 21028 22064 21060 22620
rect 20440 21520 21060 22064
rect 20440 21456 20478 21520
rect 20542 21456 20558 21520
rect 20622 21456 20638 21520
rect 20702 21456 20718 21520
rect 20782 21456 20798 21520
rect 20862 21456 20878 21520
rect 20942 21456 20958 21520
rect 21022 21456 21060 21520
rect 20440 20432 21060 21456
rect 20440 20368 20478 20432
rect 20542 20368 20558 20432
rect 20622 20368 20638 20432
rect 20702 20368 20718 20432
rect 20782 20368 20798 20432
rect 20862 20368 20878 20432
rect 20942 20368 20958 20432
rect 21022 20368 21060 20432
rect 20440 19344 21060 20368
rect 20440 19280 20478 19344
rect 20542 19280 20558 19344
rect 20622 19280 20638 19344
rect 20702 19280 20718 19344
rect 20782 19280 20798 19344
rect 20862 19280 20878 19344
rect 20942 19280 20958 19344
rect 21022 19280 21060 19344
rect 20440 18256 21060 19280
rect 20440 18192 20478 18256
rect 20542 18192 20558 18256
rect 20622 18192 20638 18256
rect 20702 18192 20718 18256
rect 20782 18192 20798 18256
rect 20862 18192 20878 18256
rect 20942 18192 20958 18256
rect 21022 18192 21060 18256
rect 20440 17168 21060 18192
rect 20440 17104 20478 17168
rect 20542 17104 20558 17168
rect 20622 17104 20638 17168
rect 20702 17104 20718 17168
rect 20782 17104 20798 17168
rect 20862 17104 20878 17168
rect 20942 17104 20958 17168
rect 21022 17104 21060 17168
rect 20440 16080 21060 17104
rect 23000 22620 23620 27744
rect 23000 22064 23032 22620
rect 23588 22064 23620 22620
rect 21265 16392 21331 16393
rect 21265 16328 21266 16392
rect 21330 16328 21331 16392
rect 21265 16327 21331 16328
rect 20440 16016 20478 16080
rect 20542 16016 20558 16080
rect 20622 16016 20638 16080
rect 20702 16016 20718 16080
rect 20782 16016 20798 16080
rect 20862 16016 20878 16080
rect 20942 16016 20958 16080
rect 21022 16016 21060 16080
rect 20440 14992 21060 16016
rect 21268 16024 21328 16327
rect 21268 15964 21604 16024
rect 20440 14928 20478 14992
rect 20542 14928 20558 14992
rect 20622 14928 20638 14992
rect 20702 14928 20718 14992
rect 20782 14928 20798 14992
rect 20862 14928 20878 14992
rect 20942 14928 20958 14992
rect 21022 14928 21060 14992
rect 20440 13904 21060 14928
rect 20440 13840 20478 13904
rect 20542 13840 20558 13904
rect 20622 13840 20638 13904
rect 20702 13840 20718 13904
rect 20782 13840 20798 13904
rect 20862 13840 20878 13904
rect 20942 13840 20958 13904
rect 21022 13840 21060 13904
rect 20440 12816 21060 13840
rect 20440 12752 20478 12816
rect 20542 12752 20558 12816
rect 20622 12752 20638 12816
rect 20702 12752 20718 12816
rect 20782 12752 20798 12816
rect 20862 12752 20878 12816
rect 20942 12752 20958 12816
rect 21022 12752 21060 12816
rect 20440 11728 21060 12752
rect 21544 12364 21604 15964
rect 21268 12304 21604 12364
rect 21268 12001 21328 12304
rect 21265 12000 21331 12001
rect 21265 11936 21266 12000
rect 21330 11936 21331 12000
rect 21265 11935 21331 11936
rect 20440 11664 20478 11728
rect 20542 11664 20558 11728
rect 20622 11664 20638 11728
rect 20702 11664 20718 11728
rect 20782 11664 20798 11728
rect 20862 11664 20878 11728
rect 20942 11664 20958 11728
rect 21022 11664 21060 11728
rect 20440 10640 21060 11664
rect 21268 11632 21328 11935
rect 21268 11572 21466 11632
rect 20440 10576 20478 10640
rect 20542 10576 20558 10640
rect 20622 10576 20638 10640
rect 20702 10576 20718 10640
rect 20782 10576 20798 10640
rect 20862 10576 20878 10640
rect 20942 10576 20958 10640
rect 21022 10576 21060 10640
rect 20440 9552 21060 10576
rect 20440 9488 20478 9552
rect 20542 9488 20558 9552
rect 20622 9488 20638 9552
rect 20702 9488 20718 9552
rect 20782 9488 20798 9552
rect 20862 9488 20878 9552
rect 20942 9488 20958 9552
rect 21022 9488 21060 9552
rect 20440 8464 21060 9488
rect 21406 8704 21466 11572
rect 20440 8400 20478 8464
rect 20542 8400 20558 8464
rect 20622 8400 20638 8464
rect 20702 8400 20718 8464
rect 20782 8400 20798 8464
rect 20862 8400 20878 8464
rect 20942 8400 20958 8464
rect 21022 8400 21060 8464
rect 20440 7376 21060 8400
rect 21268 8644 21466 8704
rect 21268 8341 21328 8644
rect 21265 8340 21331 8341
rect 21265 8276 21266 8340
rect 21330 8276 21331 8340
rect 21265 8275 21331 8276
rect 20440 7312 20478 7376
rect 20542 7312 20558 7376
rect 20622 7312 20638 7376
rect 20702 7312 20718 7376
rect 20782 7312 20798 7376
rect 20862 7312 20878 7376
rect 20942 7312 20958 7376
rect 21022 7312 21060 7376
rect 20440 6288 21060 7312
rect 20440 6224 20478 6288
rect 20542 6224 20558 6288
rect 20622 6224 20638 6288
rect 20702 6224 20718 6288
rect 20782 6224 20798 6288
rect 20862 6224 20878 6288
rect 20942 6224 20958 6288
rect 21022 6224 21060 6288
rect 20440 5680 21060 6224
rect 20440 5124 20472 5680
rect 21028 5124 21060 5680
rect 20440 5092 21060 5124
rect 23000 5680 23620 22064
rect 23000 5124 23032 5680
rect 23588 5124 23620 5680
rect 19200 3884 19232 4440
rect 19788 3884 19820 4440
rect 19200 3852 19820 3884
rect 23000 0 23620 5124
rect 24240 23860 24860 27744
rect 24240 23304 24272 23860
rect 24828 23304 24860 23860
rect 24240 4440 24860 23304
rect 24240 3884 24272 4440
rect 24828 3884 24860 4440
rect 24240 0 24860 3884
<< via4 >>
rect 3968 23304 4524 23860
rect 3968 3884 4524 4440
rect 5208 22064 5764 22620
rect 5208 5124 5764 5680
rect 8032 23304 8588 23860
rect 13632 23304 14188 23860
rect 9272 22064 9828 22620
rect 9272 5124 9828 5680
rect 19232 23304 19788 23860
rect 8032 3884 8588 4440
rect 14872 22064 15428 22620
rect 14872 5124 15428 5680
rect 13632 3884 14188 4440
rect 20472 22064 21028 22620
rect 23032 22064 23588 22620
rect 20472 5124 21028 5680
rect 23032 5124 23588 5680
rect 19232 3884 19788 4440
rect 24272 23304 24828 23860
rect 24272 3884 24828 4440
<< metal5 >>
rect 0 23860 28796 23892
rect 0 23304 3968 23860
rect 4524 23304 8032 23860
rect 8588 23304 13632 23860
rect 14188 23304 19232 23860
rect 19788 23304 24272 23860
rect 24828 23304 28796 23860
rect 0 23272 28796 23304
rect 0 22620 28796 22652
rect 0 22064 5208 22620
rect 5764 22064 9272 22620
rect 9828 22064 14872 22620
rect 15428 22064 20472 22620
rect 21028 22064 23032 22620
rect 23588 22064 28796 22620
rect 0 22032 28796 22064
rect 0 5680 28796 5712
rect 0 5124 5208 5680
rect 5764 5124 9272 5680
rect 9828 5124 14872 5680
rect 15428 5124 20472 5680
rect 21028 5124 23032 5680
rect 23588 5124 28796 5680
rect 0 5092 28796 5124
rect 0 4440 28796 4472
rect 0 3884 3968 4440
rect 4524 3884 8032 4440
rect 8588 3884 13632 4440
rect 14188 3884 19232 4440
rect 19788 3884 24272 4440
rect 24828 3884 28796 4440
rect 0 3852 28796 3884
use digital_filter_VIA3  digital_filter_VIA3_0
timestamp 1654752884
transform 1 0 20750 0 1 21488
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_1
timestamp 1654752884
transform 1 0 20750 0 1 20400
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_2
timestamp 1654752884
transform 1 0 20750 0 1 19312
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_3
timestamp 1654752884
transform 1 0 20750 0 1 18224
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_4
timestamp 1654752884
transform 1 0 20750 0 1 17136
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_5
timestamp 1654752884
transform 1 0 20750 0 1 16048
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_6
timestamp 1654752884
transform 1 0 20750 0 1 14960
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_7
timestamp 1654752884
transform 1 0 20750 0 1 13872
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_8
timestamp 1654752884
transform 1 0 20750 0 1 12784
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_9
timestamp 1654752884
transform 1 0 20750 0 1 11696
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_10
timestamp 1654752884
transform 1 0 20750 0 1 10608
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_11
timestamp 1654752884
transform 1 0 20750 0 1 9520
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_12
timestamp 1654752884
transform 1 0 20750 0 1 8432
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_13
timestamp 1654752884
transform 1 0 20750 0 1 7344
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_14
timestamp 1654752884
transform 1 0 20750 0 1 6256
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_15
timestamp 1654752884
transform 1 0 15150 0 1 21488
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_16
timestamp 1654752884
transform 1 0 15150 0 1 20400
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_17
timestamp 1654752884
transform 1 0 15150 0 1 19312
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_18
timestamp 1654752884
transform 1 0 15150 0 1 18224
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_19
timestamp 1654752884
transform 1 0 15150 0 1 17136
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_20
timestamp 1654752884
transform 1 0 15150 0 1 16048
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_21
timestamp 1654752884
transform 1 0 15150 0 1 14960
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_22
timestamp 1654752884
transform 1 0 15150 0 1 13872
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_23
timestamp 1654752884
transform 1 0 15150 0 1 12784
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_24
timestamp 1654752884
transform 1 0 15150 0 1 11696
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_25
timestamp 1654752884
transform 1 0 15150 0 1 10608
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_26
timestamp 1654752884
transform 1 0 15150 0 1 9520
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_27
timestamp 1654752884
transform 1 0 15150 0 1 8432
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_28
timestamp 1654752884
transform 1 0 15150 0 1 7344
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_29
timestamp 1654752884
transform 1 0 15150 0 1 6256
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_30
timestamp 1654752884
transform 1 0 9550 0 1 21488
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_31
timestamp 1654752884
transform 1 0 9550 0 1 20400
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_32
timestamp 1654752884
transform 1 0 9550 0 1 19312
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_33
timestamp 1654752884
transform 1 0 9550 0 1 18224
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_34
timestamp 1654752884
transform 1 0 9550 0 1 17136
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_35
timestamp 1654752884
transform 1 0 9550 0 1 16048
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_36
timestamp 1654752884
transform 1 0 9550 0 1 14960
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_37
timestamp 1654752884
transform 1 0 9550 0 1 13872
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_38
timestamp 1654752884
transform 1 0 9550 0 1 12784
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_39
timestamp 1654752884
transform 1 0 9550 0 1 11696
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_40
timestamp 1654752884
transform 1 0 9550 0 1 10608
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_41
timestamp 1654752884
transform 1 0 9550 0 1 9520
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_42
timestamp 1654752884
transform 1 0 9550 0 1 8432
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_43
timestamp 1654752884
transform 1 0 9550 0 1 7344
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_44
timestamp 1654752884
transform 1 0 9550 0 1 6256
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_45
timestamp 1654752884
transform 1 0 19510 0 1 22032
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_46
timestamp 1654752884
transform 1 0 19510 0 1 20944
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_47
timestamp 1654752884
transform 1 0 19510 0 1 19856
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_48
timestamp 1654752884
transform 1 0 19510 0 1 18768
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_49
timestamp 1654752884
transform 1 0 19510 0 1 17680
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_50
timestamp 1654752884
transform 1 0 19510 0 1 16592
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_51
timestamp 1654752884
transform 1 0 19510 0 1 15504
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_52
timestamp 1654752884
transform 1 0 19510 0 1 14416
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_53
timestamp 1654752884
transform 1 0 19510 0 1 13328
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_54
timestamp 1654752884
transform 1 0 19510 0 1 12240
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_55
timestamp 1654752884
transform 1 0 19510 0 1 11152
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_56
timestamp 1654752884
transform 1 0 19510 0 1 10064
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_57
timestamp 1654752884
transform 1 0 19510 0 1 8976
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_58
timestamp 1654752884
transform 1 0 19510 0 1 7888
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_59
timestamp 1654752884
transform 1 0 19510 0 1 6800
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_60
timestamp 1654752884
transform 1 0 19510 0 1 5712
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_61
timestamp 1654752884
transform 1 0 13910 0 1 22032
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_62
timestamp 1654752884
transform 1 0 13910 0 1 20944
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_63
timestamp 1654752884
transform 1 0 13910 0 1 19856
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_64
timestamp 1654752884
transform 1 0 13910 0 1 18768
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_65
timestamp 1654752884
transform 1 0 13910 0 1 17680
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_66
timestamp 1654752884
transform 1 0 13910 0 1 16592
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_67
timestamp 1654752884
transform 1 0 13910 0 1 15504
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_68
timestamp 1654752884
transform 1 0 13910 0 1 14416
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_69
timestamp 1654752884
transform 1 0 13910 0 1 13328
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_70
timestamp 1654752884
transform 1 0 13910 0 1 12240
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_71
timestamp 1654752884
transform 1 0 13910 0 1 11152
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_72
timestamp 1654752884
transform 1 0 13910 0 1 10064
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_73
timestamp 1654752884
transform 1 0 13910 0 1 8976
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_74
timestamp 1654752884
transform 1 0 13910 0 1 7888
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_75
timestamp 1654752884
transform 1 0 13910 0 1 6800
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_76
timestamp 1654752884
transform 1 0 13910 0 1 5712
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_77
timestamp 1654752884
transform 1 0 8310 0 1 22032
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_78
timestamp 1654752884
transform 1 0 8310 0 1 20944
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_79
timestamp 1654752884
transform 1 0 8310 0 1 19856
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_80
timestamp 1654752884
transform 1 0 8310 0 1 18768
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_81
timestamp 1654752884
transform 1 0 8310 0 1 17680
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_82
timestamp 1654752884
transform 1 0 8310 0 1 16592
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_83
timestamp 1654752884
transform 1 0 8310 0 1 15504
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_84
timestamp 1654752884
transform 1 0 8310 0 1 14416
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_85
timestamp 1654752884
transform 1 0 8310 0 1 13328
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_86
timestamp 1654752884
transform 1 0 8310 0 1 12240
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_87
timestamp 1654752884
transform 1 0 8310 0 1 11152
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_88
timestamp 1654752884
transform 1 0 8310 0 1 10064
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_89
timestamp 1654752884
transform 1 0 8310 0 1 8976
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_90
timestamp 1654752884
transform 1 0 8310 0 1 7888
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_91
timestamp 1654752884
transform 1 0 8310 0 1 6800
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_92
timestamp 1654752884
transform 1 0 8310 0 1 5712
box -310 -48 310 48
use sky130_fd_sc_hd__a21oi_1  sky130_fd_sc_hd__a21oi_1_0
timestamp 1654752884
transform -1 0 19228 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  sky130_fd_sc_hd__a21oi_1_1
timestamp 1654752884
transform -1 0 15456 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  sky130_fd_sc_hd__a21oi_1_2
timestamp 1654752884
transform 1 0 11224 0 1 18768
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  sky130_fd_sc_hd__a21oi_1_3
timestamp 1654752884
transform 1 0 6348 0 -1 12240
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  sky130_fd_sc_hd__a21oi_1_4
timestamp 1654752884
transform 1 0 6348 0 -1 10064
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  sky130_fd_sc_hd__a21oi_1_5
timestamp 1654752884
transform -1 0 7912 0 -1 6800
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_0
timestamp 1654752884
transform -1 0 20884 0 1 7888
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_1
timestamp 1654752884
transform -1 0 21068 0 1 11152
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_2
timestamp 1654752884
transform -1 0 20884 0 1 10064
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_3
timestamp 1654752884
transform -1 0 20884 0 1 8976
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_4
timestamp 1654752884
transform -1 0 22172 0 -1 13328
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_5
timestamp 1654752884
transform -1 0 20884 0 1 13328
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_6
timestamp 1654752884
transform -1 0 19688 0 -1 14416
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_7
timestamp 1654752884
transform 1 0 20240 0 1 14416
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_8
timestamp 1654752884
transform -1 0 19412 0 1 15504
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_9
timestamp 1654752884
transform 1 0 20516 0 1 16592
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_10
timestamp 1654752884
transform -1 0 19964 0 -1 17680
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_11
timestamp 1654752884
transform 1 0 17480 0 -1 18768
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_12
timestamp 1654752884
transform 1 0 15456 0 1 17680
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_13
timestamp 1654752884
transform 1 0 16652 0 -1 16592
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_14
timestamp 1654752884
transform 1 0 13708 0 1 16592
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_15
timestamp 1654752884
transform -1 0 15732 0 -1 17680
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_16
timestamp 1654752884
transform 1 0 14168 0 -1 14416
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_17
timestamp 1654752884
transform 1 0 16560 0 1 12240
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_18
timestamp 1654752884
transform 1 0 16376 0 -1 15504
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_19
timestamp 1654752884
transform 1 0 16744 0 -1 12240
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_20
timestamp 1654752884
transform -1 0 15732 0 -1 13328
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_21
timestamp 1654752884
transform 1 0 15456 0 1 11152
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_22
timestamp 1654752884
transform -1 0 14628 0 1 10064
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_23
timestamp 1654752884
transform 1 0 15272 0 -1 10064
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_24
timestamp 1654752884
transform -1 0 16836 0 1 8976
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_25
timestamp 1654752884
transform -1 0 18308 0 1 10064
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_26
timestamp 1654752884
transform -1 0 18216 0 -1 12240
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_0
timestamp 1654752884
transform 1 0 10120 0 -1 22032
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_1
timestamp 1654752884
transform 1 0 9016 0 1 15504
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_2
timestamp 1654752884
transform -1 0 10764 0 -1 19856
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_3
timestamp 1654752884
transform 1 0 10212 0 -1 17680
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_4
timestamp 1654752884
transform -1 0 7820 0 1 17680
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_5
timestamp 1654752884
transform -1 0 8280 0 -1 19856
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_6
timestamp 1654752884
transform 1 0 6532 0 1 18768
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_7
timestamp 1654752884
transform 1 0 6348 0 1 17680
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_8
timestamp 1654752884
transform 1 0 8648 0 -1 15504
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_9
timestamp 1654752884
transform 1 0 6624 0 -1 16592
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_10
timestamp 1654752884
transform 1 0 17572 0 1 5712
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_11
timestamp 1654752884
transform 1 0 18768 0 1 6800
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_12
timestamp 1654752884
transform 1 0 15180 0 1 6800
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_13
timestamp 1654752884
transform 1 0 12604 0 -1 8976
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_14
timestamp 1654752884
transform 1 0 12972 0 1 8976
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_15
timestamp 1654752884
transform 1 0 11316 0 1 10064
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_16
timestamp 1654752884
transform 1 0 11408 0 1 11152
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_17
timestamp 1654752884
transform 1 0 12880 0 1 13328
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_18
timestamp 1654752884
transform 1 0 13800 0 1 13328
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_19
timestamp 1654752884
transform 1 0 13616 0 1 14416
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_20
timestamp 1654752884
transform -1 0 13156 0 -1 16592
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_21
timestamp 1654752884
transform -1 0 13340 0 -1 17680
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_22
timestamp 1654752884
transform 1 0 12328 0 -1 19856
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_23
timestamp 1654752884
transform 1 0 15088 0 -1 19856
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_24
timestamp 1654752884
transform 1 0 15916 0 -1 19856
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_25
timestamp 1654752884
transform 1 0 16376 0 -1 19856
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_26
timestamp 1654752884
transform 1 0 21896 0 -1 18768
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_27
timestamp 1654752884
transform 1 0 21528 0 -1 20944
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_28
timestamp 1654752884
transform -1 0 22448 0 -1 16592
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_29
timestamp 1654752884
transform 1 0 22080 0 -1 15504
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_30
timestamp 1654752884
transform 1 0 21620 0 -1 10064
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_31
timestamp 1654752884
transform -1 0 21988 0 -1 12240
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_32
timestamp 1654752884
transform 1 0 21896 0 -1 7888
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_33
timestamp 1654752884
transform 1 0 22080 0 -1 10064
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_34
timestamp 1654752884
transform -1 0 18308 0 1 6800
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_35
timestamp 1654752884
transform 1 0 20700 0 1 6800
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_36
timestamp 1654752884
transform -1 0 22448 0 -1 14416
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_37
timestamp 1654752884
transform -1 0 12788 0 1 5712
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_38
timestamp 1654752884
transform 1 0 12788 0 1 5712
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_39
timestamp 1654752884
transform -1 0 12144 0 -1 7888
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_40
timestamp 1654752884
transform -1 0 11684 0 -1 7888
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_41
timestamp 1654752884
transform 1 0 8832 0 -1 7888
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_42
timestamp 1654752884
transform 1 0 9936 0 -1 10064
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_43
timestamp 1654752884
transform 1 0 8924 0 -1 11152
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_44
timestamp 1654752884
transform -1 0 10304 0 -1 12240
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_45
timestamp 1654752884
transform -1 0 10488 0 -1 13328
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_46
timestamp 1654752884
transform 1 0 9752 0 -1 16592
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_47
timestamp 1654752884
transform 1 0 9200 0 -1 16592
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_48
timestamp 1654752884
transform 1 0 10488 0 1 18768
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_49
timestamp 1654752884
transform -1 0 11868 0 1 17680
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_50
timestamp 1654752884
transform -1 0 13248 0 1 20944
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_51
timestamp 1654752884
transform -1 0 15364 0 -1 20944
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_52
timestamp 1654752884
transform -1 0 16652 0 1 20944
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_53
timestamp 1654752884
transform -1 0 19320 0 1 20944
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_54
timestamp 1654752884
transform -1 0 19780 0 1 20944
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_55
timestamp 1654752884
transform 1 0 19504 0 -1 22032
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_56
timestamp 1654752884
transform 1 0 6440 0 -1 7888
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_57
timestamp 1654752884
transform 1 0 6532 0 1 5712
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_58
timestamp 1654752884
transform 1 0 7820 0 1 5712
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_59
timestamp 1654752884
transform 1 0 6348 0 1 7888
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_60
timestamp 1654752884
transform 1 0 6440 0 1 8976
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_61
timestamp 1654752884
transform 1 0 6624 0 -1 11152
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_62
timestamp 1654752884
transform 1 0 6440 0 1 11152
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_63
timestamp 1654752884
transform 1 0 7268 0 1 13328
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_64
timestamp 1654752884
transform 1 0 6256 0 1 13328
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_0
timestamp 1654752884
transform -1 0 13340 0 -1 8976
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_1
timestamp 1654752884
transform 1 0 13616 0 1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_2
timestamp 1654752884
transform 1 0 10028 0 1 20944
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_3
timestamp 1654752884
transform -1 0 12052 0 -1 19856
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_4
timestamp 1654752884
transform 1 0 11684 0 1 15504
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_5
timestamp 1654752884
transform 1 0 15824 0 1 20944
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_6
timestamp 1654752884
transform 1 0 18032 0 1 20944
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_7
timestamp 1654752884
transform 1 0 6440 0 1 6800
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_8
timestamp 1654752884
transform 1 0 10488 0 1 5712
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_9
timestamp 1654752884
transform -1 0 7084 0 -1 10064
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_10
timestamp 1654752884
transform -1 0 7176 0 1 12240
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  sky130_fd_sc_hd__clkinv_2_0
timestamp 1654752884
transform 1 0 13984 0 1 5712
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_0
timestamp 1654752884
transform 1 0 18032 0 1 13328
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_1
timestamp 1654752884
transform 1 0 17940 0 1 14416
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_8  sky130_fd_sc_hd__clkinv_8_0
timestamp 1654752884
transform 1 0 13892 0 1 7888
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_8  sky130_fd_sc_hd__clkinv_8_1
timestamp 1654752884
transform -1 0 18676 0 -1 6800
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_8  sky130_fd_sc_hd__clkinv_8_2
timestamp 1654752884
transform 1 0 9200 0 1 6800
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_8  sky130_fd_sc_hd__clkinv_8_3
timestamp 1654752884
transform 1 0 18768 0 -1 7888
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_8  sky130_fd_sc_hd__clkinv_8_4
timestamp 1654752884
transform 1 0 20056 0 1 12240
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  sky130_fd_sc_hd__conb_1_0
timestamp 1654752884
transform -1 0 17848 0 -1 15504
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  sky130_fd_sc_hd__conb_1_1
timestamp 1654752884
transform 1 0 14536 0 -1 13328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_0
timestamp 1654752884
transform 1 0 22632 0 -1 20944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_1
timestamp 1654752884
transform 1 0 22632 0 -1 19856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_2
timestamp 1654752884
transform 1 0 22632 0 -1 18768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_3
timestamp 1654752884
transform 1 0 22632 0 -1 17680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_4
timestamp 1654752884
transform 1 0 22632 0 -1 16592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_5
timestamp 1654752884
transform 1 0 22632 0 -1 15504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_6
timestamp 1654752884
transform 1 0 22632 0 -1 14416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_7
timestamp 1654752884
transform 1 0 22632 0 -1 13328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_8
timestamp 1654752884
transform 1 0 22632 0 -1 12240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_9
timestamp 1654752884
transform 1 0 22632 0 -1 11152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_10
timestamp 1654752884
transform 1 0 22632 0 -1 10064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_11
timestamp 1654752884
transform 1 0 22632 0 -1 8976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_12
timestamp 1654752884
transform 1 0 22632 0 -1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_13
timestamp 1654752884
transform 1 0 22632 0 -1 6800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_14
timestamp 1654752884
transform 1 0 22632 0 1 5712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_15
timestamp 1654752884
transform 1 0 21344 0 1 16592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_16
timestamp 1654752884
transform 1 0 20056 0 -1 19856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_17
timestamp 1654752884
transform 1 0 19688 0 -1 14416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_18
timestamp 1654752884
transform 1 0 19228 0 -1 22032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_19
timestamp 1654752884
transform 1 0 18952 0 -1 13328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_20
timestamp 1654752884
transform 1 0 18492 0 -1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_21
timestamp 1654752884
transform 1 0 18216 0 -1 12240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_22
timestamp 1654752884
transform 1 0 17664 0 1 14416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_23
timestamp 1654752884
transform 1 0 17480 0 -1 22032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_24
timestamp 1654752884
transform 1 0 17480 0 -1 20944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_25
timestamp 1654752884
transform 1 0 17480 0 -1 16592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_26
timestamp 1654752884
transform 1 0 17480 0 -1 10064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_27
timestamp 1654752884
transform 1 0 17480 0 -1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_28
timestamp 1654752884
transform 1 0 16928 0 1 18768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_29
timestamp 1654752884
transform 1 0 16928 0 1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_30
timestamp 1654752884
transform 1 0 16192 0 1 15504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_31
timestamp 1654752884
transform 1 0 16376 0 -1 6800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_32
timestamp 1654752884
transform 1 0 15824 0 1 15504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_33
timestamp 1654752884
transform 1 0 14904 0 -1 18768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_34
timestamp 1654752884
transform 1 0 14904 0 -1 14416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_35
timestamp 1654752884
transform 1 0 14904 0 -1 11152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_36
timestamp 1654752884
transform 1 0 14536 0 -1 22032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_37
timestamp 1654752884
transform 1 0 14260 0 -1 13328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_38
timestamp 1654752884
transform 1 0 13800 0 -1 10064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_39
timestamp 1654752884
transform 1 0 13800 0 -1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_40
timestamp 1654752884
transform 1 0 13800 0 -1 6800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_41
timestamp 1654752884
transform 1 0 12328 0 -1 12240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_42
timestamp 1654752884
transform 1 0 12328 0 -1 11152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_43
timestamp 1654752884
transform 1 0 11776 0 1 20944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_44
timestamp 1654752884
transform 1 0 11040 0 -1 22032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_45
timestamp 1654752884
transform 1 0 11224 0 -1 20944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_46
timestamp 1654752884
transform 1 0 11040 0 1 16592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_47
timestamp 1654752884
transform 1 0 11040 0 1 10064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_48
timestamp 1654752884
transform 1 0 10764 0 -1 19856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_49
timestamp 1654752884
transform 1 0 10672 0 1 17680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_50
timestamp 1654752884
transform 1 0 10672 0 1 10064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_51
timestamp 1654752884
transform 1 0 10304 0 -1 12240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_52
timestamp 1654752884
transform 1 0 9752 0 1 20944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_53
timestamp 1654752884
transform 1 0 9752 0 -1 13328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_54
timestamp 1654752884
transform 1 0 9384 0 -1 11152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_55
timestamp 1654752884
transform 1 0 9384 0 -1 10064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_56
timestamp 1654752884
transform 1 0 8464 0 1 16592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_57
timestamp 1654752884
transform 1 0 8096 0 -1 22032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_58
timestamp 1654752884
transform 1 0 8096 0 1 12240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_59
timestamp 1654752884
transform 1 0 8096 0 1 10064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_60
timestamp 1654752884
transform 1 0 7176 0 -1 12240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_61
timestamp 1654752884
transform 1 0 6808 0 -1 14416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_62
timestamp 1654752884
transform 1 0 6808 0 -1 13328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_63
timestamp 1654752884
transform 1 0 6624 0 1 12240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_64
timestamp 1654752884
transform 1 0 5888 0 1 15504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_65
timestamp 1654752884
transform 1 0 5888 0 1 14416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_0
timestamp 1654752884
transform 1 0 22540 0 1 8976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_1
timestamp 1654752884
transform 1 0 22172 0 -1 13328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_2
timestamp 1654752884
transform 1 0 21620 0 -1 16592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_3
timestamp 1654752884
transform 1 0 21620 0 -1 14416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_4
timestamp 1654752884
transform 1 0 21528 0 -1 11152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_5
timestamp 1654752884
transform 1 0 20884 0 1 13328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_6
timestamp 1654752884
transform 1 0 19688 0 1 12240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_7
timestamp 1654752884
transform 1 0 19596 0 -1 6800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_8
timestamp 1654752884
transform 1 0 18308 0 1 20944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_9
timestamp 1654752884
transform 1 0 18308 0 1 16592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_10
timestamp 1654752884
transform 1 0 18308 0 1 11152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_11
timestamp 1654752884
transform 1 0 17756 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_12
timestamp 1654752884
transform 1 0 17480 0 -1 17680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_13
timestamp 1654752884
transform 1 0 17664 0 1 13328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_14
timestamp 1654752884
transform 1 0 17020 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_15
timestamp 1654752884
transform 1 0 17020 0 -1 15504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_16
timestamp 1654752884
transform 1 0 17020 0 -1 8976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_17
timestamp 1654752884
transform 1 0 16652 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_18
timestamp 1654752884
transform 1 0 16284 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_19
timestamp 1654752884
transform 1 0 16192 0 1 12240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_20
timestamp 1654752884
transform 1 0 15640 0 1 19856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_21
timestamp 1654752884
transform 1 0 14904 0 -1 10064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_22
timestamp 1654752884
transform 1 0 14444 0 -1 7888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_23
timestamp 1654752884
transform 1 0 14444 0 1 5712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_24
timestamp 1654752884
transform 1 0 14168 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_25
timestamp 1654752884
transform 1 0 14076 0 1 14416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_26
timestamp 1654752884
transform 1 0 13800 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_27
timestamp 1654752884
transform 1 0 13616 0 1 17680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_28
timestamp 1654752884
transform 1 0 13616 0 1 11152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_29
timestamp 1654752884
transform 1 0 13616 0 1 10064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_30
timestamp 1654752884
transform 1 0 13064 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_31
timestamp 1654752884
transform 1 0 12696 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_32
timestamp 1654752884
transform 1 0 12328 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_33
timestamp 1654752884
transform 1 0 12328 0 -1 16592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_34
timestamp 1654752884
transform 1 0 12328 0 -1 14416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_35
timestamp 1654752884
transform 1 0 12328 0 -1 13328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_36
timestamp 1654752884
transform 1 0 11868 0 1 5712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_37
timestamp 1654752884
transform 1 0 11684 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_38
timestamp 1654752884
transform 1 0 11316 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_39
timestamp 1654752884
transform 1 0 11040 0 1 17680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_40
timestamp 1654752884
transform 1 0 11040 0 1 11152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_41
timestamp 1654752884
transform 1 0 11132 0 1 8976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_42
timestamp 1654752884
transform 1 0 10580 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_43
timestamp 1654752884
transform 1 0 10580 0 1 19856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_44
timestamp 1654752884
transform 1 0 9752 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_45
timestamp 1654752884
transform 1 0 9844 0 -1 17680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_46
timestamp 1654752884
transform 1 0 9292 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_47
timestamp 1654752884
transform 1 0 9292 0 -1 14416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_48
timestamp 1654752884
transform 1 0 9292 0 -1 7888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_49
timestamp 1654752884
transform 1 0 8832 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_50
timestamp 1654752884
transform 1 0 8740 0 -1 17680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_51
timestamp 1654752884
transform 1 0 8464 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_52
timestamp 1654752884
transform 1 0 8464 0 1 17680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_53
timestamp 1654752884
transform 1 0 8464 0 1 5712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_54
timestamp 1654752884
transform 1 0 7728 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_55
timestamp 1654752884
transform 1 0 7360 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_56
timestamp 1654752884
transform 1 0 6716 0 -1 12240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_57
timestamp 1654752884
transform 1 0 6624 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_58
timestamp 1654752884
transform 1 0 6256 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_59
timestamp 1654752884
transform 1 0 5888 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_60
timestamp 1654752884
transform 1 0 5796 0 -1 14416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_61
timestamp 1654752884
transform 1 0 5888 0 1 12240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_62
timestamp 1654752884
transform 1 0 5888 0 1 10064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_63
timestamp 1654752884
transform 1 0 5888 0 1 7888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_0
timestamp 1654752884
transform 1 0 21988 0 -1 20944
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_1
timestamp 1654752884
transform 1 0 21988 0 -1 12240
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_2
timestamp 1654752884
transform 1 0 18124 0 1 17680
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_3
timestamp 1654752884
transform 1 0 18124 0 1 15504
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_4
timestamp 1654752884
transform 1 0 18124 0 1 5712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_5
timestamp 1654752884
transform 1 0 17940 0 -1 15504
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_6
timestamp 1654752884
transform 1 0 16836 0 -1 14416
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_7
timestamp 1654752884
transform 1 0 16192 0 1 16592
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_8
timestamp 1654752884
transform 1 0 16284 0 1 11152
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_9
timestamp 1654752884
transform 1 0 14904 0 -1 8976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_10
timestamp 1654752884
transform 1 0 14260 0 -1 19856
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_11
timestamp 1654752884
transform 1 0 14352 0 1 13328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_12
timestamp 1654752884
transform 1 0 13616 0 1 19856
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_13
timestamp 1654752884
transform 1 0 12328 0 -1 17680
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_14
timestamp 1654752884
transform 1 0 12512 0 1 7888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_15
timestamp 1654752884
transform 1 0 10396 0 1 20944
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_16
timestamp 1654752884
transform 1 0 10396 0 1 12240
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_17
timestamp 1654752884
transform 1 0 10396 0 1 6800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_18
timestamp 1654752884
transform 1 0 9752 0 -1 19856
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_19
timestamp 1654752884
transform 1 0 9844 0 -1 11152
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_20
timestamp 1654752884
transform 1 0 9108 0 -1 15504
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_21
timestamp 1654752884
transform 1 0 8556 0 1 19856
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_22
timestamp 1654752884
transform 1 0 8556 0 1 13328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_23
timestamp 1654752884
transform 1 0 8556 0 1 11152
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_24
timestamp 1654752884
transform 1 0 8556 0 1 10064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_25
timestamp 1654752884
transform 1 0 8556 0 1 8976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_26
timestamp 1654752884
transform 1 0 8556 0 1 7888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_27
timestamp 1654752884
transform 1 0 8556 0 1 6800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_28
timestamp 1654752884
transform 1 0 7820 0 1 13328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_29
timestamp 1654752884
transform 1 0 7268 0 -1 19856
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_30
timestamp 1654752884
transform 1 0 7268 0 -1 14416
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_31
timestamp 1654752884
transform 1 0 7176 0 -1 10064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_32
timestamp 1654752884
transform 1 0 7452 0 -1 8976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_33
timestamp 1654752884
transform 1 0 6808 0 1 17680
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_34
timestamp 1654752884
transform 1 0 5888 0 1 11152
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_35
timestamp 1654752884
transform 1 0 5888 0 1 8976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_36
timestamp 1654752884
transform 1 0 5796 0 -1 8976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_37
timestamp 1654752884
transform 1 0 5980 0 1 5712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_0
timestamp 1654752884
transform 1 0 21804 0 -1 8976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_1
timestamp 1654752884
transform 1 0 20424 0 1 19856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_2
timestamp 1654752884
transform 1 0 20332 0 -1 19856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_3
timestamp 1654752884
transform 1 0 20332 0 -1 17680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_4
timestamp 1654752884
transform 1 0 19228 0 -1 20944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_5
timestamp 1654752884
transform 1 0 19228 0 -1 19856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_6
timestamp 1654752884
transform 1 0 19228 0 -1 13328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_7
timestamp 1654752884
transform 1 0 18860 0 1 18768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_8
timestamp 1654752884
transform 1 0 18860 0 1 17680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_9
timestamp 1654752884
transform 1 0 18860 0 1 12240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_10
timestamp 1654752884
transform 1 0 18860 0 -1 6800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_11
timestamp 1654752884
transform 1 0 18124 0 -1 18768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_12
timestamp 1654752884
transform 1 0 17756 0 1 19856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_13
timestamp 1654752884
transform 1 0 17756 0 -1 16592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_14
timestamp 1654752884
transform 1 0 17572 0 -1 11152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_15
timestamp 1654752884
transform 1 0 17756 0 -1 7888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_16
timestamp 1654752884
transform 1 0 16652 0 -1 17680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_17
timestamp 1654752884
transform 1 0 16652 0 -1 11152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_18
timestamp 1654752884
transform 1 0 16652 0 -1 6800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_19
timestamp 1654752884
transform 1 0 16192 0 1 18768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_20
timestamp 1654752884
transform 1 0 16192 0 1 7888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_21
timestamp 1654752884
transform 1 0 15732 0 -1 17680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_22
timestamp 1654752884
transform 1 0 15364 0 1 7888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_23
timestamp 1654752884
transform 1 0 15180 0 -1 18768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_24
timestamp 1654752884
transform 1 0 15180 0 1 12240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_25
timestamp 1654752884
transform 1 0 15180 0 1 8976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_26
timestamp 1654752884
transform 1 0 14996 0 -1 7888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_27
timestamp 1654752884
transform 1 0 14076 0 -1 18768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_28
timestamp 1654752884
transform 1 0 14076 0 -1 10064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_29
timestamp 1654752884
transform 1 0 14076 0 -1 6800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_30
timestamp 1654752884
transform 1 0 13616 0 1 18768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_31
timestamp 1654752884
transform 1 0 13616 0 1 15504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_32
timestamp 1654752884
transform 1 0 12788 0 1 6800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_33
timestamp 1654752884
transform 1 0 12604 0 1 19856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_34
timestamp 1654752884
transform 1 0 12420 0 -1 15504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_35
timestamp 1654752884
transform 1 0 12604 0 1 14416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_36
timestamp 1654752884
transform 1 0 12604 0 -1 12240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_37
timestamp 1654752884
transform 1 0 12604 0 -1 11152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_38
timestamp 1654752884
transform 1 0 12052 0 1 20944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_39
timestamp 1654752884
transform 1 0 11500 0 -1 20944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_40
timestamp 1654752884
transform 1 0 11040 0 1 20944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_41
timestamp 1654752884
transform 1 0 11040 0 -1 19856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_42
timestamp 1654752884
transform 1 0 11040 0 1 12240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_43
timestamp 1654752884
transform 1 0 11040 0 1 5712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_44
timestamp 1654752884
transform 1 0 9936 0 -1 18768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_45
timestamp 1654752884
transform 1 0 9936 0 -1 14416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_46
timestamp 1654752884
transform 1 0 9752 0 -1 8976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_47
timestamp 1654752884
transform 1 0 9844 0 -1 6800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_48
timestamp 1654752884
transform 1 0 8924 0 -1 20944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_49
timestamp 1654752884
transform 1 0 8648 0 1 18768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_50
timestamp 1654752884
transform 1 0 8832 0 1 17680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_51
timestamp 1654752884
transform 1 0 8740 0 1 16592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_52
timestamp 1654752884
transform 1 0 8924 0 -1 13328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_53
timestamp 1654752884
transform 1 0 8924 0 -1 12240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_54
timestamp 1654752884
transform 1 0 8924 0 1 5712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_55
timestamp 1654752884
transform 1 0 7360 0 1 12240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_56
timestamp 1654752884
transform 1 0 7360 0 1 10064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_57
timestamp 1654752884
transform 1 0 6072 0 1 19856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_58
timestamp 1654752884
transform 1 0 6164 0 1 15504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_59
timestamp 1654752884
transform 1 0 6164 0 1 14416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_60
timestamp 1654752884
transform 1 0 5796 0 -1 13328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_61
timestamp 1654752884
transform 1 0 5796 0 -1 11152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_0
timestamp 1654752884
transform 1 0 21620 0 1 16592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_1
timestamp 1654752884
transform 1 0 14904 0 1 13328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_2
timestamp 1654752884
transform 1 0 14904 0 1 5712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_3
timestamp 1654752884
transform 1 0 8648 0 1 20944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_4
timestamp 1654752884
transform 1 0 7084 0 1 20944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_5
timestamp 1654752884
transform 1 0 7084 0 1 18768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_6
timestamp 1654752884
transform 1 0 7084 0 1 16592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_7
timestamp 1654752884
transform 1 0 5980 0 1 20944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_8
timestamp 1654752884
transform 1 0 5980 0 -1 20944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_9
timestamp 1654752884
transform 1 0 5980 0 -1 19856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_10
timestamp 1654752884
transform 1 0 5980 0 1 16592
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_0
timestamp 1654752884
transform -1 0 12512 0 1 19856
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_1
timestamp 1654752884
transform 1 0 18768 0 1 10064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_2
timestamp 1654752884
transform -1 0 11224 0 -1 7888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_3
timestamp 1654752884
transform -1 0 18676 0 1 12240
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_4
timestamp 1654752884
transform 1 0 18768 0 1 7888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_5
timestamp 1654752884
transform 1 0 18308 0 -1 11152
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_6
timestamp 1654752884
transform 1 0 20056 0 -1 10064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_7
timestamp 1654752884
transform 1 0 18492 0 -1 12240
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_8
timestamp 1654752884
transform 1 0 18768 0 1 13328
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_9
timestamp 1654752884
transform 1 0 18768 0 1 14416
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_10
timestamp 1654752884
transform -1 0 21528 0 -1 15504
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_11
timestamp 1654752884
transform 1 0 18492 0 -1 15504
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_12
timestamp 1654752884
transform -1 0 21160 0 1 15504
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_13
timestamp 1654752884
transform 1 0 18492 0 -1 16592
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_14
timestamp 1654752884
transform 1 0 18768 0 1 16592
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_15
timestamp 1654752884
transform 1 0 16192 0 1 14416
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_16
timestamp 1654752884
transform -1 0 18216 0 1 16592
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_17
timestamp 1654752884
transform 1 0 15088 0 -1 16592
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_18
timestamp 1654752884
transform -1 0 14812 0 -1 16592
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_19
timestamp 1654752884
transform -1 0 18952 0 -1 14416
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_20
timestamp 1654752884
transform -1 0 17664 0 1 13328
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_21
timestamp 1654752884
transform -1 0 18952 0 -1 13328
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_22
timestamp 1654752884
transform -1 0 17388 0 -1 13328
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_23
timestamp 1654752884
transform 1 0 14904 0 -1 12240
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_24
timestamp 1654752884
transform -1 0 17664 0 1 10064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_25
timestamp 1654752884
transform 1 0 13984 0 1 11152
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_26
timestamp 1654752884
transform -1 0 16652 0 -1 11152
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_27
timestamp 1654752884
transform -1 0 16100 0 1 10064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_28
timestamp 1654752884
transform -1 0 18308 0 1 8976
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_29
timestamp 1654752884
transform 1 0 16836 0 1 11152
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_30
timestamp 1654752884
transform 1 0 13616 0 1 6800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_31
timestamp 1654752884
transform 1 0 12328 0 -1 6800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_32
timestamp 1654752884
transform 1 0 15916 0 -1 10064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_33
timestamp 1654752884
transform -1 0 18676 0 1 7888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_34
timestamp 1654752884
transform 1 0 15456 0 -1 8976
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_35
timestamp 1654752884
transform 1 0 13340 0 -1 8976
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_36
timestamp 1654752884
transform 1 0 13616 0 1 8976
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_37
timestamp 1654752884
transform 1 0 13340 0 -1 11152
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_38
timestamp 1654752884
transform 1 0 13340 0 -1 12240
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_39
timestamp 1654752884
transform 1 0 13616 0 1 12240
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_40
timestamp 1654752884
transform 1 0 14904 0 -1 15504
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_41
timestamp 1654752884
transform 1 0 14444 0 1 14416
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_42
timestamp 1654752884
transform 1 0 14352 0 1 15504
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_43
timestamp 1654752884
transform 1 0 13340 0 -1 17680
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_44
timestamp 1654752884
transform 1 0 13984 0 1 17680
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_45
timestamp 1654752884
transform 1 0 14352 0 1 16592
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_46
timestamp 1654752884
transform -1 0 17388 0 -1 18768
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_47
timestamp 1654752884
transform 1 0 17204 0 1 18768
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_48
timestamp 1654752884
transform 1 0 20056 0 -1 18768
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_49
timestamp 1654752884
transform 1 0 19780 0 1 17680
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_50
timestamp 1654752884
transform 1 0 17848 0 -1 17680
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_51
timestamp 1654752884
transform 1 0 20056 0 -1 16592
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_52
timestamp 1654752884
transform -1 0 21620 0 -1 14416
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_53
timestamp 1654752884
transform -1 0 21528 0 -1 13328
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_54
timestamp 1654752884
transform -1 0 21528 0 -1 12240
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_55
timestamp 1654752884
transform 1 0 18768 0 1 8976
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_56
timestamp 1654752884
transform 1 0 21344 0 1 7888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_57
timestamp 1654752884
transform -1 0 21528 0 -1 11152
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_58
timestamp 1654752884
transform 1 0 21344 0 1 10064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_59
timestamp 1654752884
transform -1 0 12236 0 -1 14416
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_60
timestamp 1654752884
transform -1 0 11224 0 -1 20944
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_61
timestamp 1654752884
transform -1 0 10580 0 1 19856
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_62
timestamp 1654752884
transform -1 0 10948 0 1 16592
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_63
timestamp 1654752884
transform 1 0 6900 0 1 15504
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_64
timestamp 1654752884
transform 1 0 7268 0 -1 20944
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_65
timestamp 1654752884
transform 1 0 6808 0 1 19856
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_66
timestamp 1654752884
transform 1 0 7176 0 -1 17680
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_67
timestamp 1654752884
transform -1 0 8648 0 -1 15504
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_68
timestamp 1654752884
transform 1 0 7360 0 -1 16592
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_69
timestamp 1654752884
transform 1 0 21344 0 1 6800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_70
timestamp 1654752884
transform 1 0 19228 0 1 6800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_71
timestamp 1654752884
transform 1 0 16192 0 1 6800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_72
timestamp 1654752884
transform 1 0 12328 0 -1 10064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_73
timestamp 1654752884
transform -1 0 12972 0 1 8976
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_74
timestamp 1654752884
transform 1 0 12052 0 1 10064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_75
timestamp 1654752884
transform 1 0 12052 0 1 11152
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_76
timestamp 1654752884
transform -1 0 13340 0 1 12240
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_77
timestamp 1654752884
transform 1 0 12788 0 -1 13328
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_78
timestamp 1654752884
transform 1 0 12696 0 -1 14416
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_79
timestamp 1654752884
transform 1 0 12052 0 1 15504
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_80
timestamp 1654752884
transform 1 0 10764 0 -1 17680
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_81
timestamp 1654752884
transform 1 0 12788 0 -1 19856
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_82
timestamp 1654752884
transform -1 0 15824 0 1 20944
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_83
timestamp 1654752884
transform 1 0 16192 0 1 19856
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_84
timestamp 1654752884
transform -1 0 20240 0 1 19856
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_85
timestamp 1654752884
transform -1 0 23000 0 1 19856
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_86
timestamp 1654752884
transform -1 0 22816 0 1 17680
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_87
timestamp 1654752884
transform -1 0 22540 0 -1 17680
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_88
timestamp 1654752884
transform -1 0 22816 0 1 14416
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_89
timestamp 1654752884
transform -1 0 22540 0 -1 19856
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_90
timestamp 1654752884
transform 1 0 21344 0 1 12240
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_91
timestamp 1654752884
transform -1 0 22908 0 1 18768
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_92
timestamp 1654752884
transform -1 0 22816 0 1 13328
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_93
timestamp 1654752884
transform 1 0 18768 0 1 11152
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_94
timestamp 1654752884
transform -1 0 22816 0 1 11152
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_95
timestamp 1654752884
transform -1 0 22816 0 1 15504
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_96
timestamp 1654752884
transform 1 0 20056 0 -1 20944
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_97
timestamp 1654752884
transform 1 0 19780 0 1 20944
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_98
timestamp 1654752884
transform -1 0 19228 0 -1 20944
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_99
timestamp 1654752884
transform 1 0 15916 0 -1 20944
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_100
timestamp 1654752884
transform -1 0 15640 0 1 19856
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_101
timestamp 1654752884
transform 1 0 12328 0 -1 20944
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_102
timestamp 1654752884
transform 1 0 10672 0 -1 18768
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_103
timestamp 1654752884
transform 1 0 10304 0 -1 16592
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_104
timestamp 1654752884
transform 1 0 9476 0 1 15504
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_105
timestamp 1654752884
transform -1 0 12512 0 1 14416
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_106
timestamp 1654752884
transform 1 0 7268 0 -1 13328
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_107
timestamp 1654752884
transform 1 0 7452 0 -1 12240
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_108
timestamp 1654752884
transform 1 0 9200 0 1 10064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_109
timestamp 1654752884
transform 1 0 9292 0 1 8976
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_110
timestamp 1654752884
transform 1 0 9292 0 1 7888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_111
timestamp 1654752884
transform 1 0 11040 0 1 7888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_112
timestamp 1654752884
transform 1 0 12328 0 -1 7888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_113
timestamp 1654752884
transform 1 0 14904 0 -1 6800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_114
timestamp 1654752884
transform 1 0 7820 0 -1 14416
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_115
timestamp 1654752884
transform 1 0 6900 0 1 14416
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_116
timestamp 1654752884
transform 1 0 6900 0 1 11152
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_117
timestamp 1654752884
transform 1 0 7268 0 -1 11152
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_118
timestamp 1654752884
transform 1 0 6900 0 1 8976
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_119
timestamp 1654752884
transform 1 0 6900 0 1 7888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_120
timestamp 1654752884
transform 1 0 8188 0 -1 6800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_121
timestamp 1654752884
transform 1 0 6900 0 1 6800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_122
timestamp 1654752884
transform 1 0 7176 0 -1 7888
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_0
timestamp 1654752884
transform 1 0 21344 0 1 20944
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_1
timestamp 1654752884
transform -1 0 21252 0 1 18768
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_2
timestamp 1654752884
transform -1 0 19228 0 -1 19856
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_3
timestamp 1654752884
transform -1 0 16100 0 1 18768
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_4
timestamp 1654752884
transform -1 0 14076 0 -1 18768
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_5
timestamp 1654752884
transform -1 0 13524 0 1 18768
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_6
timestamp 1654752884
transform 1 0 11868 0 1 17680
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_7
timestamp 1654752884
transform 1 0 11868 0 1 16592
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_8
timestamp 1654752884
transform -1 0 12236 0 -1 15504
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_9
timestamp 1654752884
transform 1 0 11132 0 1 13328
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_10
timestamp 1654752884
transform 1 0 10580 0 -1 13328
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_11
timestamp 1654752884
transform 1 0 10580 0 -1 12240
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_12
timestamp 1654752884
transform 1 0 10396 0 -1 11152
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_13
timestamp 1654752884
transform 1 0 10580 0 -1 10064
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_14
timestamp 1654752884
transform 1 0 10488 0 -1 8976
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_15
timestamp 1654752884
transform 1 0 20056 0 -1 8976
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_16
timestamp 1654752884
transform 1 0 20056 0 -1 7888
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_17
timestamp 1654752884
transform -1 0 10488 0 1 14416
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_18
timestamp 1654752884
transform 1 0 9200 0 1 13328
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_19
timestamp 1654752884
transform 1 0 8648 0 1 12240
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_20
timestamp 1654752884
transform -1 0 10764 0 1 11152
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_21
timestamp 1654752884
transform -1 0 9384 0 -1 10064
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_22
timestamp 1654752884
transform -1 0 9660 0 -1 8976
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_23
timestamp 1654752884
transform 1 0 10580 0 -1 6800
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_24
timestamp 1654752884
transform 1 0 11040 0 1 6800
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_0
timestamp 1654752884
transform 1 0 18124 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_1
timestamp 1654752884
transform 1 0 16192 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_2
timestamp 1654752884
transform 1 0 12052 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_3
timestamp 1654752884
transform 1 0 9200 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_4
timestamp 1654752884
transform 1 0 10304 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_5
timestamp 1654752884
transform 1 0 8188 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_6
timestamp 1654752884
transform 1 0 5888 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_7
timestamp 1654752884
transform 1 0 22908 0 -1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_8
timestamp 1654752884
transform 1 0 18492 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_9
timestamp 1654752884
transform 1 0 17664 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_10
timestamp 1654752884
transform 1 0 13340 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_11
timestamp 1654752884
transform 1 0 12512 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_12
timestamp 1654752884
transform 1 0 8464 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_13
timestamp 1654752884
transform 1 0 22908 0 -1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_14
timestamp 1654752884
transform 1 0 7176 0 -1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_15
timestamp 1654752884
transform 1 0 18768 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_16
timestamp 1654752884
transform 1 0 8188 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_17
timestamp 1654752884
transform 1 0 6992 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_18
timestamp 1654752884
transform 1 0 22908 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_19
timestamp 1654752884
transform 1 0 19596 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_20
timestamp 1654752884
transform 1 0 18768 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_21
timestamp 1654752884
transform 1 0 18032 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_22
timestamp 1654752884
transform 1 0 22908 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_23
timestamp 1654752884
transform 1 0 20240 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_24
timestamp 1654752884
transform 1 0 9752 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_25
timestamp 1654752884
transform 1 0 8648 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_26
timestamp 1654752884
transform 1 0 22724 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_27
timestamp 1654752884
transform 1 0 18216 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_28
timestamp 1654752884
transform 1 0 8188 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_29
timestamp 1654752884
transform 1 0 5888 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_30
timestamp 1654752884
transform 1 0 22908 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_31
timestamp 1654752884
transform 1 0 21528 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_32
timestamp 1654752884
transform 1 0 22908 0 -1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_33
timestamp 1654752884
transform 1 0 17848 0 -1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_34
timestamp 1654752884
transform 1 0 12328 0 -1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_35
timestamp 1654752884
transform 1 0 13340 0 1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_36
timestamp 1654752884
transform 1 0 12512 0 1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_37
timestamp 1654752884
transform 1 0 22908 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_38
timestamp 1654752884
transform 1 0 7176 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_39
timestamp 1654752884
transform 1 0 16008 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_40
timestamp 1654752884
transform 1 0 14260 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_41
timestamp 1654752884
transform 1 0 9108 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_42
timestamp 1654752884
transform 1 0 8464 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_43
timestamp 1654752884
transform 1 0 7728 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_44
timestamp 1654752884
transform 1 0 22908 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_45
timestamp 1654752884
transform 1 0 19596 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_46
timestamp 1654752884
transform 1 0 18768 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_47
timestamp 1654752884
transform 1 0 15916 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_48
timestamp 1654752884
transform 1 0 15088 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_49
timestamp 1654752884
transform 1 0 10304 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_50
timestamp 1654752884
transform 1 0 22908 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_51
timestamp 1654752884
transform 1 0 16192 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_52
timestamp 1654752884
transform 1 0 8464 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_53
timestamp 1654752884
transform 1 0 22908 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_54
timestamp 1654752884
transform 1 0 17480 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_55
timestamp 1654752884
transform 1 0 9752 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_56
timestamp 1654752884
transform 1 0 9108 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_57
timestamp 1654752884
transform 1 0 8464 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_58
timestamp 1654752884
transform 1 0 22908 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_59
timestamp 1654752884
transform 1 0 15916 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_60
timestamp 1654752884
transform 1 0 15088 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_61
timestamp 1654752884
transform 1 0 11040 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_62
timestamp 1654752884
transform 1 0 9108 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_63
timestamp 1654752884
transform 1 0 8464 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_64
timestamp 1654752884
transform 1 0 22908 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_65
timestamp 1654752884
transform 1 0 21712 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_66
timestamp 1654752884
transform 1 0 16928 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_67
timestamp 1654752884
transform 1 0 9108 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_68
timestamp 1654752884
transform 1 0 8464 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_69
timestamp 1654752884
transform 1 0 14904 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_70
timestamp 1654752884
transform 1 0 12696 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_71
timestamp 1654752884
transform 1 0 9108 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_72
timestamp 1654752884
transform 1 0 8464 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_73
timestamp 1654752884
transform 1 0 22908 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_74
timestamp 1654752884
transform 1 0 9752 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_75
timestamp 1654752884
transform 1 0 22908 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_76
timestamp 1654752884
transform 1 0 18032 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_77
timestamp 1654752884
transform 1 0 14352 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_78
timestamp 1654752884
transform 1 0 11776 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_79
timestamp 1654752884
transform 1 0 8832 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_80
timestamp 1654752884
transform 1 0 5888 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_81
timestamp 1654752884
transform 1 0 22908 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_82
timestamp 1654752884
transform 1 0 22908 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_83
timestamp 1654752884
transform 1 0 22908 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_84
timestamp 1654752884
transform 1 0 21344 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_85
timestamp 1654752884
transform 1 0 18768 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_86
timestamp 1654752884
transform 1 0 18584 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_87
timestamp 1654752884
transform 1 0 18216 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_88
timestamp 1654752884
transform 1 0 13432 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_89
timestamp 1654752884
transform 1 0 12144 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_90
timestamp 1654752884
transform 1 0 6992 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_91
timestamp 1654752884
transform 1 0 18768 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_92
timestamp 1654752884
transform 1 0 17664 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_93
timestamp 1654752884
transform 1 0 16836 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_94
timestamp 1654752884
transform 1 0 13432 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_95
timestamp 1654752884
transform 1 0 8280 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_96
timestamp 1654752884
transform 1 0 7176 0 -1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_97
timestamp 1654752884
transform 1 0 21160 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_98
timestamp 1654752884
transform 1 0 18584 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_99
timestamp 1654752884
transform 1 0 16008 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_100
timestamp 1654752884
transform 1 0 13432 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_101
timestamp 1654752884
transform 1 0 8280 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_102
timestamp 1654752884
transform 1 0 17480 0 -1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_103
timestamp 1654752884
transform 1 0 9568 0 -1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_104
timestamp 1654752884
transform 1 0 8832 0 -1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_105
timestamp 1654752884
transform 1 0 22908 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_106
timestamp 1654752884
transform 1 0 21344 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_107
timestamp 1654752884
transform 1 0 14352 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_108
timestamp 1654752884
transform 1 0 8280 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_109
timestamp 1654752884
transform 1 0 6440 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_110
timestamp 1654752884
transform 1 0 12328 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_111
timestamp 1654752884
transform 1 0 12144 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_112
timestamp 1654752884
transform 1 0 9568 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_113
timestamp 1654752884
transform 1 0 19688 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_114
timestamp 1654752884
transform 1 0 6256 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_115
timestamp 1654752884
transform 1 0 10672 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_116
timestamp 1654752884
transform 1 0 6992 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_117
timestamp 1654752884
transform 1 0 5796 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_118
timestamp 1654752884
transform 1 0 21160 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_119
timestamp 1654752884
transform 1 0 20424 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_120
timestamp 1654752884
transform 1 0 16008 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_121
timestamp 1654752884
transform 1 0 13616 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_122
timestamp 1654752884
transform 1 0 8280 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_123
timestamp 1654752884
transform 1 0 22448 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_124
timestamp 1654752884
transform 1 0 17296 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_125
timestamp 1654752884
transform 1 0 16560 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_126
timestamp 1654752884
transform 1 0 12144 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_127
timestamp 1654752884
transform 1 0 10212 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_128
timestamp 1654752884
transform 1 0 21160 0 1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_129
timestamp 1654752884
transform 1 0 19596 0 1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_130
timestamp 1654752884
transform 1 0 11960 0 1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_131
timestamp 1654752884
transform 1 0 8924 0 1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_132
timestamp 1654752884
transform 1 0 17480 0 -1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_133
timestamp 1654752884
transform 1 0 10488 0 -1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_134
timestamp 1654752884
transform 1 0 18584 0 1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_135
timestamp 1654752884
transform 1 0 13432 0 1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_136
timestamp 1654752884
transform 1 0 10856 0 1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_137
timestamp 1654752884
transform 1 0 22448 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_138
timestamp 1654752884
transform 1 0 20056 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_139
timestamp 1654752884
transform 1 0 18952 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_140
timestamp 1654752884
transform 1 0 10672 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_141
timestamp 1654752884
transform 1 0 12788 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_142
timestamp 1654752884
transform 1 0 11040 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_143
timestamp 1654752884
transform 1 0 10856 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_144
timestamp 1654752884
transform 1 0 12696 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_145
timestamp 1654752884
transform 1 0 10488 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_146
timestamp 1654752884
transform 1 0 7176 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_147
timestamp 1654752884
transform 1 0 16008 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_148
timestamp 1654752884
transform 1 0 11776 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_149
timestamp 1654752884
transform 1 0 6256 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_150
timestamp 1654752884
transform 1 0 17480 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_151
timestamp 1654752884
transform 1 0 9752 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_152
timestamp 1654752884
transform 1 0 7176 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_153
timestamp 1654752884
transform 1 0 6532 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_154
timestamp 1654752884
transform 1 0 11960 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_155
timestamp 1654752884
transform 1 0 6532 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_156
timestamp 1654752884
transform 1 0 21528 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_157
timestamp 1654752884
transform 1 0 6716 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_158
timestamp 1654752884
transform 1 0 5796 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_159
timestamp 1654752884
transform 1 0 22908 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_160
timestamp 1654752884
transform 1 0 21344 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_161
timestamp 1654752884
transform 1 0 16008 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_162
timestamp 1654752884
transform 1 0 13432 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_163
timestamp 1654752884
transform 1 0 9200 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_164
timestamp 1654752884
transform 1 0 19872 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_165
timestamp 1654752884
transform 1 0 12512 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_166
timestamp 1654752884
transform 1 0 12144 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_167
timestamp 1654752884
transform 1 0 9200 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_168
timestamp 1654752884
transform 1 0 6808 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_169
timestamp 1654752884
transform 1 0 6256 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_170
timestamp 1654752884
transform 1 0 12144 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_171
timestamp 1654752884
transform 1 0 22816 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_172
timestamp 1654752884
transform 1 0 21160 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_173
timestamp 1654752884
transform 1 0 16008 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_174
timestamp 1654752884
transform 1 0 15088 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_175
timestamp 1654752884
transform 1 0 22448 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_176
timestamp 1654752884
transform 1 0 21344 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_177
timestamp 1654752884
transform 1 0 20056 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_178
timestamp 1654752884
transform 1 0 18768 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_179
timestamp 1654752884
transform 1 0 17480 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_180
timestamp 1654752884
transform 1 0 16192 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_181
timestamp 1654752884
transform 1 0 16008 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_182
timestamp 1654752884
transform 1 0 13616 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_183
timestamp 1654752884
transform 1 0 8280 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_184
timestamp 1654752884
transform 1 0 7728 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_185
timestamp 1654752884
transform 1 0 6992 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_0
timestamp 1654752884
transform 1 0 13616 0 -1 22032
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_1
timestamp 1654752884
transform 1 0 7176 0 -1 22032
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_2
timestamp 1654752884
transform 1 0 8464 0 1 20944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_3
timestamp 1654752884
transform 1 0 8740 0 -1 20944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_4
timestamp 1654752884
transform 1 0 5796 0 -1 20944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_5
timestamp 1654752884
transform 1 0 20240 0 1 19856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_6
timestamp 1654752884
transform 1 0 5888 0 1 19856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_7
timestamp 1654752884
transform 1 0 5796 0 -1 19856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_8
timestamp 1654752884
transform 1 0 8464 0 1 18768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_9
timestamp 1654752884
transform 1 0 9752 0 -1 18768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_10
timestamp 1654752884
transform 1 0 20056 0 -1 17680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_11
timestamp 1654752884
transform 1 0 16468 0 -1 17680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_12
timestamp 1654752884
transform 1 0 9752 0 -1 14416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_13
timestamp 1654752884
transform 1 0 8740 0 -1 13328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_14
timestamp 1654752884
transform 1 0 7176 0 1 12240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_15
timestamp 1654752884
transform 1 0 7176 0 1 10064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_16
timestamp 1654752884
transform 1 0 18676 0 -1 6800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_17
timestamp 1654752884
transform 1 0 15916 0 -1 22032
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_18
timestamp 1654752884
transform 1 0 15456 0 -1 22032
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_19
timestamp 1654752884
transform 1 0 14904 0 -1 22032
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_20
timestamp 1654752884
transform 1 0 17480 0 1 20944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_21
timestamp 1654752884
transform 1 0 16652 0 1 20944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_22
timestamp 1654752884
transform 1 0 14168 0 1 20944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_23
timestamp 1654752884
transform 1 0 13248 0 1 20944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_24
timestamp 1654752884
transform 1 0 15732 0 -1 20944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_25
timestamp 1654752884
transform 1 0 14628 0 -1 20944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_26
timestamp 1654752884
transform 1 0 14168 0 -1 20944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_27
timestamp 1654752884
transform 1 0 21344 0 1 19856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_28
timestamp 1654752884
transform 1 0 17204 0 -1 19856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_29
timestamp 1654752884
transform 1 0 14904 0 -1 19856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_30
timestamp 1654752884
transform 1 0 12052 0 -1 19856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_31
timestamp 1654752884
transform 1 0 9384 0 -1 19856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_32
timestamp 1654752884
transform 1 0 8648 0 -1 19856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_33
timestamp 1654752884
transform 1 0 11040 0 1 18768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_34
timestamp 1654752884
transform 1 0 6256 0 1 18768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_35
timestamp 1654752884
transform 1 0 22356 0 -1 18768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_36
timestamp 1654752884
transform 1 0 7176 0 -1 18768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_37
timestamp 1654752884
transform 1 0 5796 0 -1 18768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_38
timestamp 1654752884
transform 1 0 22816 0 1 17680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_39
timestamp 1654752884
transform 1 0 16192 0 1 17680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_40
timestamp 1654752884
transform 1 0 8188 0 1 17680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_41
timestamp 1654752884
transform 1 0 14904 0 -1 17680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_42
timestamp 1654752884
transform 1 0 9476 0 -1 17680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_43
timestamp 1654752884
transform 1 0 22816 0 1 16592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_44
timestamp 1654752884
transform 1 0 20240 0 1 16592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_45
timestamp 1654752884
transform 1 0 15824 0 1 16592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_46
timestamp 1654752884
transform 1 0 14904 0 -1 16592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_47
timestamp 1654752884
transform 1 0 13156 0 -1 16592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_48
timestamp 1654752884
transform 1 0 7176 0 -1 16592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_49
timestamp 1654752884
transform 1 0 5796 0 -1 16592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_50
timestamp 1654752884
transform 1 0 22816 0 1 15504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_51
timestamp 1654752884
transform 1 0 19412 0 1 15504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_52
timestamp 1654752884
transform 1 0 11500 0 1 15504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_53
timestamp 1654752884
transform 1 0 11040 0 1 15504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_54
timestamp 1654752884
transform 1 0 8740 0 1 15504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_55
timestamp 1654752884
transform 1 0 21896 0 -1 15504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_56
timestamp 1654752884
transform 1 0 9752 0 -1 15504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_57
timestamp 1654752884
transform 1 0 5796 0 -1 15504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_58
timestamp 1654752884
transform 1 0 22816 0 1 14416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_59
timestamp 1654752884
transform 1 0 15916 0 1 14416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_60
timestamp 1654752884
transform 1 0 22816 0 1 13328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_61
timestamp 1654752884
transform 1 0 13616 0 1 13328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_62
timestamp 1654752884
transform 1 0 13340 0 1 13328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_63
timestamp 1654752884
transform 1 0 15732 0 -1 13328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_64
timestamp 1654752884
transform 1 0 14904 0 -1 13328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_65
timestamp 1654752884
transform 1 0 22816 0 1 12240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_66
timestamp 1654752884
transform 1 0 13340 0 1 12240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_67
timestamp 1654752884
transform 1 0 8464 0 1 12240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_68
timestamp 1654752884
transform 1 0 6164 0 -1 12240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_69
timestamp 1654752884
transform 1 0 22816 0 1 11152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_70
timestamp 1654752884
transform 1 0 21068 0 1 11152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_71
timestamp 1654752884
transform 1 0 20240 0 1 11152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_72
timestamp 1654752884
transform 1 0 11868 0 1 11152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_73
timestamp 1654752884
transform 1 0 10764 0 1 11152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_74
timestamp 1654752884
transform 1 0 19780 0 -1 11152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_75
timestamp 1654752884
transform 1 0 12052 0 -1 11152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_76
timestamp 1654752884
transform 1 0 8740 0 -1 11152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_77
timestamp 1654752884
transform 1 0 22816 0 1 10064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_78
timestamp 1654752884
transform 1 0 11776 0 1 10064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_79
timestamp 1654752884
transform 1 0 19780 0 -1 10064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_80
timestamp 1654752884
transform 1 0 10396 0 -1 10064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_81
timestamp 1654752884
transform 1 0 9752 0 -1 10064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_82
timestamp 1654752884
transform 1 0 6164 0 -1 10064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_83
timestamp 1654752884
transform 1 0 10764 0 1 8976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_84
timestamp 1654752884
transform 1 0 12328 0 -1 8976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_85
timestamp 1654752884
transform 1 0 6900 0 -1 8976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_86
timestamp 1654752884
transform 1 0 22816 0 1 7888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_87
timestamp 1654752884
transform 1 0 13340 0 1 7888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_88
timestamp 1654752884
transform 1 0 10764 0 1 7888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_89
timestamp 1654752884
transform 1 0 22356 0 -1 7888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_90
timestamp 1654752884
transform 1 0 21712 0 -1 7888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_91
timestamp 1654752884
transform 1 0 8648 0 -1 7888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_92
timestamp 1654752884
transform 1 0 6900 0 -1 7888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_93
timestamp 1654752884
transform 1 0 17664 0 1 6800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_94
timestamp 1654752884
transform 1 0 6716 0 1 6800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_95
timestamp 1654752884
transform 1 0 21160 0 -1 6800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_96
timestamp 1654752884
transform 1 0 6348 0 -1 6800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_97
timestamp 1654752884
transform 1 0 5796 0 -1 6800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_98
timestamp 1654752884
transform 1 0 10764 0 1 5712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_99
timestamp 1654752884
transform 1 0 7544 0 1 5712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_0
timestamp 1654752884
transform 1 0 15364 0 -1 20944
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_1
timestamp 1654752884
transform 1 0 13800 0 -1 20944
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_2
timestamp 1654752884
transform 1 0 16836 0 -1 19856
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_3
timestamp 1654752884
transform 1 0 15548 0 -1 19856
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_4
timestamp 1654752884
transform 1 0 8280 0 -1 19856
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_5
timestamp 1654752884
transform 1 0 5888 0 1 18768
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_6
timestamp 1654752884
transform 1 0 21528 0 -1 18768
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_7
timestamp 1654752884
transform 1 0 7820 0 1 17680
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_8
timestamp 1654752884
transform 1 0 5888 0 1 17680
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_9
timestamp 1654752884
transform 1 0 21528 0 -1 15504
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_10
timestamp 1654752884
transform 1 0 20884 0 1 14416
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_11
timestamp 1654752884
transform 1 0 10488 0 1 14416
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_12
timestamp 1654752884
transform 1 0 8464 0 1 14416
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_13
timestamp 1654752884
transform 1 0 5888 0 1 13328
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_14
timestamp 1654752884
transform 1 0 16376 0 -1 12240
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_15
timestamp 1654752884
transform 1 0 5796 0 -1 12240
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_16
timestamp 1654752884
transform 1 0 20884 0 1 10064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_17
timestamp 1654752884
transform 1 0 18308 0 1 10064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_18
timestamp 1654752884
transform 1 0 19412 0 -1 10064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_19
timestamp 1654752884
transform 1 0 20884 0 1 8976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_20
timestamp 1654752884
transform 1 0 18308 0 1 8976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_21
timestamp 1654752884
transform 1 0 20884 0 1 7888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_22
timestamp 1654752884
transform 1 0 6072 0 -1 7888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_23
timestamp 1654752884
transform 1 0 18308 0 1 6800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_24
timestamp 1654752884
transform 1 0 15640 0 1 6800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_25
timestamp 1654752884
transform 1 0 7176 0 -1 6800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_26
timestamp 1654752884
transform 1 0 7176 0 1 5712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_0
timestamp 1654752884
transform 1 0 17480 0 -1 8976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_1
timestamp 1654752884
transform 1 0 9752 0 1 5712
box -38 -48 774 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_0
timestamp 1654752884
transform -1 0 7084 0 -1 15504
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_1
timestamp 1654752884
transform 1 0 5888 0 -1 17680
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_2
timestamp 1654752884
transform 1 0 5980 0 -1 18768
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_3
timestamp 1654752884
transform -1 0 8464 0 -1 18768
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_4
timestamp 1654752884
transform -1 0 9568 0 -1 18768
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_5
timestamp 1654752884
transform -1 0 10672 0 1 17680
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_6
timestamp 1654752884
transform -1 0 10488 0 1 18768
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_7
timestamp 1654752884
transform 1 0 20056 0 -1 6800
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_8
timestamp 1654752884
transform 1 0 18860 0 1 5712
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_9
timestamp 1654752884
transform -1 0 21252 0 1 5712
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_10
timestamp 1654752884
transform -1 0 22540 0 1 5712
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_11
timestamp 1654752884
transform -1 0 22448 0 -1 6800
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_12
timestamp 1654752884
transform 1 0 21436 0 1 8976
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_13
timestamp 1654752884
transform 1 0 18860 0 -1 18768
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_14
timestamp 1654752884
transform -1 0 22540 0 -1 22032
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_15
timestamp 1654752884
transform -1 0 17388 0 1 5712
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_0
timestamp 1654752884
transform -1 0 15364 0 1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_1
timestamp 1654752884
transform 1 0 13064 0 1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_2
timestamp 1654752884
transform 1 0 8464 0 1 15504
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_3
timestamp 1654752884
transform 1 0 11224 0 1 15504
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_4
timestamp 1654752884
transform -1 0 22908 0 -1 22032
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_5
timestamp 1654752884
transform 1 0 17756 0 1 20944
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_6
timestamp 1654752884
transform -1 0 14628 0 -1 20944
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_7
timestamp 1654752884
transform -1 0 6072 0 -1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_8
timestamp 1654752884
transform -1 0 6808 0 -1 13328
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_9
timestamp 1654752884
transform -1 0 6532 0 1 10064
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_10
timestamp 1654752884
transform 1 0 7176 0 -1 8976
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  sky130_fd_sc_hd__nand3_1_0
timestamp 1654752884
transform -1 0 9476 0 -1 17680
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  sky130_fd_sc_hd__nand3_1_1
timestamp 1654752884
transform -1 0 12144 0 -1 16592
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  sky130_fd_sc_hd__nand3_1_2
timestamp 1654752884
transform -1 0 6348 0 -1 6800
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_1  sky130_fd_sc_hd__nand4_1_0
timestamp 1654752884
transform 1 0 8924 0 -1 19856
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_0
timestamp 1654752884
transform -1 0 13524 0 1 5712
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_1
timestamp 1654752884
transform 1 0 13708 0 1 5712
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_2
timestamp 1654752884
transform -1 0 18584 0 -1 22032
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_3
timestamp 1654752884
transform 1 0 15640 0 -1 22032
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_4
timestamp 1654752884
transform 1 0 11592 0 1 18768
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_5
timestamp 1654752884
transform -1 0 6624 0 1 12240
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_6
timestamp 1654752884
transform -1 0 6164 0 -1 10064
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_7
timestamp 1654752884
transform 1 0 7912 0 -1 6800
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  sky130_fd_sc_hd__nor3_1_0
timestamp 1654752884
transform -1 0 9200 0 -1 16592
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  sky130_fd_sc_hd__o21a_1_0
timestamp 1654752884
transform 1 0 20056 0 -1 22032
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  sky130_fd_sc_hd__o21a_1_1
timestamp 1654752884
transform 1 0 16928 0 1 20944
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  sky130_fd_sc_hd__o21a_1_2
timestamp 1654752884
transform 1 0 13616 0 1 20944
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  sky130_fd_sc_hd__o21a_1_3
timestamp 1654752884
transform 1 0 11316 0 1 16592
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  sky130_fd_sc_hd__o21a_1_4
timestamp 1654752884
transform 1 0 9936 0 -1 15504
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  sky130_fd_sc_hd__o21a_1_5
timestamp 1654752884
transform -1 0 7268 0 1 13328
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  sky130_fd_sc_hd__o21a_1_6
timestamp 1654752884
transform 1 0 6624 0 1 10064
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  sky130_fd_sc_hd__o21a_1_7
timestamp 1654752884
transform 1 0 6348 0 -1 8976
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  sky130_fd_sc_hd__o21a_1_8
timestamp 1654752884
transform 1 0 6532 0 -1 6800
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  sky130_fd_sc_hd__o21a_1_9
timestamp 1654752884
transform -1 0 6440 0 1 6800
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  sky130_fd_sc_hd__o21ai_1_0
timestamp 1654752884
transform 1 0 14076 0 -1 7888
box -38 -48 406 592
use sky130_fd_sc_hd__sdlclkp_4  sky130_fd_sc_hd__sdlclkp_4_0
timestamp 1654752884
transform -1 0 16836 0 -1 14416
box -38 -48 1694 592
use sky130_fd_sc_hd__sdlclkp_4  sky130_fd_sc_hd__sdlclkp_4_1
timestamp 1654752884
transform 1 0 16468 0 1 15504
box -38 -48 1694 592
use sky130_fd_sc_hd__sdlclkp_4  sky130_fd_sc_hd__sdlclkp_4_2
timestamp 1654752884
transform -1 0 19872 0 -1 8976
box -38 -48 1694 592
use sky130_fd_sc_hd__sdlclkp_4  sky130_fd_sc_hd__sdlclkp_4_3
timestamp 1654752884
transform -1 0 17388 0 -1 7888
box -38 -48 1694 592
use sky130_fd_sc_hd__sdlclkp_4  sky130_fd_sc_hd__sdlclkp_4_4
timestamp 1654752884
transform 1 0 13156 0 -1 15504
box -38 -48 1694 592
use sky130_fd_sc_hd__sdlclkp_4  sky130_fd_sc_hd__sdlclkp_4_5
timestamp 1654752884
transform -1 0 19412 0 -1 10064
box -38 -48 1694 592
use sky130_fd_sc_hd__sdlclkp_4  sky130_fd_sc_hd__sdlclkp_4_6
timestamp 1654752884
transform 1 0 16376 0 1 17680
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1654752884
transform 1 0 22540 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1654752884
transform 1 0 21252 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1654752884
transform 1 0 19964 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1654752884
transform 1 0 18676 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1654752884
transform 1 0 17388 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1654752884
transform 1 0 16100 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1654752884
transform 1 0 14812 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1654752884
transform 1 0 13524 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_8
timestamp 1654752884
transform 1 0 12236 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_9
timestamp 1654752884
transform 1 0 10948 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_10
timestamp 1654752884
transform 1 0 9660 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_11
timestamp 1654752884
transform 1 0 8372 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_12
timestamp 1654752884
transform 1 0 7084 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_13
timestamp 1654752884
transform 1 0 5796 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_14
timestamp 1654752884
transform 1 0 21252 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_15
timestamp 1654752884
transform 1 0 18676 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_16
timestamp 1654752884
transform 1 0 16100 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_17
timestamp 1654752884
transform 1 0 13524 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_18
timestamp 1654752884
transform 1 0 10948 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_19
timestamp 1654752884
transform 1 0 8372 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_20
timestamp 1654752884
transform 1 0 5796 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_21
timestamp 1654752884
transform 1 0 22540 0 -1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_22
timestamp 1654752884
transform 1 0 19964 0 -1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_23
timestamp 1654752884
transform 1 0 17388 0 -1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_24
timestamp 1654752884
transform 1 0 14812 0 -1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_25
timestamp 1654752884
transform 1 0 12236 0 -1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_26
timestamp 1654752884
transform 1 0 9660 0 -1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_27
timestamp 1654752884
transform 1 0 7084 0 -1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_28
timestamp 1654752884
transform 1 0 21252 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_29
timestamp 1654752884
transform 1 0 18676 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_30
timestamp 1654752884
transform 1 0 16100 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_31
timestamp 1654752884
transform 1 0 13524 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_32
timestamp 1654752884
transform 1 0 10948 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_33
timestamp 1654752884
transform 1 0 8372 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_34
timestamp 1654752884
transform 1 0 5796 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_35
timestamp 1654752884
transform 1 0 22540 0 -1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_36
timestamp 1654752884
transform 1 0 19964 0 -1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_37
timestamp 1654752884
transform 1 0 17388 0 -1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_38
timestamp 1654752884
transform 1 0 14812 0 -1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_39
timestamp 1654752884
transform 1 0 12236 0 -1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_40
timestamp 1654752884
transform 1 0 9660 0 -1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_41
timestamp 1654752884
transform 1 0 7084 0 -1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_42
timestamp 1654752884
transform 1 0 21252 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_43
timestamp 1654752884
transform 1 0 18676 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_44
timestamp 1654752884
transform 1 0 16100 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_45
timestamp 1654752884
transform 1 0 13524 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_46
timestamp 1654752884
transform 1 0 10948 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_47
timestamp 1654752884
transform 1 0 8372 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_48
timestamp 1654752884
transform 1 0 5796 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_49
timestamp 1654752884
transform 1 0 22540 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_50
timestamp 1654752884
transform 1 0 19964 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_51
timestamp 1654752884
transform 1 0 17388 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_52
timestamp 1654752884
transform 1 0 14812 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_53
timestamp 1654752884
transform 1 0 12236 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_54
timestamp 1654752884
transform 1 0 9660 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_55
timestamp 1654752884
transform 1 0 7084 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_56
timestamp 1654752884
transform 1 0 21252 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_57
timestamp 1654752884
transform 1 0 18676 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_58
timestamp 1654752884
transform 1 0 16100 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_59
timestamp 1654752884
transform 1 0 13524 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_60
timestamp 1654752884
transform 1 0 10948 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_61
timestamp 1654752884
transform 1 0 8372 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_62
timestamp 1654752884
transform 1 0 5796 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_63
timestamp 1654752884
transform 1 0 22540 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_64
timestamp 1654752884
transform 1 0 19964 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_65
timestamp 1654752884
transform 1 0 17388 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_66
timestamp 1654752884
transform 1 0 14812 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_67
timestamp 1654752884
transform 1 0 12236 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_68
timestamp 1654752884
transform 1 0 9660 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_69
timestamp 1654752884
transform 1 0 7084 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_70
timestamp 1654752884
transform 1 0 21252 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_71
timestamp 1654752884
transform 1 0 18676 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_72
timestamp 1654752884
transform 1 0 16100 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_73
timestamp 1654752884
transform 1 0 13524 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_74
timestamp 1654752884
transform 1 0 10948 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_75
timestamp 1654752884
transform 1 0 8372 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_76
timestamp 1654752884
transform 1 0 5796 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_77
timestamp 1654752884
transform 1 0 22540 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_78
timestamp 1654752884
transform 1 0 19964 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_79
timestamp 1654752884
transform 1 0 17388 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_80
timestamp 1654752884
transform 1 0 14812 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_81
timestamp 1654752884
transform 1 0 12236 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_82
timestamp 1654752884
transform 1 0 9660 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_83
timestamp 1654752884
transform 1 0 7084 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_84
timestamp 1654752884
transform 1 0 21252 0 1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_85
timestamp 1654752884
transform 1 0 18676 0 1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_86
timestamp 1654752884
transform 1 0 16100 0 1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_87
timestamp 1654752884
transform 1 0 13524 0 1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_88
timestamp 1654752884
transform 1 0 10948 0 1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_89
timestamp 1654752884
transform 1 0 8372 0 1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_90
timestamp 1654752884
transform 1 0 5796 0 1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_91
timestamp 1654752884
transform 1 0 22540 0 -1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_92
timestamp 1654752884
transform 1 0 19964 0 -1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_93
timestamp 1654752884
transform 1 0 17388 0 -1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_94
timestamp 1654752884
transform 1 0 14812 0 -1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_95
timestamp 1654752884
transform 1 0 12236 0 -1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_96
timestamp 1654752884
transform 1 0 9660 0 -1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_97
timestamp 1654752884
transform 1 0 7084 0 -1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_98
timestamp 1654752884
transform 1 0 21252 0 1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_99
timestamp 1654752884
transform 1 0 18676 0 1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_100
timestamp 1654752884
transform 1 0 16100 0 1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_101
timestamp 1654752884
transform 1 0 13524 0 1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_102
timestamp 1654752884
transform 1 0 10948 0 1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_103
timestamp 1654752884
transform 1 0 8372 0 1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_104
timestamp 1654752884
transform 1 0 5796 0 1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_105
timestamp 1654752884
transform 1 0 22540 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_106
timestamp 1654752884
transform 1 0 19964 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_107
timestamp 1654752884
transform 1 0 17388 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_108
timestamp 1654752884
transform 1 0 14812 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_109
timestamp 1654752884
transform 1 0 12236 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_110
timestamp 1654752884
transform 1 0 9660 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_111
timestamp 1654752884
transform 1 0 7084 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_112
timestamp 1654752884
transform 1 0 21252 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_113
timestamp 1654752884
transform 1 0 18676 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_114
timestamp 1654752884
transform 1 0 16100 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_115
timestamp 1654752884
transform 1 0 13524 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_116
timestamp 1654752884
transform 1 0 10948 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_117
timestamp 1654752884
transform 1 0 8372 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_118
timestamp 1654752884
transform 1 0 5796 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_119
timestamp 1654752884
transform 1 0 22540 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_120
timestamp 1654752884
transform 1 0 19964 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_121
timestamp 1654752884
transform 1 0 17388 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_122
timestamp 1654752884
transform 1 0 14812 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_123
timestamp 1654752884
transform 1 0 12236 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_124
timestamp 1654752884
transform 1 0 9660 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_125
timestamp 1654752884
transform 1 0 7084 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_126
timestamp 1654752884
transform 1 0 21252 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_127
timestamp 1654752884
transform 1 0 18676 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_128
timestamp 1654752884
transform 1 0 16100 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_129
timestamp 1654752884
transform 1 0 13524 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_130
timestamp 1654752884
transform 1 0 10948 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_131
timestamp 1654752884
transform 1 0 8372 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_132
timestamp 1654752884
transform 1 0 5796 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_133
timestamp 1654752884
transform 1 0 22540 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_134
timestamp 1654752884
transform 1 0 19964 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_135
timestamp 1654752884
transform 1 0 17388 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_136
timestamp 1654752884
transform 1 0 14812 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_137
timestamp 1654752884
transform 1 0 12236 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_138
timestamp 1654752884
transform 1 0 9660 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_139
timestamp 1654752884
transform 1 0 7084 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_140
timestamp 1654752884
transform 1 0 21252 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_141
timestamp 1654752884
transform 1 0 18676 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_142
timestamp 1654752884
transform 1 0 16100 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_143
timestamp 1654752884
transform 1 0 13524 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_144
timestamp 1654752884
transform 1 0 10948 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_145
timestamp 1654752884
transform 1 0 8372 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_146
timestamp 1654752884
transform 1 0 5796 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_147
timestamp 1654752884
transform 1 0 22540 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_148
timestamp 1654752884
transform 1 0 19964 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_149
timestamp 1654752884
transform 1 0 17388 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_150
timestamp 1654752884
transform 1 0 14812 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_151
timestamp 1654752884
transform 1 0 12236 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_152
timestamp 1654752884
transform 1 0 9660 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_153
timestamp 1654752884
transform 1 0 7084 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_154
timestamp 1654752884
transform 1 0 21252 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_155
timestamp 1654752884
transform 1 0 18676 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_156
timestamp 1654752884
transform 1 0 16100 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_157
timestamp 1654752884
transform 1 0 13524 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_158
timestamp 1654752884
transform 1 0 10948 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_159
timestamp 1654752884
transform 1 0 8372 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_160
timestamp 1654752884
transform 1 0 5796 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_161
timestamp 1654752884
transform 1 0 22540 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_162
timestamp 1654752884
transform 1 0 19964 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_163
timestamp 1654752884
transform 1 0 17388 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_164
timestamp 1654752884
transform 1 0 14812 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_165
timestamp 1654752884
transform 1 0 12236 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_166
timestamp 1654752884
transform 1 0 9660 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_167
timestamp 1654752884
transform 1 0 7084 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_168
timestamp 1654752884
transform 1 0 21252 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_169
timestamp 1654752884
transform 1 0 18676 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_170
timestamp 1654752884
transform 1 0 16100 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_171
timestamp 1654752884
transform 1 0 13524 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_172
timestamp 1654752884
transform 1 0 10948 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_173
timestamp 1654752884
transform 1 0 8372 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_174
timestamp 1654752884
transform 1 0 5796 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_175
timestamp 1654752884
transform 1 0 22540 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_176
timestamp 1654752884
transform 1 0 19964 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_177
timestamp 1654752884
transform 1 0 17388 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_178
timestamp 1654752884
transform 1 0 14812 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_179
timestamp 1654752884
transform 1 0 12236 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_180
timestamp 1654752884
transform 1 0 9660 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_181
timestamp 1654752884
transform 1 0 7084 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_182
timestamp 1654752884
transform 1 0 21252 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_183
timestamp 1654752884
transform 1 0 18676 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_184
timestamp 1654752884
transform 1 0 16100 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_185
timestamp 1654752884
transform 1 0 13524 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_186
timestamp 1654752884
transform 1 0 10948 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_187
timestamp 1654752884
transform 1 0 8372 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_188
timestamp 1654752884
transform 1 0 5796 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_189
timestamp 1654752884
transform 1 0 22540 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_190
timestamp 1654752884
transform 1 0 19964 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_191
timestamp 1654752884
transform 1 0 17388 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_192
timestamp 1654752884
transform 1 0 14812 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_193
timestamp 1654752884
transform 1 0 12236 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_194
timestamp 1654752884
transform 1 0 9660 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_195
timestamp 1654752884
transform 1 0 7084 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_196
timestamp 1654752884
transform 1 0 21252 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_197
timestamp 1654752884
transform 1 0 18676 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_198
timestamp 1654752884
transform 1 0 16100 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_199
timestamp 1654752884
transform 1 0 13524 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_200
timestamp 1654752884
transform 1 0 10948 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_201
timestamp 1654752884
transform 1 0 8372 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_202
timestamp 1654752884
transform 1 0 5796 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_203
timestamp 1654752884
transform 1 0 22540 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_204
timestamp 1654752884
transform 1 0 19964 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_205
timestamp 1654752884
transform 1 0 17388 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_206
timestamp 1654752884
transform 1 0 14812 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_207
timestamp 1654752884
transform 1 0 12236 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_208
timestamp 1654752884
transform 1 0 9660 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_209
timestamp 1654752884
transform 1 0 7084 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_210
timestamp 1654752884
transform 1 0 22540 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_211
timestamp 1654752884
transform 1 0 21252 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_212
timestamp 1654752884
transform 1 0 19964 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_213
timestamp 1654752884
transform 1 0 18676 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_214
timestamp 1654752884
transform 1 0 17388 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_215
timestamp 1654752884
transform 1 0 16100 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_216
timestamp 1654752884
transform 1 0 14812 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_217
timestamp 1654752884
transform 1 0 13524 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_218
timestamp 1654752884
transform 1 0 12236 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_219
timestamp 1654752884
transform 1 0 10948 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_220
timestamp 1654752884
transform 1 0 9660 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_221
timestamp 1654752884
transform 1 0 8372 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_222
timestamp 1654752884
transform 1 0 7084 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_223
timestamp 1654752884
transform 1 0 5796 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__xnor2_1  sky130_fd_sc_hd__xnor2_1_0
timestamp 1654752884
transform -1 0 21252 0 -1 22032
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  sky130_fd_sc_hd__xnor2_1_1
timestamp 1654752884
transform -1 0 6808 0 -1 14416
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_0
timestamp 1654752884
transform 1 0 5980 0 -1 16592
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_1
timestamp 1654752884
transform 1 0 21896 0 -1 11152
box -38 -48 682 592
<< labels >>
rlabel metal2 s 28736 0 28764 97 4 clk
port 1 nsew
rlabel metal2 s 19168 0 19196 97 4 rst_n
port 2 nsew
rlabel metal2 s 9600 0 9628 97 4 sclk
port 3 nsew
rlabel metal2 s 32 0 60 97 4 cs_n
port 4 nsew
rlabel metal3 s 0 13768 160 13828 4 data_in
port 5 nsew
rlabel metal3 s 28636 104 28796 164 4 data_out[11]
port 6 nsew
rlabel metal3 s 28636 2666 28796 2726 4 data_out[10]
port 7 nsew
rlabel metal3 s 28636 5228 28796 5288 4 data_out[9]
port 8 nsew
rlabel metal3 s 28636 7668 28796 7728 4 data_out[8]
port 9 nsew
rlabel metal3 s 28636 10230 28796 10290 4 data_out[7]
port 10 nsew
rlabel metal3 s 28636 12670 28796 12730 4 data_out[6]
port 11 nsew
rlabel metal3 s 28636 15232 28796 15292 4 data_out[5]
port 12 nsew
rlabel metal3 s 28636 17672 28796 17732 4 data_out[4]
port 13 nsew
rlabel metal3 s 28636 20234 28796 20294 4 data_out[3]
port 14 nsew
rlabel metal3 s 28636 22674 28796 22734 4 data_out[2]
port 15 nsew
rlabel metal3 s 28636 25236 28796 25296 4 data_out[1]
port 16 nsew
rlabel metal3 s 28636 27676 28796 27736 4 data_out[0]
port 17 nsew
rlabel metal2 s 32 27647 60 27744 4 new_data
port 18 nsew
rlabel metal2 s 28736 27647 28764 27744 4 serial_data_out
port 19 nsew
rlabel metal5 s 0 3852 620 4472 4 VSS
port 20 nsew
rlabel metal5 s 0 5092 620 5712 4 VDD
port 21 nsew
<< properties >>
string path 451.950 281.350 456.550 281.350 
<< end >>
