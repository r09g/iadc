magic
tech sky130A
magscale 1 2
timestamp 1654720150
<< locali >>
rect -6 1174 1554 1238
rect -6 -86 58 1174
rect 214 1056 278 1174
rect 1344 1048 1408 1174
rect 1390 44 1554 108
rect -6 -150 210 -86
rect 210 -1210 274 -1100
rect 1340 -1210 1404 -1090
rect 1490 -1210 1554 44
rect -6 -1274 1554 -1210
<< viali >>
rect 697 942 731 976
rect 889 942 923 976
rect 313 131 347 165
rect 505 131 539 165
rect 307 -210 341 -176
rect 499 -210 533 -176
rect 691 -1021 725 -987
rect 883 -1021 917 -987
<< metal1 >>
rect 163 36 197 1078
rect 678 934 688 986
rect 740 934 750 986
rect 872 934 882 986
rect 934 934 944 986
rect 1444 496 1508 498
rect 1292 432 1508 496
rect 294 122 304 174
rect 356 122 366 174
rect 488 122 498 174
rect 550 122 560 174
rect 157 -1116 191 -74
rect 288 -218 298 -166
rect 350 -218 360 -166
rect 480 -220 490 -168
rect 542 -220 552 -168
rect 1444 -656 1508 432
rect 1280 -720 1508 -656
rect 672 -1030 682 -978
rect 734 -1030 744 -978
rect 864 -1030 874 -978
rect 926 -1030 936 -978
<< via1 >>
rect 688 976 740 986
rect 688 942 697 976
rect 697 942 731 976
rect 731 942 740 976
rect 688 934 740 942
rect 882 976 934 986
rect 882 942 889 976
rect 889 942 923 976
rect 923 942 934 976
rect 882 934 934 942
rect 304 165 356 174
rect 304 131 313 165
rect 313 131 347 165
rect 347 131 356 165
rect 304 122 356 131
rect 498 165 550 174
rect 498 131 505 165
rect 505 131 539 165
rect 539 131 550 165
rect 498 122 550 131
rect 298 -176 350 -166
rect 298 -210 307 -176
rect 307 -210 341 -176
rect 341 -210 350 -176
rect 298 -218 350 -210
rect 490 -176 542 -168
rect 490 -210 499 -176
rect 499 -210 533 -176
rect 533 -210 542 -176
rect 490 -220 542 -210
rect 682 -987 734 -978
rect 682 -1021 691 -987
rect 691 -1021 725 -987
rect 725 -1021 734 -987
rect 682 -1030 734 -1021
rect 874 -987 926 -978
rect 874 -1021 883 -987
rect 883 -1021 917 -987
rect 917 -1021 926 -987
rect 874 -1030 926 -1021
<< metal2 >>
rect 688 994 740 996
rect 682 986 740 994
rect 682 934 688 986
rect 882 986 934 996
rect 682 924 740 934
rect 874 934 882 980
rect 874 924 934 934
rect 682 508 734 924
rect 874 508 926 924
rect 682 456 926 508
rect 682 382 734 456
rect 102 330 734 382
rect 304 174 356 184
rect 498 174 550 184
rect 304 6 356 122
rect 490 122 498 174
rect 490 112 550 122
rect 490 6 542 112
rect 304 -46 542 6
rect 304 -156 356 -46
rect 298 -162 356 -156
rect 100 -166 356 -162
rect 100 -214 298 -166
rect 350 -218 356 -166
rect 490 -168 542 -46
rect 298 -228 350 -218
rect 490 -230 542 -220
rect 682 -654 734 330
rect 874 -654 926 456
rect 682 -706 926 -654
rect 682 -978 734 -706
rect 682 -1040 734 -1030
rect 874 -978 926 -706
rect 874 -1040 926 -1030
use transmission_gate  transmission_gate_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout_v2/transmission_gate
timestamp 1654720150
transform 1 0 216 0 1 51
box -53 -49 1241 1063
use transmission_gate  transmission_gate_1
timestamp 1654720150
transform 1 0 210 0 1 -1101
box -53 -49 1241 1063
<< labels >>
flabel metal1 178 412 178 412 1 FreeSans 400 0 0 0 v_hi
port 1 n
flabel metal1 174 -724 174 -724 1 FreeSans 400 0 0 0 v_lo
port 2 n
flabel metal2 120 354 120 354 1 FreeSans 400 0 0 0 v_b
port 4 n
flabel metal2 114 -188 114 -188 1 FreeSans 400 0 0 0 v
port 3 n
flabel metal1 1480 -6 1480 -6 1 FreeSans 400 0 0 0 out
port 5 n
flabel locali 32 1202 32 1202 1 FreeSans 400 0 0 0 VDD
port 6 n power bidirectional
flabel locali 14 -1244 14 -1244 1 FreeSans 400 0 0 0 VSS
port 7 n ground bidirectional
<< end >>
