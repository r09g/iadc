* NGSPICE file created from sc_cmfb_flat.ext - technology: sky130A

.subckt sc_cmfb_flat on cm bias_a op cmc p2_b p2 p1_b p1 VDD VSS
X0 cm p2 transmission_gate_3/out VSS sky130_fd_pr__nfet_01v8 ad=3.498e+12p pd=3.44e+07u as=1.9027e+12p ps=1.884e+07u w=530000u l=150000u
X1 transmission_gate_6/in p2_b op VDD sky130_fd_pr__pfet_01v8 ad=4.9183e+12p pd=3.732e+07u as=5.3156e+12p ps=4.064e+07u w=1.37e+06u l=150000u
X2 transmission_gate_8/in p2 cmc VSS sky130_fd_pr__nfet_01v8 ad=1.9027e+12p pd=1.884e+07u as=2.0564e+12p ps=2.048e+07u w=530000u l=150000u
X3 transmission_gate_7/in p1_b cm VDD sky130_fd_pr__pfet_01v8 ad=4.9183e+12p pd=3.732e+07u as=9.042e+12p ps=6.8e+07u w=1.37e+06u l=150000u
X4 op p2 transmission_gate_6/in VSS sky130_fd_pr__nfet_01v8 ad=2.0564e+12p pd=2.048e+07u as=1.9027e+12p ps=1.884e+07u w=530000u l=150000u
X5 transmission_gate_5/out p2 bias_a VSS sky130_fd_pr__nfet_01v8 ad=1.9027e+12p pd=1.884e+07u as=1.749e+12p ps=1.72e+07u w=530000u l=150000u
X6 cm p1_b transmission_gate_7/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X7 transmission_gate_7/in p1_b cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X8 cm p1_b transmission_gate_7/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X9 on cmc sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X10 transmission_gate_5/out p2_b bias_a VDD sky130_fd_pr__pfet_01v8 ad=4.9183e+12p pd=3.732e+07u as=4.521e+12p ps=3.4e+07u w=1.37e+06u l=150000u
X11 cmc p1_b transmission_gate_5/out VDD sky130_fd_pr__pfet_01v8 ad=5.3156e+12p pd=4.064e+07u as=0p ps=0u w=1.37e+06u l=150000u
X12 cmc p1 transmission_gate_5/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X13 c1_n1700_n1700# m3_n1800_n1800# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X14 transmission_gate_6/in p1_b cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X15 transmission_gate_7/in p1_b cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X16 cm p1_b transmission_gate_7/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X17 transmission_gate_7/in p1_b cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X18 c1_7300_5500# m3_7200_5400# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X19 c1_3700_n1700# m3_3600_n1800# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X20 on cmc sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X21 cm p2_b transmission_gate_4/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.9183e+12p ps=3.732e+07u w=1.37e+06u l=150000u
X22 cm p1 transmission_gate_6/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X23 cm p1_b transmission_gate_7/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X24 transmission_gate_7/in p1_b cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X25 c1_1900_7300# m3_1800_7200# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X26 transmission_gate_7/in p2_b on VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.3156e+12p ps=4.064e+07u w=1.37e+06u l=150000u
X27 on p2 transmission_gate_7/in VSS sky130_fd_pr__nfet_01v8 ad=2.0564e+12p pd=2.048e+07u as=1.9027e+12p ps=1.884e+07u w=530000u l=150000u
X28 op cmc sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X29 bias_a p2 transmission_gate_5/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X30 cm p2 transmission_gate_4/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.9027e+12p ps=1.884e+07u w=530000u l=150000u
X31 cmc p2 transmission_gate_8/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X32 transmission_gate_6/in p2 op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X33 cm p1_b transmission_gate_6/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X34 transmission_gate_5/out p1_b cmc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X35 on p2_b transmission_gate_7/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X36 transmission_gate_3/out p1_b on VDD sky130_fd_pr__pfet_01v8 ad=4.9183e+12p pd=3.732e+07u as=0p ps=0u w=1.37e+06u l=150000u
X37 transmission_gate_4/out p2_b cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X38 cmc p1 transmission_gate_5/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X39 transmission_gate_6/in p1 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X40 transmission_gate_8/in p2 cmc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X41 cm p2 transmission_gate_3/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X42 bias_a p1 transmission_gate_8/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X43 bias_a p1_b transmission_gate_8/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.9183e+12p ps=3.732e+07u w=1.37e+06u l=150000u
X44 on p2 transmission_gate_7/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X45 op p2 transmission_gate_6/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X46 transmission_gate_4/out p2 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X47 c1_7300_1900# m3_7200_1800# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X48 c1_n1700_5500# m3_n1800_5400# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X49 cmc p2_b transmission_gate_8/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X50 transmission_gate_4/out transmission_gate_5/out sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X51 transmission_gate_8/in p1 bias_a VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X52 cm p2_b transmission_gate_4/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X53 cmc p1_b transmission_gate_5/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X54 c1_3700_7300# m3_3600_7200# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X55 transmission_gate_8/in p1_b bias_a VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X56 cm p2_b transmission_gate_3/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X57 transmission_gate_6/in transmission_gate_8/in sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X58 transmission_gate_7/in p2_b on VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X59 transmission_gate_5/out p1 cmc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X60 cm p1 transmission_gate_6/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X61 op p2_b transmission_gate_6/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X62 cmc p2 transmission_gate_8/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X63 transmission_gate_6/in p2 op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X64 transmission_gate_3/out p2 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X65 bias_a p2 transmission_gate_5/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X66 bias_a p2_b transmission_gate_5/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X67 transmission_gate_7/in p2 on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X68 cm p2 transmission_gate_4/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X69 transmission_gate_5/out p1_b cmc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X70 cm p1_b transmission_gate_6/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X71 cm p1_b transmission_gate_7/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X72 transmission_gate_8/in p1 bias_a VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X73 transmission_gate_6/in p1 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X74 transmission_gate_8/in p1_b bias_a VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X75 cmc p2_b transmission_gate_8/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X76 transmission_gate_4/out p1 op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X77 on p2_b transmission_gate_7/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X78 transmission_gate_3/out p2_b cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X79 transmission_gate_4/out p1_b op VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X80 transmission_gate_8/in p2 cmc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X81 op p1 transmission_gate_4/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X82 op p2_b transmission_gate_6/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X83 op p2 transmission_gate_6/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X84 transmission_gate_4/out p2 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X85 c1_n1700_1900# m3_n1800_1800# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X86 op p1_b transmission_gate_4/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X87 transmission_gate_5/out p2_b bias_a VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X88 transmission_gate_5/out p2 bias_a VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X89 transmission_gate_3/out p2 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X90 c1_5500_7300# m3_5400_7200# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X91 cmc p1_b transmission_gate_5/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X92 transmission_gate_3/out transmission_gate_5/out sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X93 transmission_gate_7/in p2_b on VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X94 transmission_gate_6/in p1_b cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X95 transmission_gate_3/out p1_b on VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X96 on p1_b transmission_gate_3/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X97 cm p2_b transmission_gate_4/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X98 transmission_gate_8/in p2_b cmc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X99 cm p1 transmission_gate_6/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X100 on p1_b transmission_gate_3/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X101 transmission_gate_3/out p1_b on VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X102 on p1_b transmission_gate_3/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X103 cm p2_b transmission_gate_3/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X104 transmission_gate_5/out p1 cmc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X105 transmission_gate_3/out p1_b on VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X106 transmission_gate_3/out p1_b on VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X107 on p1_b transmission_gate_3/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X108 on p1_b transmission_gate_3/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X109 transmission_gate_7/in transmission_gate_8/in sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X110 op p1 transmission_gate_4/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X111 transmission_gate_6/in p2 op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X112 cm p2 transmission_gate_4/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X113 op p1_b transmission_gate_4/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X114 transmission_gate_6/in p2_b op VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X115 transmission_gate_7/in p2 on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X116 transmission_gate_7/in p1 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X117 bias_a p2_b transmission_gate_5/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X118 transmission_gate_5/out p2 bias_a VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X119 transmission_gate_3/out p2_b cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X120 transmission_gate_5/out p1_b cmc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X121 transmission_gate_4/out p1 op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X122 cm p1 transmission_gate_7/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X123 transmission_gate_7/in p1 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X124 cm p1 transmission_gate_7/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X125 on p2_b transmission_gate_7/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X126 cmc p1 transmission_gate_5/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X127 transmission_gate_4/out p1_b op VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X128 cm p1 transmission_gate_7/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X129 transmission_gate_7/in p1 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X130 transmission_gate_4/out p2_b cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X131 transmission_gate_6/in p1_b cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X132 transmission_gate_6/in p1 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X133 transmission_gate_7/in p1 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X134 transmission_gate_7/in p1 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X135 cm p1 transmission_gate_7/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X136 transmission_gate_7/in transmission_gate_8/in sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X137 transmission_gate_5/out p2_b bias_a VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X138 on p2 transmission_gate_7/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X139 c1_7300_7300# m3_7200_7200# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X140 transmission_gate_4/out p2 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X141 op cmc sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X142 transmission_gate_4/out p1 op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X143 cm p1 transmission_gate_6/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X144 c1_5500_n1700# m3_5400_n1800# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X145 transmission_gate_4/out p1_b op VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X146 transmission_gate_7/in p2_b on VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X147 cm p2_b transmission_gate_3/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X148 c1_n1700_100# m3_n1800_0# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X149 transmission_gate_8/in p2_b cmc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X150 transmission_gate_5/out p1 cmc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X151 op p1 transmission_gate_4/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X152 transmission_gate_3/out p1 on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X153 transmission_gate_4/out p2_b cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X154 cmc p2 transmission_gate_8/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X155 op p1_b transmission_gate_4/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X156 bias_a p2_b transmission_gate_5/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X157 cm p2 transmission_gate_4/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X158 transmission_gate_4/out p1 op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X159 transmission_gate_7/in p2 on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X160 cm p2 transmission_gate_3/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X161 transmission_gate_4/out p1_b op VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X162 transmission_gate_6/in p2_b op VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X163 bias_a p1 transmission_gate_8/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X164 cmc p2_b transmission_gate_8/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X165 bias_a p1_b transmission_gate_8/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X166 transmission_gate_3/out p2_b cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X167 transmission_gate_8/in p1 bias_a VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X168 cmc p1 transmission_gate_5/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X169 c1_1900_n1700# m3_1800_n1800# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X170 transmission_gate_8/in p1_b bias_a VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X171 op cmc sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X172 c1_7300_3700# m3_7200_3600# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X173 c1_n1700_7300# m3_n1800_7200# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X174 bias_a p1 transmission_gate_8/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X175 op p2_b transmission_gate_6/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X176 op p2 transmission_gate_6/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X177 cmc p2 transmission_gate_8/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X178 op cmc sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X179 bias_a p1_b transmission_gate_8/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X180 transmission_gate_5/out p2_b bias_a VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X181 on p2 transmission_gate_7/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X182 transmission_gate_3/out p2 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X183 bias_a p2 transmission_gate_5/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X184 cmc p1_b transmission_gate_5/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X185 transmission_gate_5/out p1 cmc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X186 cm p2_b transmission_gate_3/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X187 cm p1_b transmission_gate_6/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X188 cm p1 transmission_gate_6/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X189 transmission_gate_8/in p2_b cmc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X190 cm p1 transmission_gate_7/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X191 bias_a p2_b transmission_gate_5/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X192 transmission_gate_7/in p2 on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X193 c1_7300_100# m3_7200_0# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X194 bias_a p1 transmission_gate_8/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X195 transmission_gate_6/in p2_b op VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X196 cm p2 transmission_gate_4/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X197 transmission_gate_8/in p2 cmc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X198 bias_a p1_b transmission_gate_8/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X199 cm p2 transmission_gate_3/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X200 op p2 transmission_gate_6/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X201 transmission_gate_5/out p2 bias_a VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X202 on p2_b transmission_gate_7/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X203 transmission_gate_8/in p1 bias_a VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X204 cmc p1_b transmission_gate_5/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X205 cmc p1 transmission_gate_5/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X206 transmission_gate_8/in p1_b bias_a VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X207 on p1 transmission_gate_3/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X208 cmc p2_b transmission_gate_8/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X209 transmission_gate_6/in p1_b cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X210 transmission_gate_6/in p1 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X211 transmission_gate_3/out p1 on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X212 cm p2_b transmission_gate_4/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X213 c1_n1700_3700# m3_n1800_3600# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X214 on p1 transmission_gate_3/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X215 transmission_gate_3/out p1 on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X216 on p1 transmission_gate_3/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X217 on cmc sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X218 transmission_gate_3/out p1 on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X219 on p1 transmission_gate_3/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X220 transmission_gate_3/out p1 on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X221 on p2 transmission_gate_7/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X222 transmission_gate_3/out p2 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X223 transmission_gate_3/out transmission_gate_5/out sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X224 transmission_gate_4/out p2 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X225 on cmc sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X226 on p1 transmission_gate_3/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X227 op p2_b transmission_gate_6/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X228 transmission_gate_6/in p2 op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X229 transmission_gate_8/in p2_b cmc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X230 bias_a p2 transmission_gate_5/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X231 cm p2_b transmission_gate_3/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X232 c1_100_n1700# m3_0_n1800# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X233 transmission_gate_8/in p1 bias_a VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X234 transmission_gate_8/in p1_b bias_a VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X235 transmission_gate_5/out p1_b cmc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X236 transmission_gate_5/out p1 cmc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X237 cm p1_b transmission_gate_6/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X238 on p2_b transmission_gate_7/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X239 transmission_gate_4/out p2_b cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X240 transmission_gate_6/in p1 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X241 bias_a p1 transmission_gate_8/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X242 bias_a p1_b transmission_gate_8/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X243 transmission_gate_6/in p2_b op VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X244 bias_a p2_b transmission_gate_5/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X245 cm p2 transmission_gate_3/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X246 op p1 transmission_gate_4/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X247 transmission_gate_5/out p2 bias_a VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X248 transmission_gate_7/in p2 on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X249 transmission_gate_8/in p2 cmc VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X250 op p1_b transmission_gate_4/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X251 transmission_gate_4/out p2 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X252 cmc p2_b transmission_gate_8/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X253 transmission_gate_6/in p1_b cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X254 c1_100_7300# m3_0_7200# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X255 transmission_gate_3/out p2_b cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X256 transmission_gate_7/in p2_b on VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X257 transmission_gate_6/in transmission_gate_8/in sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X258 transmission_gate_4/out transmission_gate_5/out sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X259 cm p2_b transmission_gate_4/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X260 op p2_b transmission_gate_6/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X261 transmission_gate_5/out p2_b bias_a VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X262 cmc p2 transmission_gate_8/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X263 op p1 transmission_gate_4/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X264 transmission_gate_3/out p2 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X265 op p1_b transmission_gate_4/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X266 bias_a p2 transmission_gate_5/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X267 transmission_gate_6/in p2 op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X268 c1_7300_n1700# m3_7200_n1800# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X269 transmission_gate_8/in p2_b cmc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X270 cm p1_b transmission_gate_6/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X271 transmission_gate_4/out p1 op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=530000u l=150000u
X272 transmission_gate_4/out p2_b cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X273 transmission_gate_5/out p1_b cmc VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X274 transmission_gate_4/out p1_b op VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
X275 transmission_gate_3/out p2_b cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.37e+06u l=150000u
.ends

