magic
tech sky130A
magscale 1 2
timestamp 1654720771
<< nwell >>
rect -2386 -1234 -1092 -1157
<< pwell >>
rect -528 -702 -409 -700
rect -548 -855 -231 -702
rect -548 -1692 -405 -1537
rect -548 -1693 -429 -1692
<< locali >>
rect -2626 115 3466 243
rect -2599 -493 -2335 -429
rect -2599 -2678 -2535 -493
rect -1186 -1162 -1122 -1123
rect -870 -1162 -806 115
rect -626 -684 -510 -620
rect -74 -1077 -10 115
rect 1637 -51 3236 13
rect 1637 -169 1701 -51
rect 3172 -102 3236 -51
rect 3038 -166 3236 -102
rect -74 -1141 348 -1077
rect -1186 -1226 -371 -1162
rect -74 -1195 -10 -1141
rect 1647 -1195 1711 -1074
rect -1186 -1269 -1122 -1226
rect -74 -1259 1711 -1195
rect -697 -1718 -501 -1710
rect -697 -1779 -690 -1718
rect -626 -1779 -501 -1718
rect -626 -1782 -625 -1779
rect -1204 -2678 -1140 -2268
rect -689 -2678 -625 -1782
rect -74 -2410 -10 -1259
rect 3172 -1336 3236 -166
rect 1645 -1400 3236 -1336
rect 1645 -1488 1709 -1400
rect 3172 -1442 3236 -1400
rect 3034 -1506 3236 -1442
rect -74 -2474 334 -2410
rect -74 -2529 -10 -2474
rect 1643 -2529 1707 -2423
rect -74 -2593 1707 -2529
rect 3172 -2678 3236 -1506
rect -2626 -2806 3466 -2678
<< viali >>
rect -1276 -231 -1242 -197
rect -1276 -1042 -1242 -1008
rect -690 -684 -626 -620
rect -298 -812 -264 -778
rect -381 -907 -347 -873
rect -1276 -1386 -1242 -1352
rect -299 -1382 -265 -1348
rect -382 -1520 -348 -1486
rect -690 -1782 -626 -1718
rect -1276 -2197 -1242 -2163
<< metal1 >>
rect -1297 -240 -1287 -188
rect -1235 -240 -1225 -188
rect -1046 -479 104 -445
rect -1046 -513 -1012 -479
rect -2638 -547 -2375 -513
rect -1271 -547 -1012 -513
rect 70 -503 104 -479
rect 70 -547 296 -503
rect 3055 -547 3258 -513
rect 71 -555 296 -547
rect -702 -620 -614 -614
rect -702 -684 -690 -620
rect -626 -684 -614 -620
rect -702 -690 -614 -684
rect -528 -700 -522 -604
rect -43 -772 -33 -769
rect -310 -778 -33 -772
rect -310 -812 -298 -778
rect -264 -812 -33 -778
rect -310 -818 -33 -812
rect -43 -821 -33 -818
rect 19 -821 29 -769
rect -401 -917 -391 -865
rect -339 -917 -329 -865
rect 139 -1000 149 -997
rect -1298 -1052 -1288 -1000
rect -1236 -1052 -1226 -1000
rect -176 -1052 -166 -1000
rect -114 -1049 149 -1000
rect 201 -1049 211 -997
rect -114 -1052 198 -1049
rect 3224 -1270 3258 -547
rect 3224 -1304 3429 -1270
rect -1295 -1395 -1285 -1343
rect -1233 -1395 -1223 -1343
rect -1025 -1394 -1015 -1342
rect -963 -1348 -253 -1342
rect -963 -1382 -299 -1348
rect -265 -1382 -253 -1348
rect -963 -1388 -253 -1382
rect -963 -1394 -953 -1388
rect -401 -1530 -391 -1478
rect -339 -1530 -329 -1478
rect -702 -1718 -614 -1712
rect -702 -1782 -690 -1718
rect -626 -1782 -614 -1718
rect -702 -1788 -614 -1782
rect -2638 -1881 -2375 -1847
rect -1272 -1881 -989 -1847
rect -1023 -2007 -989 -1881
rect -875 -1910 -865 -1858
rect -813 -1910 -390 -1858
rect -338 -1910 -328 -1858
rect 69 -1889 303 -1837
rect 3224 -1847 3258 -1304
rect 3052 -1881 3258 -1847
rect 69 -2007 103 -1889
rect -1023 -2041 103 -2007
rect -1296 -2206 -1286 -2154
rect -1234 -2206 -1224 -2154
<< via1 >>
rect -1287 -197 -1235 -188
rect -1287 -231 -1276 -197
rect -1276 -231 -1242 -197
rect -1242 -231 -1235 -197
rect -1287 -240 -1235 -231
rect -690 -684 -626 -620
rect -33 -821 19 -769
rect -391 -873 -339 -865
rect -391 -907 -381 -873
rect -381 -907 -347 -873
rect -347 -907 -339 -873
rect -391 -917 -339 -907
rect -1288 -1008 -1236 -1000
rect -1288 -1042 -1276 -1008
rect -1276 -1042 -1242 -1008
rect -1242 -1042 -1236 -1008
rect -1288 -1052 -1236 -1042
rect -166 -1052 -114 -1000
rect 149 -1049 201 -997
rect -1285 -1352 -1233 -1343
rect -1285 -1386 -1276 -1352
rect -1276 -1386 -1242 -1352
rect -1242 -1386 -1233 -1352
rect -1285 -1395 -1233 -1386
rect -1015 -1394 -963 -1342
rect -391 -1486 -339 -1478
rect -391 -1520 -382 -1486
rect -382 -1520 -348 -1486
rect -348 -1520 -339 -1486
rect -391 -1530 -339 -1520
rect -690 -1782 -626 -1718
rect -865 -1910 -813 -1858
rect -390 -1910 -338 -1858
rect -1286 -2163 -1234 -2154
rect -1286 -2197 -1276 -2163
rect -1276 -2197 -1242 -2163
rect -1242 -2197 -1234 -2163
rect -1286 -2206 -1234 -2197
<< metal2 >>
rect -1287 -188 -1235 -178
rect -1306 -240 -1287 -192
rect -1235 -240 -813 -192
rect -1306 -244 -813 -240
rect -1287 -250 -1235 -244
rect -1288 -1000 -1236 -990
rect -1312 -1052 -1288 -1000
rect -1236 -1052 -963 -1000
rect -1288 -1062 -1236 -1052
rect -1285 -1342 -1233 -1333
rect -1015 -1342 -963 -1052
rect -1285 -1343 -1015 -1342
rect -1233 -1394 -1015 -1343
rect -1285 -1405 -1233 -1395
rect -1015 -1404 -963 -1394
rect -865 -1858 -813 -244
rect -690 -620 -626 -610
rect -690 -1718 -626 -684
rect -391 -865 -339 115
rect -391 -1000 -339 -917
rect -33 -245 261 -193
rect -33 -769 19 -245
rect -166 -1000 -114 -990
rect -391 -1052 -166 -1000
rect -166 -1062 -114 -1052
rect -690 -1792 -626 -1782
rect -391 -1478 -339 -1468
rect -1286 -2149 -1234 -2144
rect -865 -2149 -813 -1910
rect -1297 -2154 -813 -2149
rect -1297 -2201 -1286 -2154
rect -1234 -2201 -813 -2154
rect -391 -1848 -339 -1530
rect -391 -1858 -338 -1848
rect -391 -1910 -390 -1858
rect -391 -1920 -338 -1910
rect -1286 -2216 -1234 -2206
rect -391 -2457 -339 -1920
rect -33 -2334 19 -821
rect 149 -997 201 -987
rect 201 -1049 259 -1000
rect 149 -1052 259 -1049
rect 149 -1527 201 -1052
rect 149 -1579 305 -1527
rect 149 -1589 201 -1579
rect -33 -2386 261 -2334
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1654309566
transform 1 0 -459 0 1 -1740
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1654309566
transform 1 0 -459 0 -1 -652
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1650294714
transform 1 0 -551 0 1 -1740
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1650294714
transform -1 0 -459 0 -1 -652
box -38 -48 130 592
use switch_5t_mux2  switch_5t_mux2_0
timestamp 1654720150
transform 1 0 123 0 -1 -1396
box 92 4 2977 1118
use switch_5t_mux2  switch_5t_mux2_1
timestamp 1654720150
transform 1 0 123 0 -1 -62
box 92 4 2977 1118
use transmission_gate  transmission_gate_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout_v2/transmission_gate
timestamp 1654720150
transform 1 0 -2333 0 -1 -117
box -53 -49 1241 1063
use transmission_gate  transmission_gate_1
timestamp 1654720150
transform 1 0 -2333 0 1 -2277
box -53 -49 1241 1063
<< labels >>
flabel metal1 -2635 -530 -2635 -530 3 FreeSans 400 0 0 0 in0
port 3 e
flabel metal1 -2634 -1864 -2634 -1864 3 FreeSans 400 0 0 0 in1
port 4 e
flabel metal2 -365 -2445 -365 -2445 1 FreeSans 400 0 0 0 en
port 1 n
flabel metal1 3423 -1288 3423 -1288 1 FreeSans 400 0 0 0 out
port 5 n
flabel metal2 -366 110 -366 110 5 FreeSans 400 0 0 0 s0
port 2 s
flabel locali -2575 182 -2575 182 1 FreeSans 400 0 0 0 VDD
port 6 n power bidirectional
flabel locali -2569 -2738 -2569 -2738 1 FreeSans 400 0 0 0 VSS
port 7 n power bidirectional
<< end >>
