magic
tech sky130A
magscale 1 2
timestamp 1654583406
<< nwell >>
rect -38 261 2246 582
<< pwell >>
rect 347 21 1863 157
rect 29 -17 63 17
<< scnmos >>
rect 426 47 456 131
rect 512 47 542 131
rect 598 47 628 131
rect 684 47 714 131
rect 770 47 800 131
rect 856 47 886 131
rect 949 47 979 131
rect 1066 47 1096 131
rect 1152 47 1182 131
rect 1238 47 1268 131
rect 1324 47 1354 131
rect 1410 47 1440 131
rect 1496 47 1526 131
rect 1582 47 1612 131
rect 1668 47 1698 131
rect 1754 47 1784 131
<< scpmoshvt >>
rect 82 297 112 497
rect 168 297 198 497
rect 254 297 284 497
rect 340 297 370 497
rect 426 297 456 497
rect 512 297 542 497
rect 598 297 628 497
rect 684 297 714 497
rect 770 297 800 497
rect 856 297 886 497
rect 949 297 979 497
rect 1066 297 1096 497
rect 1152 297 1182 497
rect 1238 297 1268 497
rect 1324 297 1354 497
rect 1410 297 1440 497
rect 1496 297 1526 497
rect 1582 297 1612 497
rect 1668 297 1698 497
rect 1754 297 1784 497
rect 1840 297 1870 497
rect 1926 297 1956 497
rect 2012 297 2042 497
rect 2098 297 2128 497
<< ndiff >>
rect 373 106 426 131
rect 373 72 381 106
rect 415 72 426 106
rect 373 47 426 72
rect 456 106 512 131
rect 456 72 467 106
rect 501 72 512 106
rect 456 47 512 72
rect 542 106 598 131
rect 542 72 553 106
rect 587 72 598 106
rect 542 47 598 72
rect 628 106 684 131
rect 628 72 639 106
rect 673 72 684 106
rect 628 47 684 72
rect 714 106 770 131
rect 714 72 725 106
rect 759 72 770 106
rect 714 47 770 72
rect 800 106 856 131
rect 800 72 811 106
rect 845 72 856 106
rect 800 47 856 72
rect 886 106 949 131
rect 886 72 902 106
rect 936 72 949 106
rect 886 47 949 72
rect 979 106 1066 131
rect 979 72 996 106
rect 1030 72 1066 106
rect 979 47 1066 72
rect 1096 106 1152 131
rect 1096 72 1107 106
rect 1141 72 1152 106
rect 1096 47 1152 72
rect 1182 106 1238 131
rect 1182 72 1193 106
rect 1227 72 1238 106
rect 1182 47 1238 72
rect 1268 106 1324 131
rect 1268 72 1279 106
rect 1313 72 1324 106
rect 1268 47 1324 72
rect 1354 106 1410 131
rect 1354 72 1365 106
rect 1399 72 1410 106
rect 1354 47 1410 72
rect 1440 106 1496 131
rect 1440 72 1451 106
rect 1485 72 1496 106
rect 1440 47 1496 72
rect 1526 106 1582 131
rect 1526 72 1537 106
rect 1571 72 1582 106
rect 1526 47 1582 72
rect 1612 106 1668 131
rect 1612 72 1623 106
rect 1657 72 1668 106
rect 1612 47 1668 72
rect 1698 106 1754 131
rect 1698 72 1709 106
rect 1743 72 1754 106
rect 1698 47 1754 72
rect 1784 106 1837 131
rect 1784 72 1795 106
rect 1829 72 1837 106
rect 1784 47 1837 72
<< pdiff >>
rect 27 485 82 497
rect 27 451 38 485
rect 72 451 82 485
rect 27 417 82 451
rect 27 383 38 417
rect 72 383 82 417
rect 27 349 82 383
rect 27 315 38 349
rect 72 315 82 349
rect 27 297 82 315
rect 112 477 168 497
rect 112 443 123 477
rect 157 443 168 477
rect 112 409 168 443
rect 112 375 123 409
rect 157 375 168 409
rect 112 341 168 375
rect 112 307 123 341
rect 157 307 168 341
rect 112 297 168 307
rect 198 485 254 497
rect 198 451 209 485
rect 243 451 254 485
rect 198 417 254 451
rect 198 383 209 417
rect 243 383 254 417
rect 198 297 254 383
rect 284 474 340 497
rect 284 440 295 474
rect 329 440 340 474
rect 284 341 340 440
rect 284 307 295 341
rect 329 307 340 341
rect 284 297 340 307
rect 370 485 426 497
rect 370 451 381 485
rect 415 451 426 485
rect 370 417 426 451
rect 370 383 381 417
rect 415 383 426 417
rect 370 297 426 383
rect 456 474 512 497
rect 456 440 467 474
rect 501 440 512 474
rect 456 341 512 440
rect 456 307 467 341
rect 501 307 512 341
rect 456 297 512 307
rect 542 485 598 497
rect 542 451 553 485
rect 587 451 598 485
rect 542 417 598 451
rect 542 383 553 417
rect 587 383 598 417
rect 542 297 598 383
rect 628 474 684 497
rect 628 440 639 474
rect 673 440 684 474
rect 628 341 684 440
rect 628 307 639 341
rect 673 307 684 341
rect 628 297 684 307
rect 714 485 770 497
rect 714 451 725 485
rect 759 451 770 485
rect 714 417 770 451
rect 714 383 725 417
rect 759 383 770 417
rect 714 297 770 383
rect 800 474 856 497
rect 800 440 811 474
rect 845 440 856 474
rect 800 341 856 440
rect 800 307 811 341
rect 845 307 856 341
rect 800 297 856 307
rect 886 485 949 497
rect 886 451 901 485
rect 935 451 949 485
rect 886 417 949 451
rect 886 383 901 417
rect 935 383 949 417
rect 886 297 949 383
rect 979 474 1066 497
rect 979 440 1016 474
rect 1050 440 1066 474
rect 979 341 1066 440
rect 979 307 1016 341
rect 1050 307 1066 341
rect 979 297 1066 307
rect 1096 485 1152 497
rect 1096 451 1106 485
rect 1140 451 1152 485
rect 1096 417 1152 451
rect 1096 383 1106 417
rect 1140 383 1152 417
rect 1096 297 1152 383
rect 1182 474 1238 497
rect 1182 440 1193 474
rect 1227 440 1238 474
rect 1182 341 1238 440
rect 1182 307 1193 341
rect 1227 307 1238 341
rect 1182 297 1238 307
rect 1268 485 1324 497
rect 1268 451 1279 485
rect 1313 451 1324 485
rect 1268 417 1324 451
rect 1268 383 1279 417
rect 1313 383 1324 417
rect 1268 297 1324 383
rect 1354 474 1410 497
rect 1354 440 1365 474
rect 1399 440 1410 474
rect 1354 341 1410 440
rect 1354 307 1365 341
rect 1399 307 1410 341
rect 1354 297 1410 307
rect 1440 485 1496 497
rect 1440 451 1451 485
rect 1485 451 1496 485
rect 1440 417 1496 451
rect 1440 383 1451 417
rect 1485 383 1496 417
rect 1440 297 1496 383
rect 1526 474 1582 497
rect 1526 440 1537 474
rect 1571 440 1582 474
rect 1526 341 1582 440
rect 1526 307 1537 341
rect 1571 307 1582 341
rect 1526 297 1582 307
rect 1612 485 1668 497
rect 1612 451 1623 485
rect 1657 451 1668 485
rect 1612 417 1668 451
rect 1612 383 1623 417
rect 1657 383 1668 417
rect 1612 297 1668 383
rect 1698 474 1754 497
rect 1698 440 1709 474
rect 1743 440 1754 474
rect 1698 341 1754 440
rect 1698 307 1709 341
rect 1743 307 1754 341
rect 1698 297 1754 307
rect 1784 485 1840 497
rect 1784 451 1795 485
rect 1829 451 1840 485
rect 1784 417 1840 451
rect 1784 383 1795 417
rect 1829 383 1840 417
rect 1784 297 1840 383
rect 1870 474 1926 497
rect 1870 440 1881 474
rect 1915 440 1926 474
rect 1870 341 1926 440
rect 1870 307 1881 341
rect 1915 307 1926 341
rect 1870 297 1926 307
rect 1956 485 2012 497
rect 1956 451 1967 485
rect 2001 451 2012 485
rect 1956 417 2012 451
rect 1956 383 1967 417
rect 2001 383 2012 417
rect 1956 297 2012 383
rect 2042 474 2098 497
rect 2042 440 2053 474
rect 2087 440 2098 474
rect 2042 341 2098 440
rect 2042 307 2053 341
rect 2087 307 2098 341
rect 2042 297 2098 307
rect 2128 485 2181 497
rect 2128 451 2138 485
rect 2172 451 2181 485
rect 2128 417 2181 451
rect 2128 383 2138 417
rect 2172 383 2181 417
rect 2128 297 2181 383
<< ndiffc >>
rect 381 72 415 106
rect 467 72 501 106
rect 553 72 587 106
rect 639 72 673 106
rect 725 72 759 106
rect 811 72 845 106
rect 902 72 936 106
rect 996 72 1030 106
rect 1107 72 1141 106
rect 1193 72 1227 106
rect 1279 72 1313 106
rect 1365 72 1399 106
rect 1451 72 1485 106
rect 1537 72 1571 106
rect 1623 72 1657 106
rect 1709 72 1743 106
rect 1795 72 1829 106
<< pdiffc >>
rect 38 451 72 485
rect 38 383 72 417
rect 38 315 72 349
rect 123 443 157 477
rect 123 375 157 409
rect 123 307 157 341
rect 209 451 243 485
rect 209 383 243 417
rect 295 440 329 474
rect 295 307 329 341
rect 381 451 415 485
rect 381 383 415 417
rect 467 440 501 474
rect 467 307 501 341
rect 553 451 587 485
rect 553 383 587 417
rect 639 440 673 474
rect 639 307 673 341
rect 725 451 759 485
rect 725 383 759 417
rect 811 440 845 474
rect 811 307 845 341
rect 901 451 935 485
rect 901 383 935 417
rect 1016 440 1050 474
rect 1016 307 1050 341
rect 1106 451 1140 485
rect 1106 383 1140 417
rect 1193 440 1227 474
rect 1193 307 1227 341
rect 1279 451 1313 485
rect 1279 383 1313 417
rect 1365 440 1399 474
rect 1365 307 1399 341
rect 1451 451 1485 485
rect 1451 383 1485 417
rect 1537 440 1571 474
rect 1537 307 1571 341
rect 1623 451 1657 485
rect 1623 383 1657 417
rect 1709 440 1743 474
rect 1709 307 1743 341
rect 1795 451 1829 485
rect 1795 383 1829 417
rect 1881 440 1915 474
rect 1881 307 1915 341
rect 1967 451 2001 485
rect 1967 383 2001 417
rect 2053 440 2087 474
rect 2053 307 2087 341
rect 2138 451 2172 485
rect 2138 383 2172 417
<< poly >>
rect 82 497 112 523
rect 168 497 198 523
rect 254 497 284 523
rect 340 497 370 523
rect 426 497 456 523
rect 512 497 542 523
rect 598 497 628 523
rect 684 497 714 523
rect 770 497 800 523
rect 856 497 886 523
rect 949 497 979 523
rect 1066 497 1096 523
rect 1152 497 1182 523
rect 1238 497 1268 523
rect 1324 497 1354 523
rect 1410 497 1440 523
rect 1496 497 1526 523
rect 1582 497 1612 523
rect 1668 497 1698 523
rect 1754 497 1784 523
rect 1840 497 1870 523
rect 1926 497 1956 523
rect 2012 497 2042 523
rect 2098 497 2128 523
rect 82 270 112 297
rect 168 270 198 297
rect 254 270 284 297
rect 340 270 370 297
rect 426 270 456 297
rect 512 270 542 297
rect 598 270 628 297
rect 684 270 714 297
rect 770 270 800 297
rect 856 270 886 297
rect 949 270 979 297
rect 1066 270 1096 297
rect 1152 270 1182 297
rect 1238 270 1268 297
rect 1324 270 1354 297
rect 1410 270 1440 297
rect 1496 270 1526 297
rect 1582 270 1612 297
rect 1668 270 1698 297
rect 1754 270 1784 297
rect 1840 270 1870 297
rect 1926 270 1956 297
rect 2012 270 2042 297
rect 2098 270 2128 297
rect 82 249 2128 270
rect 82 215 101 249
rect 135 215 169 249
rect 203 215 237 249
rect 271 215 305 249
rect 339 215 373 249
rect 407 215 1803 249
rect 1837 215 1871 249
rect 1905 215 1939 249
rect 1973 215 2007 249
rect 2041 215 2075 249
rect 2109 215 2128 249
rect 82 198 2128 215
rect 426 131 456 198
rect 512 131 542 198
rect 598 131 628 198
rect 684 131 714 198
rect 770 131 800 198
rect 856 131 886 198
rect 949 131 979 198
rect 1066 131 1096 198
rect 1152 131 1182 198
rect 1238 131 1268 198
rect 1324 131 1354 198
rect 1410 131 1440 198
rect 1496 131 1526 198
rect 1582 131 1612 198
rect 1668 131 1698 198
rect 1754 131 1784 198
rect 426 21 456 47
rect 512 21 542 47
rect 598 21 628 47
rect 684 21 714 47
rect 770 21 800 47
rect 856 21 886 47
rect 949 21 979 47
rect 1066 21 1096 47
rect 1152 21 1182 47
rect 1238 21 1268 47
rect 1324 21 1354 47
rect 1410 21 1440 47
rect 1496 21 1526 47
rect 1582 21 1612 47
rect 1668 21 1698 47
rect 1754 21 1784 47
<< polycont >>
rect 101 215 135 249
rect 169 215 203 249
rect 237 215 271 249
rect 305 215 339 249
rect 373 215 407 249
rect 1803 215 1837 249
rect 1871 215 1905 249
rect 1939 215 1973 249
rect 2007 215 2041 249
rect 2075 215 2109 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 28 485 81 527
rect 28 451 38 485
rect 72 451 81 485
rect 28 417 81 451
rect 28 383 38 417
rect 72 383 81 417
rect 28 349 81 383
rect 28 315 38 349
rect 72 315 81 349
rect 28 299 81 315
rect 115 477 166 493
rect 115 443 123 477
rect 157 443 166 477
rect 115 409 166 443
rect 115 375 123 409
rect 157 375 166 409
rect 115 341 166 375
rect 200 485 252 527
rect 200 451 209 485
rect 243 451 252 485
rect 200 417 252 451
rect 200 383 209 417
rect 243 383 252 417
rect 200 367 252 383
rect 287 474 338 490
rect 287 440 295 474
rect 329 440 338 474
rect 115 307 123 341
rect 157 333 166 341
rect 287 341 338 440
rect 373 485 424 527
rect 373 451 381 485
rect 415 451 424 485
rect 373 417 424 451
rect 373 383 381 417
rect 415 383 424 417
rect 373 367 424 383
rect 465 474 510 493
rect 465 440 467 474
rect 501 440 510 474
rect 287 333 295 341
rect 157 307 295 333
rect 329 333 338 341
rect 465 341 510 440
rect 544 485 596 527
rect 544 451 553 485
rect 587 451 596 485
rect 544 417 596 451
rect 544 383 553 417
rect 587 383 596 417
rect 544 367 596 383
rect 631 474 682 490
rect 631 440 639 474
rect 673 440 682 474
rect 465 333 467 341
rect 329 307 467 333
rect 501 333 510 341
rect 631 341 682 440
rect 717 485 768 527
rect 717 451 725 485
rect 759 451 768 485
rect 717 417 768 451
rect 717 383 725 417
rect 759 383 768 417
rect 717 367 768 383
rect 803 474 851 490
rect 803 440 811 474
rect 845 440 851 474
rect 631 333 639 341
rect 501 307 639 333
rect 673 333 682 341
rect 803 341 851 440
rect 893 485 944 527
rect 893 451 901 485
rect 935 451 944 485
rect 893 417 944 451
rect 893 383 901 417
rect 935 383 944 417
rect 893 367 944 383
rect 981 474 1056 490
rect 981 440 1016 474
rect 1050 440 1056 474
rect 803 333 811 341
rect 673 307 811 333
rect 845 333 851 341
rect 981 341 1056 440
rect 1098 485 1150 527
rect 1098 451 1106 485
rect 1140 451 1150 485
rect 1098 424 1150 451
rect 1185 474 1235 490
rect 1185 440 1193 474
rect 1227 440 1235 474
rect 1098 417 1149 424
rect 1098 383 1106 417
rect 1140 383 1149 417
rect 1098 367 1149 383
rect 981 333 1016 341
rect 845 307 1016 333
rect 1050 333 1056 341
rect 1185 341 1235 440
rect 1271 485 1322 527
rect 1271 451 1279 485
rect 1313 451 1322 485
rect 1271 417 1322 451
rect 1271 383 1279 417
rect 1313 383 1322 417
rect 1271 367 1322 383
rect 1357 474 1407 490
rect 1357 440 1365 474
rect 1399 440 1407 474
rect 1185 333 1193 341
rect 1050 307 1193 333
rect 1227 333 1235 341
rect 1357 341 1407 440
rect 1443 485 1494 527
rect 1443 451 1451 485
rect 1485 451 1494 485
rect 1443 417 1494 451
rect 1443 383 1451 417
rect 1485 383 1494 417
rect 1443 367 1494 383
rect 1529 474 1579 490
rect 1529 440 1537 474
rect 1571 440 1579 474
rect 1357 333 1365 341
rect 1227 307 1365 333
rect 1399 333 1407 341
rect 1529 341 1579 440
rect 1615 485 1666 527
rect 1615 451 1623 485
rect 1657 451 1666 485
rect 1615 417 1666 451
rect 1615 383 1623 417
rect 1657 383 1666 417
rect 1615 367 1666 383
rect 1701 474 1751 490
rect 1701 440 1709 474
rect 1743 440 1751 474
rect 1529 333 1537 341
rect 1399 307 1537 333
rect 1571 333 1579 341
rect 1701 341 1751 440
rect 1787 485 1838 527
rect 1787 451 1795 485
rect 1829 451 1838 485
rect 1787 417 1838 451
rect 1787 383 1795 417
rect 1829 383 1838 417
rect 1787 367 1838 383
rect 1873 474 1921 490
rect 1873 440 1881 474
rect 1915 440 1921 474
rect 1701 333 1709 341
rect 1571 307 1709 333
rect 1743 333 1751 341
rect 1873 341 1921 440
rect 1959 485 2010 527
rect 1959 451 1967 485
rect 2001 451 2010 485
rect 1959 417 2010 451
rect 1959 383 1967 417
rect 2001 383 2010 417
rect 1959 367 2010 383
rect 2045 474 2096 490
rect 2045 440 2053 474
rect 2087 440 2096 474
rect 1873 333 1881 341
rect 1743 307 1881 333
rect 1915 333 1921 341
rect 2045 341 2096 440
rect 2130 485 2182 527
rect 2130 451 2138 485
rect 2172 451 2182 485
rect 2130 417 2182 451
rect 2130 383 2138 417
rect 2172 383 2182 417
rect 2130 367 2182 383
rect 2045 333 2053 341
rect 1915 307 2053 333
rect 2087 307 2096 341
rect 115 291 2096 307
rect 465 283 1751 291
rect 69 249 305 255
rect 339 249 397 255
rect 69 215 101 249
rect 135 215 169 249
rect 203 215 237 249
rect 271 215 305 249
rect 339 215 373 249
rect 407 215 431 221
rect 69 179 431 215
rect 371 106 425 122
rect 371 72 381 106
rect 415 72 425 106
rect 371 17 425 72
rect 465 106 510 283
rect 465 72 467 106
rect 501 72 510 106
rect 465 56 510 72
rect 544 106 597 122
rect 544 72 553 106
rect 587 72 597 106
rect 544 17 597 72
rect 631 106 682 283
rect 631 72 639 106
rect 673 72 682 106
rect 631 56 682 72
rect 716 106 769 122
rect 716 72 725 106
rect 759 72 769 106
rect 716 17 769 72
rect 803 106 851 283
rect 803 72 811 106
rect 845 72 851 106
rect 803 56 851 72
rect 893 106 946 122
rect 893 72 902 106
rect 936 72 946 106
rect 893 17 946 72
rect 981 106 1051 283
rect 981 72 996 106
rect 1030 72 1051 106
rect 981 56 1051 72
rect 1098 106 1151 122
rect 1098 72 1107 106
rect 1141 72 1151 106
rect 1098 17 1151 72
rect 1185 106 1235 283
rect 1185 72 1193 106
rect 1227 72 1235 106
rect 1185 56 1235 72
rect 1270 106 1315 122
rect 1270 72 1279 106
rect 1313 72 1315 106
rect 1270 17 1315 72
rect 1357 106 1407 283
rect 1357 72 1365 106
rect 1399 72 1407 106
rect 1357 56 1407 72
rect 1442 106 1495 122
rect 1442 72 1451 106
rect 1485 72 1495 106
rect 1442 17 1495 72
rect 1529 106 1579 283
rect 1529 72 1537 106
rect 1571 72 1579 106
rect 1529 56 1579 72
rect 1614 106 1667 122
rect 1614 72 1623 106
rect 1657 72 1667 106
rect 1614 17 1667 72
rect 1701 106 1751 283
rect 1786 249 1869 255
rect 1903 249 1961 255
rect 1995 249 2142 255
rect 1786 215 1803 249
rect 1837 221 1869 249
rect 1837 215 1871 221
rect 1905 215 1939 249
rect 1995 221 2007 249
rect 1973 215 2007 221
rect 2041 215 2075 249
rect 2109 215 2142 249
rect 1786 179 2142 215
rect 1701 72 1709 106
rect 1743 72 1751 106
rect 1701 56 1751 72
rect 1786 106 1839 122
rect 1786 72 1795 106
rect 1829 72 1839 106
rect 1786 17 1839 72
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 305 249 339 255
rect 397 249 431 255
rect 305 221 339 249
rect 397 221 407 249
rect 407 221 431 249
rect 1869 249 1903 255
rect 1961 249 1995 255
rect 1869 221 1871 249
rect 1871 221 1903 249
rect 1961 221 1973 249
rect 1973 221 1995 249
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
<< metal1 >>
rect 0 561 2208 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 0 496 2208 527
rect 293 255 443 261
rect 293 221 305 255
rect 339 221 397 255
rect 431 252 443 255
rect 1857 255 2007 261
rect 1857 252 1869 255
rect 431 224 1869 252
rect 431 221 443 224
rect 293 215 443 221
rect 1857 221 1869 224
rect 1903 221 1961 255
rect 1995 221 2007 255
rect 1857 215 2007 221
rect 0 17 2208 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
rect 0 -48 2208 -17
<< labels >>
flabel locali s 1041 289 1075 323 0 FreeSans 400 0 0 0 Y
port 1 nsew
flabel locali s 397 221 431 255 0 FreeSans 400 0 0 0 A
port 2 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 4 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew
rlabel comment s 0 0 0 0 4 clkinv_16
<< properties >>
string FIXED_BBOX 0 0 2208 544
string path 0.000 0.000 11.040 0.000 
<< end >>
