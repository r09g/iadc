magic
tech sky130A
timestamp 1654711401
<< metal3 >>
rect -515 -490 464 490
<< mimcap >>
rect -465 420 414 440
rect -465 -420 -445 420
rect 394 -420 414 420
rect -465 -440 414 -420
<< mimcapcontact >>
rect -445 -420 394 420
<< metal4 >>
rect -446 -420 -445 420
rect 394 -420 395 420
<< properties >>
string FIXED_BBOX -515 -490 465 490
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 8.8 l 8.8 val 161.568 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 1 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
