magic
tech sky130A
timestamp 1654517900
<< nwell >>
rect -744 -120 744 120
<< pmoslvt >>
rect -697 -70 -637 70
rect -608 -70 -548 70
rect -519 -70 -459 70
rect -430 -70 -370 70
rect -341 -70 -281 70
rect -252 -70 -192 70
rect -163 -70 -103 70
rect -74 -70 -14 70
rect 14 -70 74 70
rect 103 -70 163 70
rect 192 -70 252 70
rect 281 -70 341 70
rect 370 -70 430 70
rect 459 -70 519 70
rect 548 -70 608 70
rect 637 -70 697 70
<< pdiff >>
rect -726 64 -697 70
rect -726 -64 -720 64
rect -703 -64 -697 64
rect -726 -70 -697 -64
rect -637 64 -608 70
rect -637 -64 -631 64
rect -614 -64 -608 64
rect -637 -70 -608 -64
rect -548 64 -519 70
rect -548 -64 -542 64
rect -525 -64 -519 64
rect -548 -70 -519 -64
rect -459 64 -430 70
rect -459 -64 -453 64
rect -436 -64 -430 64
rect -459 -70 -430 -64
rect -370 64 -341 70
rect -370 -64 -364 64
rect -347 -64 -341 64
rect -370 -70 -341 -64
rect -281 64 -252 70
rect -281 -64 -275 64
rect -258 -64 -252 64
rect -281 -70 -252 -64
rect -192 64 -163 70
rect -192 -64 -186 64
rect -169 -64 -163 64
rect -192 -70 -163 -64
rect -103 64 -74 70
rect -103 -64 -97 64
rect -80 -64 -74 64
rect -103 -70 -74 -64
rect -14 64 14 70
rect -14 -64 -8 64
rect 8 -64 14 64
rect -14 -70 14 -64
rect 74 64 103 70
rect 74 -64 80 64
rect 97 -64 103 64
rect 74 -70 103 -64
rect 163 64 192 70
rect 163 -64 169 64
rect 186 -64 192 64
rect 163 -70 192 -64
rect 252 64 281 70
rect 252 -64 258 64
rect 275 -64 281 64
rect 252 -70 281 -64
rect 341 64 370 70
rect 341 -64 347 64
rect 364 -64 370 64
rect 341 -70 370 -64
rect 430 64 459 70
rect 430 -64 436 64
rect 453 -64 459 64
rect 430 -70 459 -64
rect 519 64 548 70
rect 519 -64 525 64
rect 542 -64 548 64
rect 519 -70 548 -64
rect 608 64 637 70
rect 608 -64 614 64
rect 631 -64 637 64
rect 608 -70 637 -64
rect 697 64 726 70
rect 697 -64 703 64
rect 720 -64 726 64
rect 697 -70 726 -64
<< pdiffc >>
rect -720 -64 -703 64
rect -631 -64 -614 64
rect -542 -64 -525 64
rect -453 -64 -436 64
rect -364 -64 -347 64
rect -275 -64 -258 64
rect -186 -64 -169 64
rect -97 -64 -80 64
rect -8 -64 8 64
rect 80 -64 97 64
rect 169 -64 186 64
rect 258 -64 275 64
rect 347 -64 364 64
rect 436 -64 453 64
rect 525 -64 542 64
rect 614 -64 631 64
rect 703 -64 720 64
<< poly >>
rect -686 110 -648 118
rect -686 102 -678 110
rect -697 93 -678 102
rect -656 102 -648 110
rect -597 110 -559 118
rect -597 102 -589 110
rect -656 93 -637 102
rect -697 70 -637 93
rect -608 93 -589 102
rect -567 102 -559 110
rect -508 110 -470 118
rect -508 102 -500 110
rect -567 93 -548 102
rect -608 70 -548 93
rect -519 93 -500 102
rect -478 102 -470 110
rect -419 110 -381 118
rect -419 102 -411 110
rect -478 93 -459 102
rect -519 70 -459 93
rect -430 93 -411 102
rect -389 102 -381 110
rect -330 110 -292 118
rect -330 102 -322 110
rect -389 93 -370 102
rect -430 70 -370 93
rect -341 93 -322 102
rect -300 102 -292 110
rect -241 110 -203 118
rect -241 102 -233 110
rect -300 93 -281 102
rect -341 70 -281 93
rect -252 93 -233 102
rect -211 102 -203 110
rect -152 110 -114 118
rect -152 102 -144 110
rect -211 93 -192 102
rect -252 70 -192 93
rect -163 93 -144 102
rect -122 102 -114 110
rect -63 110 -25 118
rect -63 102 -55 110
rect -122 93 -103 102
rect -163 70 -103 93
rect -74 93 -55 102
rect -33 102 -25 110
rect 25 110 63 118
rect 25 102 33 110
rect -33 93 -14 102
rect -74 70 -14 93
rect 14 93 33 102
rect 55 102 63 110
rect 114 110 152 118
rect 114 102 122 110
rect 55 93 74 102
rect 14 70 74 93
rect 103 93 122 102
rect 144 102 152 110
rect 203 110 241 118
rect 203 102 211 110
rect 144 93 163 102
rect 103 70 163 93
rect 192 93 211 102
rect 233 102 241 110
rect 292 110 330 118
rect 292 102 300 110
rect 233 93 252 102
rect 192 70 252 93
rect 281 93 300 102
rect 322 102 330 110
rect 381 110 419 118
rect 381 102 389 110
rect 322 93 341 102
rect 281 70 341 93
rect 370 93 389 102
rect 411 102 419 110
rect 470 110 508 118
rect 470 102 478 110
rect 411 93 430 102
rect 370 70 430 93
rect 459 93 478 102
rect 500 102 508 110
rect 559 110 597 118
rect 559 102 567 110
rect 500 93 519 102
rect 459 70 519 93
rect 548 93 567 102
rect 589 102 597 110
rect 648 110 686 118
rect 648 102 656 110
rect 589 93 608 102
rect 548 70 608 93
rect 637 93 656 102
rect 678 102 686 110
rect 678 93 697 102
rect 637 70 697 93
rect -697 -93 -637 -70
rect -697 -102 -678 -93
rect -686 -110 -678 -102
rect -656 -102 -637 -93
rect -608 -93 -548 -70
rect -608 -102 -589 -93
rect -656 -110 -648 -102
rect -686 -118 -648 -110
rect -597 -110 -589 -102
rect -567 -102 -548 -93
rect -519 -93 -459 -70
rect -519 -102 -500 -93
rect -567 -110 -559 -102
rect -597 -118 -559 -110
rect -508 -110 -500 -102
rect -478 -102 -459 -93
rect -430 -93 -370 -70
rect -430 -102 -411 -93
rect -478 -110 -470 -102
rect -508 -118 -470 -110
rect -419 -110 -411 -102
rect -389 -102 -370 -93
rect -341 -93 -281 -70
rect -341 -102 -322 -93
rect -389 -110 -381 -102
rect -419 -118 -381 -110
rect -330 -110 -322 -102
rect -300 -102 -281 -93
rect -252 -93 -192 -70
rect -252 -102 -233 -93
rect -300 -110 -292 -102
rect -330 -118 -292 -110
rect -241 -110 -233 -102
rect -211 -102 -192 -93
rect -163 -93 -103 -70
rect -163 -102 -144 -93
rect -211 -110 -203 -102
rect -241 -118 -203 -110
rect -152 -110 -144 -102
rect -122 -102 -103 -93
rect -74 -93 -14 -70
rect -74 -102 -55 -93
rect -122 -110 -114 -102
rect -152 -118 -114 -110
rect -63 -110 -55 -102
rect -33 -102 -14 -93
rect 14 -93 74 -70
rect 14 -102 33 -93
rect -33 -110 -25 -102
rect -63 -118 -25 -110
rect 25 -110 33 -102
rect 55 -102 74 -93
rect 103 -93 163 -70
rect 103 -102 122 -93
rect 55 -110 63 -102
rect 25 -118 63 -110
rect 114 -110 122 -102
rect 144 -102 163 -93
rect 192 -93 252 -70
rect 192 -102 211 -93
rect 144 -110 152 -102
rect 114 -118 152 -110
rect 203 -110 211 -102
rect 233 -102 252 -93
rect 281 -93 341 -70
rect 281 -102 300 -93
rect 233 -110 241 -102
rect 203 -118 241 -110
rect 292 -110 300 -102
rect 322 -102 341 -93
rect 370 -93 430 -70
rect 370 -102 389 -93
rect 322 -110 330 -102
rect 292 -118 330 -110
rect 381 -110 389 -102
rect 411 -102 430 -93
rect 459 -93 519 -70
rect 459 -102 478 -93
rect 411 -110 419 -102
rect 381 -118 419 -110
rect 470 -110 478 -102
rect 500 -102 519 -93
rect 548 -93 608 -70
rect 548 -102 567 -93
rect 500 -110 508 -102
rect 470 -118 508 -110
rect 559 -110 567 -102
rect 589 -102 608 -93
rect 637 -93 697 -70
rect 637 -102 656 -93
rect 589 -110 597 -102
rect 559 -118 597 -110
rect 648 -110 656 -102
rect 678 -102 697 -93
rect 678 -110 686 -102
rect 648 -118 686 -110
<< polycont >>
rect -678 93 -656 110
rect -589 93 -567 110
rect -500 93 -478 110
rect -411 93 -389 110
rect -322 93 -300 110
rect -233 93 -211 110
rect -144 93 -122 110
rect -55 93 -33 110
rect 33 93 55 110
rect 122 93 144 110
rect 211 93 233 110
rect 300 93 322 110
rect 389 93 411 110
rect 478 93 500 110
rect 567 93 589 110
rect 656 93 678 110
rect -678 -110 -656 -93
rect -589 -110 -567 -93
rect -500 -110 -478 -93
rect -411 -110 -389 -93
rect -322 -110 -300 -93
rect -233 -110 -211 -93
rect -144 -110 -122 -93
rect -55 -110 -33 -93
rect 33 -110 55 -93
rect 122 -110 144 -93
rect 211 -110 233 -93
rect 300 -110 322 -93
rect 389 -110 411 -93
rect 478 -110 500 -93
rect 567 -110 589 -93
rect 656 -110 678 -93
<< locali >>
rect -686 93 -678 110
rect -656 93 -648 110
rect -597 93 -589 110
rect -567 93 -559 110
rect -508 93 -500 110
rect -478 93 -470 110
rect -419 93 -411 110
rect -389 93 -381 110
rect -330 93 -322 110
rect -300 93 -292 110
rect -241 93 -233 110
rect -211 93 -203 110
rect -152 93 -144 110
rect -122 93 -114 110
rect -63 93 -55 110
rect -33 93 -25 110
rect 25 93 33 110
rect 55 93 63 110
rect 114 93 122 110
rect 144 93 152 110
rect 203 93 211 110
rect 233 93 241 110
rect 292 93 300 110
rect 322 93 330 110
rect 381 93 389 110
rect 411 93 419 110
rect 470 93 478 110
rect 500 93 508 110
rect 559 93 567 110
rect 589 93 597 110
rect 648 93 656 110
rect 678 93 686 110
rect -720 64 -703 72
rect -720 -72 -703 -64
rect -631 64 -614 72
rect -631 -72 -614 -64
rect -542 64 -525 72
rect -542 -72 -525 -64
rect -453 64 -436 72
rect -453 -72 -436 -64
rect -364 64 -347 72
rect -364 -72 -347 -64
rect -275 64 -258 72
rect -275 -72 -258 -64
rect -186 64 -169 72
rect -186 -72 -169 -64
rect -97 64 -80 72
rect -97 -72 -80 -64
rect -8 64 8 72
rect -8 -72 8 -64
rect 80 64 97 72
rect 80 -72 97 -64
rect 169 64 186 72
rect 169 -72 186 -64
rect 258 64 275 72
rect 258 -72 275 -64
rect 347 64 364 72
rect 347 -72 364 -64
rect 436 64 453 72
rect 436 -72 453 -64
rect 525 64 542 72
rect 525 -72 542 -64
rect 614 64 631 72
rect 614 -72 631 -64
rect 703 64 720 72
rect 703 -72 720 -64
rect -686 -110 -678 -93
rect -656 -110 -648 -93
rect -597 -110 -589 -93
rect -567 -110 -559 -93
rect -508 -110 -500 -93
rect -478 -110 -470 -93
rect -419 -110 -411 -93
rect -389 -110 -381 -93
rect -330 -110 -322 -93
rect -300 -110 -292 -93
rect -241 -110 -233 -93
rect -211 -110 -203 -93
rect -152 -110 -144 -93
rect -122 -110 -114 -93
rect -63 -110 -55 -93
rect -33 -110 -25 -93
rect 25 -110 33 -93
rect 55 -110 63 -93
rect 114 -110 122 -93
rect 144 -110 152 -93
rect 203 -110 211 -93
rect 233 -110 241 -93
rect 292 -110 300 -93
rect 322 -110 330 -93
rect 381 -110 389 -93
rect 411 -110 419 -93
rect 470 -110 478 -93
rect 500 -110 508 -93
rect 559 -110 567 -93
rect 589 -110 597 -93
rect 648 -110 656 -93
rect 678 -110 686 -93
<< viali >>
rect -678 93 -656 110
rect -589 93 -567 110
rect -500 93 -478 110
rect -411 93 -389 110
rect -322 93 -300 110
rect -233 93 -211 110
rect -144 93 -122 110
rect -55 93 -33 110
rect 33 93 55 110
rect 122 93 144 110
rect 211 93 233 110
rect 300 93 322 110
rect 389 93 411 110
rect 478 93 500 110
rect 567 93 589 110
rect 656 93 678 110
rect -720 -64 -703 64
rect -631 -64 -614 64
rect -542 -64 -525 64
rect -453 -64 -436 64
rect -364 -64 -347 64
rect -275 -64 -258 64
rect -186 -64 -169 64
rect -97 -64 -80 64
rect -8 -64 8 64
rect 80 -64 97 64
rect 169 -64 186 64
rect 258 -64 275 64
rect 347 -64 364 64
rect 436 -64 453 64
rect 525 -64 542 64
rect 614 -64 631 64
rect 703 -64 720 64
rect -678 -110 -656 -93
rect -589 -110 -567 -93
rect -500 -110 -478 -93
rect -411 -110 -389 -93
rect -322 -110 -300 -93
rect -233 -110 -211 -93
rect -144 -110 -122 -93
rect -55 -110 -33 -93
rect 33 -110 55 -93
rect 122 -110 144 -93
rect 211 -110 233 -93
rect 300 -110 322 -93
rect 389 -110 411 -93
rect 478 -110 500 -93
rect 567 -110 589 -93
rect 656 -110 678 -93
<< metal1 >>
rect -686 110 -648 118
rect -686 93 -678 110
rect -656 93 -648 110
rect -686 90 -648 93
rect -597 110 -559 118
rect -597 93 -589 110
rect -567 93 -559 110
rect -597 90 -559 93
rect -508 110 -470 118
rect -508 93 -500 110
rect -478 93 -470 110
rect -508 90 -470 93
rect -419 110 -381 118
rect -419 93 -411 110
rect -389 93 -381 110
rect -419 90 -381 93
rect -330 110 -292 118
rect -330 93 -322 110
rect -300 93 -292 110
rect -330 90 -292 93
rect -241 110 -203 118
rect -241 93 -233 110
rect -211 93 -203 110
rect -241 90 -203 93
rect -152 110 -114 118
rect -152 93 -144 110
rect -122 93 -114 110
rect -152 90 -114 93
rect -63 110 -25 118
rect -63 93 -55 110
rect -33 93 -25 110
rect -63 90 -25 93
rect 25 110 63 118
rect 25 93 33 110
rect 55 93 63 110
rect 25 90 63 93
rect 114 110 152 118
rect 114 93 122 110
rect 144 93 152 110
rect 114 90 152 93
rect 203 110 241 118
rect 203 93 211 110
rect 233 93 241 110
rect 203 90 241 93
rect 292 110 330 118
rect 292 93 300 110
rect 322 93 330 110
rect 292 90 330 93
rect 381 110 419 118
rect 381 93 389 110
rect 411 93 419 110
rect 381 90 419 93
rect 470 110 508 118
rect 470 93 478 110
rect 500 93 508 110
rect 470 90 508 93
rect 559 110 597 118
rect 559 93 567 110
rect 589 93 597 110
rect 559 90 597 93
rect 648 110 686 118
rect 648 93 656 110
rect 678 93 686 110
rect 648 90 686 93
rect -723 64 -700 70
rect -723 -64 -720 64
rect -703 -64 -700 64
rect -723 -70 -700 -64
rect -634 64 -611 70
rect -634 -64 -631 64
rect -614 -64 -611 64
rect -634 -70 -611 -64
rect -545 64 -522 70
rect -545 -64 -542 64
rect -525 -64 -522 64
rect -545 -70 -522 -64
rect -456 64 -433 70
rect -456 -64 -453 64
rect -436 -64 -433 64
rect -456 -70 -433 -64
rect -367 64 -344 70
rect -367 -64 -364 64
rect -347 -64 -344 64
rect -367 -70 -344 -64
rect -278 64 -255 70
rect -278 -64 -275 64
rect -258 -64 -255 64
rect -278 -70 -255 -64
rect -189 64 -166 70
rect -189 -64 -186 64
rect -169 -64 -166 64
rect -189 -70 -166 -64
rect -100 64 -77 70
rect -100 -64 -97 64
rect -80 -64 -77 64
rect -100 -70 -77 -64
rect -11 64 11 70
rect -11 -64 -8 64
rect 8 -64 11 64
rect -11 -70 11 -64
rect 77 64 100 70
rect 77 -64 80 64
rect 97 -64 100 64
rect 77 -70 100 -64
rect 166 64 189 70
rect 166 -64 169 64
rect 186 -64 189 64
rect 166 -70 189 -64
rect 255 64 278 70
rect 255 -64 258 64
rect 275 -64 278 64
rect 255 -70 278 -64
rect 344 64 367 70
rect 344 -64 347 64
rect 364 -64 367 64
rect 344 -70 367 -64
rect 433 64 456 70
rect 433 -64 436 64
rect 453 -64 456 64
rect 433 -70 456 -64
rect 522 64 545 70
rect 522 -64 525 64
rect 542 -64 545 64
rect 522 -70 545 -64
rect 611 64 634 70
rect 611 -64 614 64
rect 631 -64 634 64
rect 611 -70 634 -64
rect 700 64 723 70
rect 700 -64 703 64
rect 720 -64 723 64
rect 700 -70 723 -64
rect -686 -93 -648 -90
rect -686 -110 -678 -93
rect -656 -110 -648 -93
rect -686 -118 -648 -110
rect -597 -93 -559 -90
rect -597 -110 -589 -93
rect -567 -110 -559 -93
rect -597 -118 -559 -110
rect -508 -93 -470 -90
rect -508 -110 -500 -93
rect -478 -110 -470 -93
rect -508 -118 -470 -110
rect -419 -93 -381 -90
rect -419 -110 -411 -93
rect -389 -110 -381 -93
rect -419 -118 -381 -110
rect -330 -93 -292 -90
rect -330 -110 -322 -93
rect -300 -110 -292 -93
rect -330 -118 -292 -110
rect -241 -93 -203 -90
rect -241 -110 -233 -93
rect -211 -110 -203 -93
rect -241 -118 -203 -110
rect -152 -93 -114 -90
rect -152 -110 -144 -93
rect -122 -110 -114 -93
rect -152 -118 -114 -110
rect -63 -93 -25 -90
rect -63 -110 -55 -93
rect -33 -110 -25 -93
rect -63 -118 -25 -110
rect 25 -93 63 -90
rect 25 -110 33 -93
rect 55 -110 63 -93
rect 25 -118 63 -110
rect 114 -93 152 -90
rect 114 -110 122 -93
rect 144 -110 152 -93
rect 114 -118 152 -110
rect 203 -93 241 -90
rect 203 -110 211 -93
rect 233 -110 241 -93
rect 203 -118 241 -110
rect 292 -93 330 -90
rect 292 -110 300 -93
rect 322 -110 330 -93
rect 292 -118 330 -110
rect 381 -93 419 -90
rect 381 -110 389 -93
rect 411 -110 419 -93
rect 381 -118 419 -110
rect 470 -93 508 -90
rect 470 -110 478 -93
rect 500 -110 508 -93
rect 470 -118 508 -110
rect 559 -93 597 -90
rect 559 -110 567 -93
rect 589 -110 597 -93
rect 559 -118 597 -110
rect 648 -93 686 -90
rect 648 -110 656 -93
rect 678 -110 686 -93
rect 648 -118 686 -110
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 1.4 l 0.6 m 1 nf 16 diffcov 100 polycov 50 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
